module real_jpeg_1140_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_62),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_1),
.B(n_35),
.Y(n_203)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_62),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_2),
.B(n_44),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_2),
.B(n_35),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_2),
.B(n_32),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_2),
.B(n_77),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_4),
.B(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_50),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_26),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_4),
.B(n_41),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_4),
.B(n_44),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_32),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_4),
.B(n_35),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_4),
.B(n_77),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_50),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_5),
.B(n_26),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_5),
.B(n_41),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_44),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_32),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_10),
.B(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_41),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_10),
.B(n_77),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_11),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_11),
.B(n_35),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_32),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_77),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_12),
.B(n_26),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_12),
.B(n_50),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_12),
.B(n_41),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_12),
.B(n_44),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_32),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_14),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_14),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_41),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_26),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_121),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_19),
.B(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_80),
.C(n_91),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_20),
.B(n_80),
.CI(n_91),
.CON(n_148),
.SN(n_148)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_59),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_21),
.B(n_60),
.C(n_71),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.C(n_46),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_22),
.A2(n_23),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_24),
.B(n_33),
.C(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_26),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_31),
.A2(n_38),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_31),
.B(n_212),
.C(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_31),
.A2(n_38),
.B1(n_212),
.B2(n_218),
.Y(n_217)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_32),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_33),
.A2(n_34),
.B1(n_76),
.B2(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_33),
.A2(n_34),
.B1(n_173),
.B2(n_251),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_74),
.C(n_76),
.Y(n_73)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_36),
.B(n_170),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_38),
.B(n_84),
.C(n_85),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_39),
.B(n_46),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_40),
.B(n_43),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_41),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_42),
.A2(n_83),
.B1(n_84),
.B2(n_94),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_42),
.B(n_84),
.C(n_192),
.Y(n_231)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_56),
.C(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_56),
.A2(n_57),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_138),
.C(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_66),
.C(n_68),
.Y(n_131)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_62),
.Y(n_171)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_114),
.C(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_67),
.B1(n_114),
.B2(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_73),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_76),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_76),
.A2(n_100),
.B1(n_268),
.B2(n_269),
.Y(n_281)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_79),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_113),
.C(n_119),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_79),
.A2(n_110),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_110),
.B1(n_119),
.B2(n_120),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_84),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_107),
.C(n_112),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_92),
.B(n_107),
.CI(n_112),
.CON(n_150),
.SN(n_150)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_103),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_93),
.B(n_97),
.Y(n_357)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_98),
.A2(n_99),
.B1(n_208),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_100),
.B(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_101),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_102),
.A2(n_184),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_103),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_115),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_115),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_142),
.B2(n_143),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_141),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_137),
.A2(n_138),
.B1(n_160),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_176),
.B(n_371),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_148),
.B(n_149),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_148),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.C(n_154),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_150),
.B(n_151),
.Y(n_359)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_150),
.Y(n_375)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_154),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.C(n_166),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_155),
.A2(n_156),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_157),
.B(n_159),
.CI(n_161),
.CON(n_333),
.SN(n_333)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_160),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_164),
.B(n_166),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.C(n_175),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_167),
.A2(n_168),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_169),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_172),
.A2(n_173),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_172),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_173),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_174),
.A2(n_175),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_174),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_175),
.Y(n_345)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI31xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_347),
.A3(n_360),
.B(n_365),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_327),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_252),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_225),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_181),
.B(n_225),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_195),
.C(n_215),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_182),
.B(n_324),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_182),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.CI(n_191),
.CON(n_182),
.SN(n_182)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_187),
.C(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_185),
.B(n_186),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_190),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_193),
.B(n_209),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_193),
.B(n_236),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_195),
.B(n_215),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_205),
.B2(n_214),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_206),
.C(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_202),
.C(n_204),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_223),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_216),
.B(n_219),
.CI(n_223),
.CON(n_314),
.SN(n_314)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_222),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_263),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_225),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_242),
.CI(n_243),
.CON(n_225),
.SN(n_225)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_226),
.B(n_242),
.C(n_243),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_227),
.B(n_230),
.C(n_237),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_237),
.B2(n_238),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_322),
.B(n_326),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_310),
.B(n_321),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_282),
.B(n_309),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_273),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_273),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_260),
.CI(n_261),
.CON(n_274),
.SN(n_274)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_262),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.C(n_281),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_306),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_274),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_303),
.B(n_308),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_294),
.B(n_302),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_297),
.B(n_301),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_299),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_317),
.C(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_328),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_346),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_346),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_332),
.C(n_335),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_340),
.C(n_341),
.Y(n_354)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g365 ( 
.A1(n_348),
.A2(n_361),
.B(n_366),
.C(n_369),
.D(n_370),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_358),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_358),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.C(n_355),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_350),
.A2(n_351),
.B1(n_355),
.B2(n_356),
.Y(n_363)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_363),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_364),
.Y(n_369)
);


endmodule