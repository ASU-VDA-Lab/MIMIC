module fake_jpeg_22576_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_22),
.Y(n_65)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_22),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_20),
.B1(n_32),
.B2(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_64),
.A2(n_29),
.B1(n_25),
.B2(n_47),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_76),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_20),
.B1(n_36),
.B2(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_20),
.B1(n_32),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_44),
.B1(n_43),
.B2(n_29),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_42),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_19),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_33),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_103),
.C(n_26),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_46),
.B1(n_33),
.B2(n_31),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_90),
.B(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_95),
.B1(n_105),
.B2(n_46),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_96),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_42),
.B1(n_38),
.B2(n_46),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_98),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_28),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_107),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_67),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_44),
.B1(n_43),
.B2(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_43),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_114),
.B1(n_26),
.B2(n_31),
.Y(n_137)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_52),
.A2(n_25),
.B1(n_42),
.B2(n_33),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_56),
.B1(n_79),
.B2(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_30),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_143),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_124),
.B1(n_133),
.B2(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_125),
.Y(n_159)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_130),
.B1(n_95),
.B2(n_94),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_132),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_68),
.B1(n_66),
.B2(n_58),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_83),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_79),
.B1(n_56),
.B2(n_18),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_68),
.B1(n_58),
.B2(n_52),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_136),
.B1(n_95),
.B2(n_86),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_26),
.B(n_13),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_9),
.B(n_16),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_101),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_96),
.A2(n_21),
.B1(n_23),
.B2(n_17),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_17),
.B1(n_37),
.B2(n_23),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_24),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_113),
.C(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_149),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_78),
.C(n_73),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_0),
.Y(n_181)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

XOR2x1_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_12),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_85),
.B(n_84),
.C(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_85),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_181),
.B(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_173),
.B1(n_179),
.B2(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_171),
.B1(n_146),
.B2(n_153),
.Y(n_212)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_121),
.A2(n_95),
.B1(n_108),
.B2(n_94),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_93),
.B(n_21),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_120),
.B(n_131),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_23),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_182),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_93),
.B1(n_21),
.B2(n_37),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_104),
.B1(n_38),
.B2(n_106),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_120),
.B(n_24),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_193),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_136),
.B1(n_143),
.B2(n_126),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_206),
.B1(n_212),
.B2(n_179),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_211),
.B(n_216),
.Y(n_229)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_203),
.Y(n_233)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_202),
.B1(n_127),
.B2(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_130),
.B1(n_151),
.B2(n_127),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_214),
.B1(n_169),
.B2(n_170),
.Y(n_219)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_207),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_151),
.B1(n_145),
.B2(n_125),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_158),
.B(n_146),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_166),
.B1(n_170),
.B2(n_163),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_1),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_181),
.B(n_185),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g216 ( 
.A(n_157),
.B(n_141),
.C(n_123),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_9),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_162),
.B(n_167),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_231),
.B1(n_237),
.B2(n_206),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_226),
.B1(n_199),
.B2(n_240),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_199),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_178),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_239),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_182),
.C(n_176),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_196),
.C(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_232),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_167),
.B1(n_162),
.B2(n_144),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_205),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_38),
.B1(n_1),
.B2(n_3),
.Y(n_237)
);

FAx1_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_38),
.CI(n_1),
.CON(n_239),
.SN(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_16),
.B(n_3),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_211),
.B1(n_201),
.B2(n_189),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_208),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_213),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_247),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_214),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_201),
.C(n_189),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_260),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_224),
.B1(n_235),
.B2(n_218),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_251),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_255),
.B(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_197),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_216),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_262),
.C(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_215),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_261),
.B1(n_247),
.B2(n_224),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_267),
.B1(n_272),
.B2(n_215),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_274),
.C(n_278),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_265),
.B(n_225),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_223),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_270),
.B(n_280),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_218),
.B(n_230),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_244),
.A2(n_239),
.B1(n_233),
.B2(n_203),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_258),
.C(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_229),
.C(n_237),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_229),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_16),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_282),
.B(n_287),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_248),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_241),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_289),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_291),
.B1(n_278),
.B2(n_270),
.Y(n_298)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_195),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_225),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_193),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_274),
.C(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_264),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_2),
.B(n_3),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_280),
.B1(n_271),
.B2(n_272),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_283),
.B1(n_285),
.B2(n_289),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_273),
.B1(n_279),
.B2(n_5),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_2),
.C(n_4),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_297),
.B(n_299),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_283),
.B(n_275),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_296),
.B(n_304),
.Y(n_315)
);

AOI31xp33_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_4),
.Y(n_312)
);

FAx1_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_303),
.CI(n_6),
.CON(n_313),
.SN(n_313)
);

AOI31xp67_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_316),
.A3(n_317),
.B(n_8),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_296),
.B(n_305),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_320),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_311),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_319),
.B(n_11),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_322),
.B1(n_11),
.B2(n_13),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_8),
.B(n_14),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_14),
.Y(n_327)
);


endmodule