module fake_jpeg_138_n_118 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_2),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_1),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_54),
.B(n_51),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_37),
.B1(n_39),
.B2(n_33),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_38),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_38),
.B1(n_33),
.B2(n_44),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_32),
.B1(n_15),
.B2(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_45),
.C(n_44),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_20),
.C(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_27),
.B(n_26),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_81),
.B1(n_74),
.B2(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_8),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_86),
.C(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_14),
.C(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_94),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_91),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_31),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_22),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_6),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.C(n_107),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_90),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_95),
.B1(n_12),
.B2(n_13),
.C(n_11),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_109),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_103),
.B1(n_101),
.B2(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_112),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_112),
.Y(n_118)
);


endmodule