module fake_netlist_5_1665_n_2084 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2084);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2084;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_8),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_139),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_22),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_86),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_0),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_87),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_90),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_57),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_40),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_116),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_66),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_104),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_191),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_123),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_40),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_51),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_119),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_35),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_70),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_82),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_138),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_126),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_106),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_175),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_69),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_151),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_48),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_37),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_84),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_22),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_67),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_74),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_128),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_15),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_44),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_32),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_74),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_115),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_32),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_54),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_107),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_166),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_81),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_102),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_85),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_77),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_113),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_142),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_91),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_66),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_89),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_62),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_98),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_82),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_122),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_67),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_48),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_78),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_16),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_8),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_95),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_177),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_162),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_144),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_45),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_44),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_120),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_135),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_133),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_61),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_12),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_154),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_64),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_28),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_20),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_27),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_47),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_26),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_155),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_17),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_77),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_140),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_99),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_92),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_153),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_36),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_55),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_187),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_168),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_63),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_21),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_165),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_178),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_34),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_9),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_33),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_52),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_27),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_96),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_172),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_20),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_167),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_103),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_149),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_161),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_7),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_53),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_94),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_148),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_52),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_30),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_58),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_110),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_19),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_109),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_9),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_194),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_6),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_111),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_35),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_5),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_6),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_134),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_73),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_59),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_164),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_189),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_18),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_81),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_105),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_2),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_58),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_51),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_50),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_124),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_93),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_42),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_1),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_285),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_226),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_219),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_285),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_227),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_285),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_199),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_2),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_285),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_200),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_305),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_201),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_285),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_260),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_222),
.B(n_5),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_285),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_391),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_212),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_227),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_285),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_285),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_285),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_216),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_217),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_220),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_221),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_267),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_202),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_208),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_232),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_359),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_234),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_202),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_202),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_222),
.B(n_7),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_202),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_202),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_202),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_218),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_218),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_250),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_218),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_218),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_218),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_265),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_250),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_265),
.B(n_10),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_231),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_310),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_218),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_245),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_248),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_243),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_247),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_251),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_339),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_255),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_271),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_339),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_274),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_281),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_339),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_339),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_283),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_288),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_390),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_279),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_237),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_237),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_293),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_237),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_237),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_237),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_215),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_215),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_243),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_289),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_292),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_379),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_233),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_233),
.B(n_13),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_268),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_268),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_296),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_361),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_298),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_312),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_197),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_315),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_197),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_205),
.B(n_13),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_321),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_293),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_205),
.B(n_14),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_399),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_204),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_467),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_398),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_441),
.B(n_207),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_393),
.B(n_229),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_402),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_404),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_247),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_449),
.B(n_264),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_469),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_394),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_203),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_469),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_411),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_416),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_466),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

CKINVDCx8_ASAP7_75t_R g523 ( 
.A(n_448),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_475),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_417),
.Y(n_529)
);

CKINVDCx11_ASAP7_75t_R g530 ( 
.A(n_422),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_429),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_418),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_466),
.B(n_204),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_419),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_423),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_432),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_425),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_466),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_445),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_447),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_433),
.B(n_330),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_396),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_450),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_454),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_433),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_434),
.B(n_335),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_401),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_442),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_438),
.B(n_340),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_401),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_457),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_462),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_443),
.B(n_240),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_405),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_444),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_407),
.B(n_207),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_407),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_446),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_460),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_403),
.B(n_211),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_547),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_523),
.B(n_395),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_501),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_508),
.B(n_473),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_521),
.B(n_213),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_507),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_502),
.B(n_480),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_448),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

INVx4_ASAP7_75t_SL g585 ( 
.A(n_503),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_521),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_521),
.B(n_489),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_521),
.B(n_484),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_526),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_508),
.B(n_572),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_528),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_502),
.B(n_485),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_526),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_526),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_513),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_487),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_521),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_513),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_490),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_569),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_530),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_513),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_543),
.Y(n_607)
);

NOR2x1p5_ASAP7_75t_L g608 ( 
.A(n_494),
.B(n_397),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_501),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_543),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_497),
.B(n_203),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_543),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_512),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_536),
.B(n_489),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_536),
.B(n_412),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_501),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_497),
.B(n_463),
.C(n_439),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_543),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_530),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_532),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_546),
.B(n_446),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_569),
.B(n_229),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_543),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_553),
.Y(n_627)
);

BUFx8_ASAP7_75t_SL g628 ( 
.A(n_511),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_563),
.B(n_472),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_410),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_501),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_536),
.B(n_470),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_532),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_505),
.B(n_453),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_518),
.B(n_456),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_497),
.B(n_470),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_552),
.B(n_451),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_563),
.B(n_520),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_541),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_552),
.B(n_451),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_501),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_559),
.B(n_452),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_554),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_501),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_529),
.B(n_461),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_535),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_547),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_512),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_553),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_537),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_553),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_559),
.B(n_553),
.Y(n_655)
);

BUFx4f_ASAP7_75t_L g656 ( 
.A(n_547),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_534),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_568),
.B(n_472),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_553),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_547),
.B(n_452),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_506),
.B(n_213),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_455),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_538),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_540),
.B(n_474),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_519),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_568),
.B(n_408),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_544),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_471),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_561),
.B(n_455),
.Y(n_672)
);

AND2x6_ASAP7_75t_SL g673 ( 
.A(n_565),
.B(n_209),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_561),
.B(n_458),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_519),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_541),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_503),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_524),
.Y(n_679)
);

OR2x2_ASAP7_75t_SL g680 ( 
.A(n_500),
.B(n_492),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_566),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_534),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_524),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_555),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_493),
.B(n_471),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_555),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_514),
.B(n_492),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_495),
.B(n_496),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_495),
.B(n_476),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_525),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_522),
.B(n_554),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_525),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_561),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_503),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_561),
.B(n_230),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_545),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_548),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_566),
.B(n_458),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_541),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_541),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_527),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_555),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_496),
.B(n_498),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_503),
.A2(n_477),
.B1(n_428),
.B2(n_214),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_527),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_531),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_531),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_229),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_533),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_503),
.B(n_229),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_549),
.B(n_406),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_566),
.B(n_459),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_533),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_562),
.B(n_420),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_556),
.Y(n_716)
);

INVxp33_ASAP7_75t_SL g717 ( 
.A(n_571),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_539),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_522),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_566),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_566),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_566),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_556),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_523),
.B(n_207),
.Y(n_725)
);

AND2x6_ASAP7_75t_SL g726 ( 
.A(n_631),
.B(n_209),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_586),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_596),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_615),
.B(n_498),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_596),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_582),
.A2(n_430),
.B1(n_424),
.B2(n_257),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_615),
.B(n_499),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_599),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_593),
.B(n_506),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_599),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_655),
.B(n_523),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_720),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_720),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_600),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_615),
.B(n_499),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_662),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_587),
.B(n_229),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_665),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_587),
.B(n_323),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_592),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_611),
.A2(n_230),
.B1(n_333),
.B2(n_301),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_611),
.A2(n_333),
.B1(n_301),
.B2(n_238),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_687),
.B(n_329),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_600),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_602),
.B(n_597),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_628),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_591),
.A2(n_477),
.B(n_400),
.C(n_224),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_587),
.B(n_323),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_586),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_641),
.B(n_223),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_598),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_579),
.B(n_323),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_611),
.A2(n_238),
.B1(n_246),
.B2(n_223),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_624),
.B(n_509),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_337),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_601),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_601),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

CKINVDCx11_ASAP7_75t_R g765 ( 
.A(n_697),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_579),
.B(n_323),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_639),
.B(n_509),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_642),
.B(n_515),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_579),
.B(n_323),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_579),
.B(n_500),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_633),
.B(n_246),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_592),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_644),
.B(n_515),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_603),
.B(n_486),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_665),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_671),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_611),
.A2(n_309),
.B1(n_371),
.B2(n_244),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_638),
.B(n_539),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_638),
.B(n_542),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_671),
.Y(n_781)
);

NOR2x2_ASAP7_75t_L g782 ( 
.A(n_673),
.B(n_500),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_687),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_611),
.B(n_542),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_611),
.B(n_550),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_685),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_685),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_689),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_659),
.A2(n_278),
.B1(n_282),
.B2(n_252),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_611),
.A2(n_278),
.B1(n_282),
.B2(n_252),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_663),
.A2(n_291),
.B1(n_300),
.B2(n_287),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_584),
.B(n_500),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_663),
.A2(n_224),
.B(n_235),
.C(n_214),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_616),
.B(n_550),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_692),
.B(n_279),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_616),
.B(n_551),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_668),
.B(n_551),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_614),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_668),
.B(n_557),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_676),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_676),
.B(n_557),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_576),
.A2(n_357),
.B1(n_344),
.B2(n_345),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_584),
.B(n_500),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_SL g805 ( 
.A(n_629),
.B(n_210),
.C(n_198),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_669),
.B(n_225),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_679),
.B(n_558),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_663),
.A2(n_348),
.B(n_254),
.C(n_256),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_679),
.B(n_558),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_669),
.B(n_228),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_633),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_683),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_688),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_619),
.B(n_236),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_683),
.B(n_560),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_583),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_690),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_688),
.Y(n_818)
);

NOR2x1p5_ASAP7_75t_L g819 ( 
.A(n_659),
.B(n_239),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_583),
.A2(n_351),
.B1(n_341),
.B2(n_311),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_690),
.B(n_560),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_590),
.B(n_352),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_608),
.A2(n_358),
.B1(n_355),
.B2(n_356),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_693),
.Y(n_824)
);

AND2x6_ASAP7_75t_SL g825 ( 
.A(n_636),
.B(n_235),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_704),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_704),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_590),
.B(n_362),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_693),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_702),
.B(n_570),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_650),
.A2(n_291),
.B1(n_351),
.B2(n_300),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_702),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_608),
.A2(n_367),
.B1(n_363),
.B2(n_389),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_594),
.B(n_369),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_706),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_706),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_707),
.B(n_708),
.Y(n_837)
);

BUFx12f_ASAP7_75t_L g838 ( 
.A(n_697),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_588),
.A2(n_381),
.B1(n_377),
.B2(n_206),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_594),
.B(n_405),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_692),
.B(n_486),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_707),
.B(n_570),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_725),
.B(n_241),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_708),
.B(n_503),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_719),
.B(n_488),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_710),
.B(n_714),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_710),
.B(n_503),
.Y(n_847)
);

AND2x6_ASAP7_75t_SL g848 ( 
.A(n_637),
.B(n_647),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_691),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_714),
.B(n_503),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_718),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_700),
.B(n_701),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_595),
.B(n_409),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_648),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_718),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_607),
.B(n_287),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_645),
.B(n_488),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_607),
.B(n_311),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_610),
.B(n_318),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_663),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_697),
.B(n_476),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_630),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_610),
.B(n_318),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_613),
.B(n_319),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_595),
.B(n_409),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_613),
.B(n_319),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_648),
.B(n_652),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_620),
.B(n_334),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_620),
.B(n_334),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_626),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_626),
.B(n_413),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_627),
.B(n_242),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_598),
.A2(n_380),
.B1(n_336),
.B2(n_341),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_627),
.B(n_336),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_651),
.B(n_249),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_651),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_654),
.B(n_253),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_654),
.B(n_373),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_660),
.A2(n_373),
.B1(n_380),
.B2(n_206),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_717),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_660),
.B(n_413),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_577),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_581),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_720),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_577),
.Y(n_885)
);

BUFx5_ASAP7_75t_L g886 ( 
.A(n_696),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_581),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_618),
.B(n_510),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_575),
.B(n_609),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_667),
.B(n_254),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_678),
.B(n_414),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_575),
.B(n_609),
.Y(n_892)
);

CKINVDCx11_ASAP7_75t_R g893 ( 
.A(n_717),
.Y(n_893)
);

BUFx8_ASAP7_75t_L g894 ( 
.A(n_700),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_575),
.B(n_510),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_640),
.B(n_262),
.C(n_258),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_652),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_724),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_751),
.B(n_609),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_SL g900 ( 
.A1(n_806),
.A2(n_666),
.B1(n_698),
.B2(n_670),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_728),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_740),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_783),
.B(n_666),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_857),
.B(n_670),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_755),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_734),
.B(n_643),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_854),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_794),
.B(n_643),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_746),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_740),
.Y(n_910)
);

AO22x1_ASAP7_75t_L g911 ( 
.A1(n_843),
.A2(n_698),
.B1(n_715),
.B2(n_712),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_730),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_742),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_733),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_860),
.A2(n_705),
.B1(n_625),
.B2(n_578),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_742),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_744),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_755),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_755),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_796),
.B(n_643),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_775),
.B(n_574),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_727),
.A2(n_656),
.B(n_589),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_838),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_845),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_838),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_727),
.B(n_649),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_816),
.B(n_680),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_772),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_755),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_735),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_744),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_897),
.Y(n_932)
);

INVx3_ASAP7_75t_SL g933 ( 
.A(n_752),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_849),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_776),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_776),
.Y(n_937)
);

NAND2x1_ASAP7_75t_L g938 ( 
.A(n_737),
.B(n_738),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_750),
.A2(n_578),
.B1(n_580),
.B2(n_701),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_SL g940 ( 
.A(n_820),
.B(n_621),
.C(n_605),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_801),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_801),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_757),
.B(n_678),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_835),
.B(n_649),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_836),
.B(n_851),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_757),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_757),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_762),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_855),
.B(n_649),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_R g950 ( 
.A(n_893),
.B(n_605),
.Y(n_950)
);

BUFx6f_ASAP7_75t_SL g951 ( 
.A(n_880),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_763),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_764),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_805),
.B(n_261),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_799),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_765),
.B(n_621),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_774),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_757),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_898),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_813),
.A2(n_818),
.B1(n_827),
.B2(n_826),
.Y(n_960)
);

CKINVDCx14_ASAP7_75t_R g961 ( 
.A(n_867),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_898),
.Y(n_962)
);

INVx3_ASAP7_75t_SL g963 ( 
.A(n_782),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_792),
.B(n_290),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_795),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_837),
.B(n_721),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_795),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_737),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_736),
.B(n_680),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_738),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_736),
.A2(n_822),
.B1(n_834),
.B2(n_828),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_812),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_817),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_SL g975 ( 
.A(n_792),
.B(n_327),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_824),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_862),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_811),
.B(n_641),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_SL g979 ( 
.A(n_831),
.B(n_266),
.C(n_263),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_777),
.B(n_657),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_884),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_824),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_829),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_848),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_761),
.B(n_806),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_771),
.A2(n_580),
.B1(n_696),
.B2(n_604),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_829),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_884),
.Y(n_988)
);

CKINVDCx11_ASAP7_75t_R g989 ( 
.A(n_825),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_832),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_880),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_832),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_810),
.A2(n_326),
.B(n_325),
.C(n_324),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_894),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_849),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_771),
.A2(n_696),
.B1(n_604),
.B2(n_612),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_795),
.B(n_657),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_890),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_870),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_846),
.B(n_721),
.Y(n_1000)
);

BUFx4f_ASAP7_75t_L g1001 ( 
.A(n_890),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_779),
.B(n_721),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_780),
.B(n_630),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_781),
.B(n_677),
.Y(n_1004)
);

CKINVDCx6p67_ASAP7_75t_R g1005 ( 
.A(n_890),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_882),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_761),
.B(n_786),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_SL g1008 ( 
.A(n_789),
.B(n_270),
.C(n_269),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_876),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_787),
.B(n_630),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_729),
.A2(n_656),
.B(n_589),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_R g1012 ( 
.A(n_749),
.B(n_841),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_810),
.B(n_573),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_731),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_788),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_882),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_886),
.B(n_678),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_756),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_814),
.A2(n_677),
.B(n_275),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_798),
.B(n_585),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_771),
.B(n_585),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_885),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_885),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_756),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_883),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_861),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_887),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_852),
.B(n_272),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_732),
.Y(n_1029)
);

AO22x1_ASAP7_75t_L g1030 ( 
.A1(n_843),
.A2(n_814),
.B1(n_896),
.B2(n_894),
.Y(n_1030)
);

AO22x1_ASAP7_75t_L g1031 ( 
.A1(n_894),
.A2(n_320),
.B1(n_322),
.B2(n_317),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_756),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_797),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_741),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_800),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_791),
.A2(n_324),
.B1(n_313),
.B2(n_302),
.C(n_284),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_802),
.Y(n_1037)
);

BUFx8_ASAP7_75t_SL g1038 ( 
.A(n_726),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_753),
.B(n_277),
.C(n_276),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_R g1040 ( 
.A(n_756),
.B(n_280),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_886),
.B(n_678),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_756),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_803),
.B(n_294),
.C(n_286),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_872),
.B(n_573),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_807),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_760),
.B(n_630),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_889),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_822),
.A2(n_681),
.B1(n_573),
.B2(n_694),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_892),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_759),
.A2(n_696),
.B1(n_612),
.B2(n_617),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_767),
.B(n_630),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_872),
.B(n_622),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_886),
.B(n_678),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_886),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_768),
.B(n_632),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_886),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_773),
.B(n_632),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_809),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_770),
.B(n_585),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_871),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_815),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_821),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_819),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_830),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_875),
.B(n_622),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_842),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_871),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_753),
.B(n_297),
.C(n_295),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_881),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_875),
.B(n_877),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_877),
.B(n_632),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_881),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_840),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_873),
.B(n_632),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_770),
.B(n_585),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_828),
.A2(n_622),
.B1(n_634),
.B2(n_694),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_834),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_840),
.B(n_632),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_853),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_853),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_804),
.B(n_634),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_823),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_793),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_793),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_R g1086 ( 
.A(n_784),
.B(n_785),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_808),
.A2(n_709),
.B(n_711),
.C(n_713),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_808),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_865),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_856),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_865),
.B(n_646),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1054),
.A2(n_1057),
.B(n_1056),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_985),
.A2(n_804),
.B(n_743),
.C(n_754),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_985),
.B(n_839),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1037),
.B(n_778),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_922),
.A2(n_859),
.B(n_858),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_902),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_L g1098 ( 
.A(n_1014),
.B(n_833),
.C(n_790),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_935),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_904),
.B(n_743),
.Y(n_1100)
);

CKINVDCx14_ASAP7_75t_R g1101 ( 
.A(n_950),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1011),
.A2(n_864),
.B(n_863),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1054),
.A2(n_868),
.B(n_866),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_932),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1054),
.A2(n_656),
.B(n_589),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_902),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1056),
.A2(n_1057),
.B(n_926),
.Y(n_1107)
);

AND2x2_ASAP7_75t_SL g1108 ( 
.A(n_1071),
.B(n_748),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_1013),
.A2(n_754),
.B(n_745),
.C(n_766),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_1072),
.A2(n_874),
.B(n_869),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_899),
.A2(n_745),
.B(n_844),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1056),
.A2(n_878),
.B(n_850),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1057),
.A2(n_675),
.B(n_747),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_972),
.B(n_847),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1044),
.A2(n_766),
.B(n_758),
.Y(n_1115)
);

AO21x1_ASAP7_75t_L g1116 ( 
.A1(n_964),
.A2(n_769),
.B(n_758),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_969),
.Y(n_1117)
);

OA22x2_ASAP7_75t_L g1118 ( 
.A1(n_924),
.A2(n_256),
.B1(n_259),
.B2(n_273),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_910),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1045),
.B(n_1059),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_993),
.A2(n_769),
.B(n_348),
.C(n_347),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_970),
.A2(n_879),
.B(n_259),
.C(n_273),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_969),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1003),
.A2(n_895),
.B(n_888),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_945),
.A2(n_664),
.B(n_661),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_969),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1091),
.A2(n_674),
.B(n_672),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1063),
.B(n_891),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1079),
.A2(n_699),
.B(n_891),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_995),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_910),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_991),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1026),
.B(n_478),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1044),
.A2(n_675),
.B(n_634),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_900),
.A2(n_302),
.B(n_284),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1052),
.A2(n_675),
.B(n_623),
.Y(n_1136)
);

OA22x2_ASAP7_75t_L g1137 ( 
.A1(n_1083),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_913),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_913),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_984),
.A2(n_306),
.B1(n_299),
.B2(n_303),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_973),
.A2(n_682),
.B(n_617),
.Y(n_1141)
);

NAND2x1_ASAP7_75t_L g1142 ( 
.A(n_969),
.B(n_646),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_SL g1143 ( 
.A1(n_1061),
.A2(n_332),
.B(n_342),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_906),
.A2(n_686),
.B(n_623),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_973),
.A2(n_684),
.B(n_635),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_973),
.A2(n_684),
.B(n_635),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_955),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_971),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1012),
.B(n_304),
.C(n_307),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1052),
.A2(n_686),
.B(n_653),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1067),
.B(n_1033),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_921),
.B(n_903),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_991),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1012),
.B(n_392),
.C(n_346),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_992),
.A2(n_653),
.B(n_658),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_992),
.A2(n_658),
.B(n_682),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_993),
.A2(n_703),
.A3(n_716),
.B(n_332),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_992),
.A2(n_703),
.B(n_716),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1066),
.A2(n_724),
.B(n_694),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_724),
.B(n_342),
.C(n_343),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1066),
.A2(n_646),
.B(n_722),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_909),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_908),
.A2(n_920),
.B(n_1002),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_646),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1061),
.A2(n_343),
.B(n_365),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1035),
.B(n_1062),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_970),
.A2(n_383),
.B(n_347),
.C(n_365),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1046),
.A2(n_646),
.B(n_722),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1035),
.B(n_720),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1062),
.B(n_720),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_928),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_916),
.A2(n_459),
.B(n_556),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_1007),
.A2(n_376),
.B(n_308),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_903),
.Y(n_1174)
);

CKINVDCx11_ASAP7_75t_R g1175 ( 
.A(n_933),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_916),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_907),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_932),
.B(n_83),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_954),
.A2(n_378),
.B1(n_314),
.B2(n_331),
.C(n_338),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_950),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1065),
.A2(n_1034),
.B1(n_1029),
.B2(n_1061),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1065),
.B(n_722),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_901),
.B(n_722),
.Y(n_1183)
);

INVx3_ASAP7_75t_SL g1184 ( 
.A(n_933),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_912),
.B(n_722),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1084),
.A2(n_368),
.A3(n_374),
.B(n_382),
.Y(n_1186)
);

AOI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1083),
.A2(n_1078),
.B(n_1019),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1051),
.A2(n_723),
.B(n_678),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1055),
.A2(n_723),
.B(n_695),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1073),
.A2(n_723),
.B1(n_695),
.B2(n_316),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1080),
.B(n_723),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_917),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_917),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_911),
.B(n_328),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_914),
.B(n_723),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1073),
.A2(n_695),
.B1(n_386),
.B2(n_350),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_930),
.B(n_353),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_931),
.A2(n_564),
.B(n_567),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_934),
.B(n_948),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_952),
.B(n_953),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1058),
.A2(n_695),
.B(n_567),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_957),
.B(n_354),
.Y(n_1202)
);

AOI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_954),
.A2(n_388),
.B1(n_360),
.B2(n_364),
.C(n_366),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_960),
.B(n_370),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_931),
.A2(n_564),
.B(n_567),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1068),
.A2(n_696),
.B(n_414),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_961),
.B(n_478),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1015),
.B(n_479),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_936),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_977),
.A2(n_1000),
.B(n_967),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_961),
.B(n_479),
.Y(n_1211)
);

OAI22x1_ASAP7_75t_L g1212 ( 
.A1(n_927),
.A2(n_375),
.B1(n_372),
.B2(n_374),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_929),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_936),
.A2(n_990),
.A3(n_942),
.B(n_941),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1090),
.B(n_510),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1090),
.B(n_510),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_999),
.B(n_368),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1009),
.B(n_382),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_937),
.A2(n_564),
.B(n_415),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_937),
.A2(n_415),
.B(n_482),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_941),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_942),
.A2(n_482),
.B(n_481),
.Y(n_1222)
);

AND2x6_ASAP7_75t_SL g1223 ( 
.A(n_927),
.B(n_383),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_984),
.A2(n_387),
.B1(n_385),
.B2(n_481),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_1043),
.B(n_88),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_976),
.A2(n_385),
.B(n_387),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1075),
.A2(n_695),
.B(n_696),
.Y(n_1227)
);

AO21x1_ASAP7_75t_L g1228 ( 
.A1(n_964),
.A2(n_207),
.B(n_696),
.Y(n_1228)
);

AOI21xp33_ASAP7_75t_L g1229 ( 
.A1(n_1070),
.A2(n_14),
.B(n_15),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_976),
.A2(n_160),
.B(n_196),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_982),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_982),
.A2(n_159),
.B(n_195),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_971),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1088),
.B(n_695),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_965),
.B(n_17),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1080),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_990),
.A2(n_193),
.B(n_188),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_966),
.B(n_19),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_1086),
.A2(n_183),
.B(n_182),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_974),
.B(n_21),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_944),
.A2(n_181),
.B(n_174),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_983),
.B(n_23),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_949),
.A2(n_171),
.B(n_170),
.Y(n_1243)
);

NOR2xp67_ASAP7_75t_L g1244 ( 
.A(n_907),
.B(n_152),
.Y(n_1244)
);

NAND3x1_ASAP7_75t_L g1245 ( 
.A(n_1036),
.B(n_23),
.C(n_24),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_SL g1246 ( 
.A1(n_1073),
.A2(n_146),
.B(n_141),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_987),
.B(n_24),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1074),
.A2(n_28),
.A3(n_29),
.B(n_30),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1047),
.B(n_29),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_971),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_938),
.A2(n_132),
.B(n_130),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_975),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1022),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1016),
.A2(n_117),
.B(n_114),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_971),
.A2(n_108),
.B(n_101),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1148),
.B(n_980),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1100),
.B(n_1039),
.Y(n_1257)
);

INVx8_ASAP7_75t_L g1258 ( 
.A(n_1148),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1198),
.A2(n_1010),
.B(n_1023),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1198),
.A2(n_1205),
.B(n_1172),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1205),
.A2(n_1023),
.B(n_1016),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1200),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1103),
.A2(n_1027),
.B(n_1025),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1104),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1180),
.B(n_925),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1214),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1152),
.A2(n_975),
.B1(n_1001),
.B2(n_998),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1214),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1166),
.B(n_1069),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1214),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1252),
.A2(n_1008),
.B(n_1064),
.C(n_979),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1120),
.B(n_978),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1252),
.A2(n_963),
.B(n_940),
.C(n_968),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1172),
.A2(n_1016),
.B(n_1023),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1099),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1214),
.Y(n_1276)
);

CKINVDCx9p33_ASAP7_75t_R g1277 ( 
.A(n_1132),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1151),
.B(n_978),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1219),
.A2(n_1087),
.B(n_1006),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1175),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1108),
.B(n_1006),
.Y(n_1281)
);

AOI221xp5_ASAP7_75t_L g1282 ( 
.A1(n_1135),
.A2(n_1212),
.B1(n_1194),
.B2(n_1187),
.C(n_1167),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1174),
.B(n_1005),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1116),
.A2(n_1074),
.A3(n_918),
.B(n_919),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1131),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1148),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1108),
.B(n_1020),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1219),
.A2(n_1048),
.B(n_962),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1098),
.A2(n_1085),
.B1(n_1001),
.B2(n_998),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1148),
.B(n_980),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1136),
.A2(n_1086),
.B(n_1077),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1094),
.A2(n_1095),
.B1(n_1199),
.B2(n_1181),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1130),
.B(n_1147),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1131),
.Y(n_1294)
);

AOI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1144),
.A2(n_1114),
.B(n_1134),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1253),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1236),
.B(n_1020),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1194),
.A2(n_1085),
.B1(n_978),
.B2(n_1004),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1249),
.B(n_1030),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1107),
.A2(n_959),
.B(n_962),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1117),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_SL g1302 ( 
.A1(n_1143),
.A2(n_1074),
.B(n_918),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1175),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1097),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1093),
.A2(n_915),
.B(n_1082),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1228),
.A2(n_918),
.A3(n_919),
.B(n_1082),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1107),
.A2(n_962),
.B(n_959),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_SL g1308 ( 
.A1(n_1165),
.A2(n_919),
.B(n_939),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1199),
.B(n_980),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1210),
.A2(n_1018),
.B(n_1032),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1106),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1220),
.A2(n_1145),
.B(n_1141),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1117),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1128),
.A2(n_947),
.B1(n_929),
.B2(n_958),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1138),
.B(n_1020),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1220),
.A2(n_959),
.B(n_905),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1138),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1103),
.A2(n_1082),
.B(n_943),
.Y(n_1318)
);

BUFx2_ASAP7_75t_SL g1319 ( 
.A(n_1117),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1115),
.A2(n_929),
.B1(n_958),
.B2(n_1018),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1176),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1226),
.A2(n_1050),
.B(n_996),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1117),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1176),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1204),
.A2(n_929),
.B1(n_958),
.B2(n_1018),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1141),
.A2(n_946),
.B(n_905),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1192),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1192),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1123),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1217),
.B(n_1004),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1213),
.B(n_1004),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1119),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1213),
.B(n_1021),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1231),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_1099),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1226),
.A2(n_986),
.B(n_943),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1145),
.A2(n_905),
.B(n_946),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1162),
.A2(n_958),
.B1(n_1032),
.B2(n_1018),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1101),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1213),
.B(n_1021),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1231),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1159),
.A2(n_1040),
.B(n_1028),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1109),
.A2(n_1076),
.B(n_1060),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1139),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1146),
.A2(n_946),
.B(n_1017),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1193),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1114),
.A2(n_1076),
.B(n_1060),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1218),
.B(n_1049),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1173),
.B(n_1049),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1209),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1221),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1146),
.A2(n_1017),
.B(n_1053),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1163),
.A2(n_1040),
.B(n_1028),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1149),
.A2(n_951),
.B1(n_956),
.B2(n_994),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1222),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1164),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1169),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1155),
.A2(n_1053),
.B(n_1041),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1208),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1222),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1155),
.A2(n_1041),
.B(n_1049),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1162),
.A2(n_1032),
.B1(n_981),
.B2(n_988),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1160),
.A2(n_1076),
.B(n_1060),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1156),
.A2(n_1049),
.B(n_1047),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1161),
.A2(n_997),
.B(n_1021),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1156),
.A2(n_1047),
.B(n_1032),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1133),
.B(n_1047),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1207),
.A2(n_951),
.B1(n_923),
.B2(n_997),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1211),
.A2(n_997),
.B1(n_963),
.B2(n_1031),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1158),
.A2(n_1042),
.B(n_1024),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1123),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1167),
.B(n_988),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1238),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1123),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1177),
.B(n_994),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1170),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1251),
.B(n_988),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1123),
.B(n_1042),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1153),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1182),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1158),
.A2(n_1042),
.B(n_1024),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1234),
.A2(n_988),
.B1(n_981),
.B2(n_1024),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1154),
.A2(n_956),
.B1(n_925),
.B2(n_1024),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1240),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1112),
.A2(n_1042),
.B(n_981),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1179),
.A2(n_989),
.B1(n_1038),
.B2(n_981),
.C(n_42),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1126),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1112),
.A2(n_97),
.B(n_39),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1127),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1125),
.A2(n_38),
.B(n_39),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1126),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1113),
.A2(n_989),
.B1(n_1038),
.B2(n_43),
.Y(n_1392)
);

CKINVDCx6p67_ASAP7_75t_R g1393 ( 
.A(n_1184),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1137),
.B(n_38),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1096),
.A2(n_41),
.B(n_43),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1171),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1171),
.B(n_41),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1127),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1150),
.A2(n_46),
.B(n_49),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1102),
.A2(n_46),
.B(n_49),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1126),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1129),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1129),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1096),
.A2(n_53),
.B(n_54),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1246),
.A2(n_56),
.B(n_57),
.Y(n_1405)
);

AOI222xp33_ASAP7_75t_L g1406 ( 
.A1(n_1140),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.C1(n_61),
.C2(n_63),
.Y(n_1406)
);

NAND2x1_ASAP7_75t_L g1407 ( 
.A(n_1126),
.B(n_80),
.Y(n_1407)
);

AOI22x1_ASAP7_75t_L g1408 ( 
.A1(n_1111),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1203),
.B(n_65),
.C(n_68),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1102),
.A2(n_1191),
.B(n_1124),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1229),
.A2(n_1202),
.B1(n_1197),
.B2(n_1235),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1242),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1137),
.B(n_71),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1124),
.A2(n_71),
.B(n_73),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1247),
.A2(n_75),
.B(n_76),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1105),
.A2(n_75),
.B(n_76),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1157),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1191),
.A2(n_79),
.B(n_80),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1230),
.A2(n_1237),
.B(n_1232),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1230),
.A2(n_1237),
.B(n_1232),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1215),
.A2(n_1216),
.B(n_1122),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1157),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1104),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1122),
.A2(n_1225),
.B(n_1121),
.C(n_1244),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1184),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1178),
.A2(n_1118),
.B1(n_1180),
.B2(n_1224),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1359),
.B(n_1118),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1257),
.B(n_1101),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1292),
.B(n_1250),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1275),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1305),
.A2(n_1239),
.B(n_1168),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1275),
.B(n_1186),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1257),
.B(n_1186),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1331),
.B(n_1250),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1406),
.A2(n_1239),
.B1(n_1245),
.B2(n_1255),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1386),
.A2(n_1245),
.B1(n_1195),
.B2(n_1185),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1296),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1269),
.B(n_1186),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1424),
.A2(n_1342),
.B(n_1353),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1309),
.B(n_1223),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1304),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_R g1442 ( 
.A(n_1287),
.B(n_1110),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1286),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1408),
.A2(n_1251),
.B1(n_1254),
.B2(n_1206),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1311),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1399),
.A2(n_1254),
.B(n_1243),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_L g1447 ( 
.A(n_1262),
.B(n_1233),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1264),
.Y(n_1448)
);

INVxp33_ASAP7_75t_L g1449 ( 
.A(n_1293),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1335),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1331),
.B(n_1233),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1280),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1379),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1267),
.A2(n_1196),
.B1(n_1190),
.B2(n_1183),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1408),
.A2(n_1248),
.B1(n_1243),
.B2(n_1241),
.Y(n_1455)
);

AO21x1_ASAP7_75t_L g1456 ( 
.A1(n_1418),
.A2(n_1241),
.B(n_1092),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1282),
.B(n_1409),
.C(n_1411),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1272),
.B(n_1250),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1394),
.A2(n_1110),
.B1(n_1250),
.B2(n_1233),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1394),
.A2(n_1110),
.B1(n_1201),
.B2(n_1227),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1269),
.B(n_1186),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1289),
.A2(n_1142),
.B1(n_1188),
.B2(n_1189),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1285),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1367),
.B(n_1396),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1373),
.B(n_1157),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1264),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1421),
.A2(n_1157),
.B(n_1248),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1280),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1332),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1286),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1367),
.B(n_1248),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1313),
.B(n_1248),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1277),
.Y(n_1473)
);

AOI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1384),
.A2(n_1412),
.B(n_1271),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1344),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1278),
.B(n_1375),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1392),
.A2(n_1369),
.B1(n_1273),
.B2(n_1298),
.C(n_1354),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1413),
.A2(n_1415),
.B1(n_1426),
.B2(n_1342),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1346),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1425),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1413),
.B(n_1287),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1283),
.A2(n_1330),
.B1(n_1375),
.B2(n_1368),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1310),
.A2(n_1291),
.B(n_1342),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1423),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1291),
.A2(n_1353),
.B(n_1320),
.Y(n_1485)
);

CKINVDCx6p67_ASAP7_75t_R g1486 ( 
.A(n_1393),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1425),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1258),
.B(n_1347),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1350),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1317),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1351),
.B(n_1348),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1281),
.B(n_1356),
.Y(n_1492)
);

INVx4_ASAP7_75t_SL g1493 ( 
.A(n_1286),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1281),
.B(n_1299),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1397),
.A2(n_1415),
.B1(n_1416),
.B2(n_1405),
.C(n_1372),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1315),
.B(n_1331),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1353),
.A2(n_1390),
.B1(n_1265),
.B2(n_1291),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1294),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1256),
.B(n_1290),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1266),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1303),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1419),
.A2(n_1420),
.B(n_1260),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1315),
.B(n_1297),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1299),
.A2(n_1390),
.B1(n_1405),
.B2(n_1297),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1299),
.A2(n_1390),
.B1(n_1400),
.B2(n_1356),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1303),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1357),
.B(n_1376),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1258),
.B(n_1299),
.Y(n_1508)
);

AO31x2_ASAP7_75t_L g1509 ( 
.A1(n_1417),
.A2(n_1422),
.A3(n_1389),
.B(n_1398),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1383),
.A2(n_1393),
.B1(n_1339),
.B2(n_1349),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1294),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1400),
.A2(n_1343),
.B1(n_1322),
.B2(n_1258),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1400),
.A2(n_1380),
.B1(n_1376),
.B2(n_1357),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1382),
.A2(n_1377),
.B(n_1325),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1324),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1380),
.A2(n_1256),
.B1(n_1290),
.B2(n_1339),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1258),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1333),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1321),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1327),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1256),
.B(n_1290),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1328),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1407),
.A2(n_1422),
.B1(n_1417),
.B2(n_1308),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1328),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1407),
.A2(n_1308),
.B1(n_1334),
.B2(n_1341),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1419),
.A2(n_1420),
.B(n_1414),
.Y(n_1526)
);

AOI22x1_ASAP7_75t_L g1527 ( 
.A1(n_1302),
.A2(n_1377),
.B1(n_1398),
.B2(n_1389),
.Y(n_1527)
);

OAI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1314),
.A2(n_1365),
.B1(n_1377),
.B2(n_1362),
.C(n_1338),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1341),
.B(n_1334),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1365),
.A2(n_1363),
.B1(n_1295),
.B2(n_1263),
.C(n_1329),
.Y(n_1530)
);

NAND4xp25_ASAP7_75t_L g1531 ( 
.A(n_1371),
.B(n_1333),
.C(n_1340),
.D(n_1374),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1387),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1333),
.B(n_1340),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1268),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1340),
.B(n_1378),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1260),
.A2(n_1312),
.B(n_1385),
.Y(n_1536)
);

NAND2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1286),
.B(n_1378),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1387),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1268),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1302),
.A2(n_1363),
.B1(n_1414),
.B2(n_1276),
.Y(n_1540)
);

OAI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1363),
.A2(n_1295),
.B1(n_1263),
.B2(n_1329),
.C(n_1323),
.Y(n_1541)
);

OAI22x1_ASAP7_75t_L g1542 ( 
.A1(n_1263),
.A2(n_1402),
.B1(n_1403),
.B2(n_1270),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1371),
.B(n_1323),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1371),
.B(n_1378),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1270),
.A2(n_1276),
.B1(n_1395),
.B2(n_1404),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1279),
.Y(n_1546)
);

INVx4_ASAP7_75t_SL g1547 ( 
.A(n_1286),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_SL g1548 ( 
.A1(n_1402),
.A2(n_1403),
.B(n_1355),
.C(n_1360),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1284),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1313),
.A2(n_1319),
.B1(n_1387),
.B2(n_1322),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1387),
.A2(n_1374),
.B1(n_1319),
.B2(n_1318),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1322),
.A2(n_1313),
.B1(n_1374),
.B2(n_1401),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1313),
.B(n_1391),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1301),
.Y(n_1554)
);

AO31x2_ASAP7_75t_L g1555 ( 
.A1(n_1355),
.A2(n_1360),
.A3(n_1410),
.B(n_1395),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1301),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1318),
.A2(n_1401),
.B1(n_1391),
.B2(n_1301),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1313),
.B(n_1401),
.Y(n_1558)
);

AO21x1_ASAP7_75t_L g1559 ( 
.A1(n_1404),
.A2(n_1388),
.B(n_1288),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1388),
.A2(n_1336),
.B1(n_1401),
.B2(n_1391),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1318),
.A2(n_1336),
.B1(n_1279),
.B2(n_1410),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1284),
.Y(n_1562)
);

AOI222xp33_ASAP7_75t_L g1563 ( 
.A1(n_1301),
.A2(n_1391),
.B1(n_1401),
.B2(n_1288),
.C1(n_1307),
.C2(n_1300),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1391),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1336),
.A2(n_1410),
.B1(n_1307),
.B2(n_1300),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1568)
);

INVx8_ASAP7_75t_L g1569 ( 
.A(n_1306),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1306),
.A2(n_1385),
.B1(n_1361),
.B2(n_1370),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1366),
.A2(n_1364),
.B(n_1370),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1361),
.B(n_1337),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1274),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1381),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1381),
.B(n_1316),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1326),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1366),
.A2(n_1364),
.B1(n_1274),
.B2(n_1316),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_L g1578 ( 
.A(n_1326),
.B(n_1337),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1345),
.B(n_1261),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1261),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1259),
.B(n_1345),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1259),
.B(n_1358),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1352),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1352),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1358),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1312),
.Y(n_1586)
);

CKINVDCx6p67_ASAP7_75t_R g1587 ( 
.A(n_1393),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1262),
.B(n_985),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1457),
.A2(n_1477),
.B1(n_1435),
.B2(n_1440),
.C(n_1495),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1440),
.A2(n_1435),
.B1(n_1436),
.B2(n_1474),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1588),
.A2(n_1510),
.B1(n_1449),
.B2(n_1473),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1478),
.A2(n_1485),
.B(n_1447),
.C(n_1454),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1436),
.A2(n_1478),
.B1(n_1427),
.B2(n_1482),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1437),
.Y(n_1594)
);

AND4x1_ASAP7_75t_L g1595 ( 
.A(n_1428),
.B(n_1504),
.C(n_1439),
.D(n_1438),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1467),
.A2(n_1504),
.B1(n_1449),
.B2(n_1433),
.C(n_1461),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1516),
.A2(n_1508),
.B1(n_1450),
.B2(n_1453),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1476),
.B(n_1492),
.Y(n_1599)
);

OAI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1508),
.A2(n_1507),
.B1(n_1488),
.B2(n_1484),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1508),
.A2(n_1488),
.B1(n_1587),
.B2(n_1486),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1488),
.A2(n_1432),
.B1(n_1471),
.B2(n_1430),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1429),
.A2(n_1489),
.B1(n_1469),
.B2(n_1441),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1502),
.A2(n_1536),
.B(n_1527),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1483),
.A2(n_1429),
.B(n_1552),
.Y(n_1605)
);

OAI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1531),
.A2(n_1491),
.B1(n_1487),
.B2(n_1480),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1466),
.Y(n_1607)
);

AOI211xp5_ASAP7_75t_L g1608 ( 
.A1(n_1446),
.A2(n_1456),
.B(n_1528),
.C(n_1462),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1499),
.A2(n_1521),
.B1(n_1468),
.B2(n_1506),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1497),
.A2(n_1444),
.B1(n_1460),
.B2(n_1505),
.C(n_1455),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1466),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1465),
.B(n_1445),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1499),
.A2(n_1521),
.B1(n_1501),
.B2(n_1452),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1480),
.Y(n_1614)
);

AOI222xp33_ASAP7_75t_L g1615 ( 
.A1(n_1475),
.A2(n_1479),
.B1(n_1496),
.B2(n_1458),
.C1(n_1487),
.C2(n_1505),
.Y(n_1615)
);

AOI321xp33_ASAP7_75t_L g1616 ( 
.A1(n_1460),
.A2(n_1513),
.A3(n_1459),
.B1(n_1525),
.B2(n_1523),
.C(n_1550),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1443),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1518),
.A2(n_1497),
.B1(n_1535),
.B2(n_1533),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1537),
.A2(n_1518),
.B1(n_1448),
.B2(n_1451),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1444),
.A2(n_1431),
.B1(n_1498),
.B2(n_1522),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1511),
.B(n_1515),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1431),
.A2(n_1524),
.B1(n_1520),
.B2(n_1455),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1569),
.A2(n_1514),
.B1(n_1517),
.B2(n_1472),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1512),
.A2(n_1532),
.B1(n_1472),
.B2(n_1538),
.Y(n_1624)
);

OAI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1513),
.A2(n_1512),
.B(n_1560),
.C(n_1551),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1557),
.A2(n_1530),
.B(n_1529),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1517),
.A2(n_1434),
.B1(n_1451),
.B2(n_1553),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1543),
.B(n_1434),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1537),
.A2(n_1463),
.B1(n_1519),
.B2(n_1490),
.Y(n_1629)
);

AOI321xp33_ASAP7_75t_L g1630 ( 
.A1(n_1552),
.A2(n_1541),
.A3(n_1567),
.B1(n_1540),
.B2(n_1566),
.C(n_1568),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1490),
.A2(n_1519),
.B1(n_1549),
.B2(n_1562),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_SL g1632 ( 
.A1(n_1569),
.A2(n_1443),
.B1(n_1470),
.B2(n_1566),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1534),
.A2(n_1539),
.B1(n_1500),
.B2(n_1470),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1443),
.A2(n_1470),
.B1(n_1560),
.B2(n_1556),
.Y(n_1634)
);

AO221x2_ASAP7_75t_L g1635 ( 
.A1(n_1570),
.A2(n_1542),
.B1(n_1442),
.B2(n_1581),
.C(n_1572),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1500),
.A2(n_1470),
.B1(n_1546),
.B2(n_1556),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1554),
.B(n_1564),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1558),
.B(n_1493),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1546),
.A2(n_1559),
.B1(n_1573),
.B2(n_1558),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1493),
.B(n_1547),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1545),
.B2(n_1547),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1545),
.A2(n_1561),
.B1(n_1565),
.B2(n_1586),
.C(n_1582),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1561),
.A2(n_1577),
.B1(n_1565),
.B2(n_1576),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1526),
.A2(n_1584),
.B1(n_1583),
.B2(n_1579),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1442),
.A2(n_1586),
.B1(n_1574),
.B2(n_1585),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1526),
.A2(n_1579),
.B1(n_1575),
.B2(n_1574),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1577),
.A2(n_1548),
.B1(n_1578),
.B2(n_1585),
.C(n_1571),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1548),
.A2(n_1509),
.B(n_1526),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1509),
.B(n_1555),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1575),
.A2(n_985),
.B1(n_1406),
.B2(n_1457),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1555),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1555),
.B(n_1544),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1481),
.B(n_1503),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1654)
);

CKINVDCx11_ASAP7_75t_R g1655 ( 
.A(n_1486),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1452),
.Y(n_1656)
);

AO21x2_ASAP7_75t_L g1657 ( 
.A1(n_1483),
.A2(n_1485),
.B(n_1548),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1437),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1659)
);

BUFx4f_ASAP7_75t_SL g1660 ( 
.A(n_1486),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_751),
.B2(n_1386),
.C(n_591),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1477),
.A2(n_985),
.B1(n_1457),
.B2(n_1194),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1477),
.A2(n_985),
.B1(n_1457),
.B2(n_1194),
.Y(n_1663)
);

AOI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1457),
.A2(n_985),
.B(n_1071),
.Y(n_1664)
);

AND2x4_ASAP7_75t_SL g1665 ( 
.A(n_1486),
.B(n_1393),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1440),
.A2(n_985),
.B1(n_1014),
.B2(n_637),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1437),
.Y(n_1667)
);

OAI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1477),
.A2(n_1435),
.B1(n_985),
.B2(n_1478),
.C1(n_1436),
.C2(n_1408),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1500),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1437),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1671)
);

OAI21xp33_ASAP7_75t_L g1672 ( 
.A1(n_1457),
.A2(n_985),
.B(n_751),
.Y(n_1672)
);

AO31x2_ASAP7_75t_L g1673 ( 
.A1(n_1559),
.A2(n_1446),
.A3(n_1570),
.B(n_1483),
.Y(n_1673)
);

OAI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1477),
.A2(n_1408),
.B1(n_502),
.B2(n_985),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_751),
.B2(n_1386),
.C(n_591),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1481),
.B(n_1503),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1677)
);

BUFx8_ASAP7_75t_SL g1678 ( 
.A(n_1452),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1466),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1457),
.B(n_985),
.C(n_1282),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_591),
.B2(n_1386),
.C(n_572),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1386),
.B2(n_1194),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1386),
.B2(n_1194),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1437),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1588),
.B(n_1476),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1466),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1457),
.A2(n_985),
.B(n_1071),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1481),
.B(n_1503),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1485),
.A2(n_1505),
.B(n_1483),
.Y(n_1692)
);

AOI33xp33_ASAP7_75t_L g1693 ( 
.A1(n_1427),
.A2(n_900),
.A3(n_1386),
.B1(n_337),
.B2(n_329),
.B3(n_831),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1477),
.A2(n_985),
.B1(n_1457),
.B2(n_1194),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1588),
.B(n_1476),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_751),
.B2(n_1386),
.C(n_591),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1499),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1499),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1588),
.B(n_1476),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1435),
.A2(n_985),
.B1(n_1014),
.B2(n_1289),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1440),
.A2(n_985),
.B1(n_1014),
.B2(n_637),
.Y(n_1703)
);

AOI222xp33_ASAP7_75t_L g1704 ( 
.A1(n_1457),
.A2(n_1386),
.B1(n_985),
.B2(n_502),
.C1(n_591),
.C2(n_810),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_591),
.B2(n_1386),
.C(n_572),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1437),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_751),
.B2(n_1386),
.C(n_591),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_1406),
.B2(n_1282),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1477),
.A2(n_985),
.B1(n_1457),
.B2(n_1194),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1439),
.A2(n_1071),
.B(n_1310),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1443),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1457),
.A2(n_985),
.B1(n_591),
.B2(n_1386),
.C(n_572),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1477),
.A2(n_985),
.B1(n_1457),
.B2(n_1194),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1466),
.Y(n_1715)
);

INVx4_ASAP7_75t_SL g1716 ( 
.A(n_1508),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1669),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1649),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1634),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1612),
.B(n_1599),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1594),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1711),
.A2(n_1605),
.B(n_1674),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1604),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1658),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1667),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1670),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1635),
.B(n_1652),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1687),
.B(n_1697),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1635),
.B(n_1692),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1635),
.B(n_1652),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1646),
.B(n_1692),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1601),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1626),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1645),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1686),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1648),
.Y(n_1736)
);

INVx4_ASAP7_75t_R g1737 ( 
.A(n_1614),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1646),
.B(n_1644),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1603),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1673),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1673),
.B(n_1657),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1644),
.B(n_1642),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1673),
.B(n_1622),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1603),
.B(n_1707),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1673),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1596),
.B(n_1615),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1704),
.A2(n_1663),
.B1(n_1696),
.B2(n_1714),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1622),
.B(n_1620),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1620),
.B(n_1639),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1639),
.A2(n_1592),
.B(n_1625),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1643),
.B(n_1651),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1689),
.B(n_1680),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1621),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1657),
.B(n_1631),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1597),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1682),
.A2(n_1705),
.B1(n_1713),
.B2(n_1709),
.C1(n_1654),
.C2(n_1695),
.Y(n_1756)
);

AO21x2_ASAP7_75t_L g1757 ( 
.A1(n_1645),
.A2(n_1610),
.B(n_1647),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1602),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1671),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1631),
.B(n_1641),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1662),
.A2(n_1710),
.B1(n_1654),
.B2(n_1709),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1683),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1706),
.B(n_1602),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1716),
.B(n_1641),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1624),
.B(n_1618),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1653),
.B(n_1676),
.Y(n_1766)
);

AOI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1659),
.A2(n_1677),
.B1(n_1681),
.B2(n_1691),
.C1(n_1695),
.C2(n_1694),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1668),
.A2(n_1600),
.B(n_1664),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1600),
.B(n_1636),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1611),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1633),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1633),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1690),
.B(n_1608),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1589),
.B(n_1606),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1595),
.B(n_1623),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1616),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1630),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1632),
.B(n_1636),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_1715),
.Y(n_1779)
);

OAI321xp33_ASAP7_75t_L g1780 ( 
.A1(n_1659),
.A2(n_1677),
.A3(n_1694),
.B1(n_1691),
.B2(n_1681),
.C(n_1590),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1593),
.B(n_1628),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1593),
.B(n_1629),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1780),
.B(n_1661),
.C(n_1675),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1733),
.B(n_1606),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1720),
.B(n_1590),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1727),
.B(n_1730),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1747),
.A2(n_1685),
.B1(n_1684),
.B2(n_1672),
.Y(n_1787)
);

OAI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1747),
.A2(n_1756),
.B(n_1761),
.C(n_1767),
.Y(n_1788)
);

NOR4xp25_ASAP7_75t_L g1789 ( 
.A(n_1780),
.B(n_1708),
.C(n_1698),
.D(n_1650),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1720),
.B(n_1591),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1718),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_L g1792 ( 
.A(n_1756),
.B(n_1650),
.C(n_1666),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1767),
.A2(n_1702),
.B1(n_1703),
.B2(n_1598),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1724),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1722),
.A2(n_1629),
.B(n_1619),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1725),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1717),
.Y(n_1797)
);

OAI31xp33_ASAP7_75t_L g1798 ( 
.A1(n_1761),
.A2(n_1693),
.A3(n_1665),
.B(n_1627),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1723),
.A2(n_1640),
.B(n_1638),
.Y(n_1799)
);

AOI222xp33_ASAP7_75t_L g1800 ( 
.A1(n_1746),
.A2(n_1660),
.B1(n_1655),
.B2(n_1700),
.C1(n_1699),
.C2(n_1607),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1776),
.A2(n_1699),
.B1(n_1700),
.B2(n_1660),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1688),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1776),
.A2(n_1679),
.B1(n_1613),
.B2(n_1609),
.C(n_1637),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1733),
.A2(n_1617),
.B1(n_1712),
.B2(n_1656),
.C(n_1678),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1779),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1733),
.A2(n_1617),
.B1(n_1712),
.B2(n_1752),
.C(n_1777),
.Y(n_1806)
);

OAI33xp33_ASAP7_75t_L g1807 ( 
.A1(n_1752),
.A2(n_1746),
.A3(n_1777),
.B1(n_1739),
.B2(n_1744),
.B3(n_1735),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1779),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1727),
.B(n_1730),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1774),
.A2(n_1719),
.B1(n_1775),
.B2(n_1765),
.Y(n_1810)
);

OAI31xp33_ASAP7_75t_L g1811 ( 
.A1(n_1765),
.A2(n_1722),
.A3(n_1775),
.B(n_1782),
.Y(n_1811)
);

AOI33xp33_ASAP7_75t_L g1812 ( 
.A1(n_1751),
.A2(n_1742),
.A3(n_1748),
.B1(n_1773),
.B2(n_1749),
.B3(n_1743),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1742),
.A2(n_1751),
.B1(n_1748),
.B2(n_1749),
.C(n_1734),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1774),
.A2(n_1750),
.B(n_1765),
.C(n_1742),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1751),
.A2(n_1748),
.B1(n_1749),
.B2(n_1734),
.C(n_1739),
.Y(n_1815)
);

OAI31xp33_ASAP7_75t_L g1816 ( 
.A1(n_1775),
.A2(n_1782),
.A3(n_1719),
.B(n_1760),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1770),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1727),
.B(n_1730),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1762),
.B(n_1755),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1820)
);

AOI222xp33_ASAP7_75t_L g1821 ( 
.A1(n_1782),
.A2(n_1760),
.B1(n_1719),
.B2(n_1758),
.C1(n_1759),
.C2(n_1773),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1760),
.A2(n_1743),
.B1(n_1719),
.B2(n_1771),
.C(n_1772),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1721),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1762),
.B(n_1718),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1750),
.A2(n_1732),
.B1(n_1758),
.B2(n_1769),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1721),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1728),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1750),
.A2(n_1729),
.B(n_1743),
.C(n_1736),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1759),
.B(n_1728),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1729),
.B(n_1718),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1771),
.A2(n_1772),
.B1(n_1744),
.B2(n_1758),
.C(n_1773),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1738),
.B(n_1729),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1738),
.B(n_1731),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1732),
.A2(n_1764),
.B(n_1769),
.C(n_1736),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1726),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1731),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1830),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1833),
.B(n_1731),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1832),
.B(n_1820),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1819),
.Y(n_1840)
);

OAI31xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1788),
.A2(n_1764),
.A3(n_1778),
.B(n_1781),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1807),
.B(n_1792),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1832),
.B(n_1736),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1794),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1819),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1809),
.B(n_1818),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1830),
.Y(n_1847)
);

NAND2x1_ASAP7_75t_SL g1848 ( 
.A(n_1784),
.B(n_1740),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1809),
.B(n_1754),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1796),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1818),
.B(n_1754),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1799),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1827),
.B(n_1753),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1791),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1786),
.B(n_1824),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1786),
.B(n_1745),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1797),
.B(n_1741),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1829),
.B(n_1735),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1717),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1828),
.B(n_1741),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1823),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1799),
.B(n_1723),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1826),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1805),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1855),
.B(n_1808),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1840),
.B(n_1802),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1864),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1863),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1842),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1855),
.B(n_1817),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1836),
.B(n_1812),
.Y(n_1872)
);

NAND4xp25_ASAP7_75t_L g1873 ( 
.A(n_1842),
.B(n_1792),
.C(n_1787),
.D(n_1810),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1864),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1836),
.B(n_1817),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1836),
.B(n_1757),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1861),
.A2(n_1814),
.B(n_1750),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1862),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1862),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1861),
.A2(n_1750),
.B1(n_1825),
.B2(n_1784),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1844),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1848),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1854),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1838),
.B(n_1822),
.Y(n_1885)
);

NOR2xp67_ASAP7_75t_L g1886 ( 
.A(n_1861),
.B(n_1835),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1844),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1838),
.B(n_1831),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1859),
.B(n_1790),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1841),
.A2(n_1793),
.B1(n_1783),
.B2(n_1813),
.Y(n_1890)
);

OAI31xp33_ASAP7_75t_L g1891 ( 
.A1(n_1843),
.A2(n_1811),
.A3(n_1816),
.B(n_1798),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1860),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1850),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1838),
.B(n_1757),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1859),
.B(n_1815),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1850),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1845),
.B(n_1763),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1845),
.B(n_1763),
.Y(n_1898)
);

CKINVDCx16_ASAP7_75t_R g1899 ( 
.A(n_1890),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1879),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1870),
.B(n_1843),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1870),
.B(n_1843),
.Y(n_1902)
);

AND2x2_ASAP7_75t_SL g1903 ( 
.A(n_1883),
.B(n_1789),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1883),
.B(n_1849),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1882),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1876),
.B(n_1849),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1878),
.B(n_1877),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1876),
.B(n_1894),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1882),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1879),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1872),
.B(n_1839),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1873),
.B(n_1853),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1887),
.Y(n_1913)
);

NAND3xp33_ASAP7_75t_L g1914 ( 
.A(n_1890),
.B(n_1798),
.C(n_1816),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1872),
.B(n_1839),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1873),
.B(n_1806),
.C(n_1785),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1887),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1868),
.B(n_1858),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1894),
.B(n_1849),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1895),
.B(n_1839),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1893),
.Y(n_1923)
);

INVxp67_ASAP7_75t_SL g1924 ( 
.A(n_1884),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1869),
.B(n_1851),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1884),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1895),
.B(n_1853),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1879),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_L g1929 ( 
.A(n_1878),
.B(n_1852),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1869),
.B(n_1875),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1869),
.B(n_1857),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1880),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1889),
.B(n_1847),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1875),
.B(n_1857),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1880),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1874),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1880),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1871),
.B(n_1857),
.Y(n_1938)
);

NAND2x1_ASAP7_75t_L g1939 ( 
.A(n_1868),
.B(n_1837),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1865),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1888),
.B(n_1892),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1885),
.B(n_1766),
.Y(n_1942)
);

AND5x1_ASAP7_75t_L g1943 ( 
.A(n_1891),
.B(n_1804),
.C(n_1803),
.D(n_1834),
.E(n_1848),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1926),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1926),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1903),
.B(n_1885),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1903),
.B(n_1888),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1907),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1924),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1846),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1939),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1903),
.B(n_1891),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1899),
.B(n_1865),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1914),
.A2(n_1881),
.B(n_1821),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1905),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1903),
.B(n_1866),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1904),
.B(n_1846),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1916),
.B(n_1866),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1899),
.A2(n_1757),
.B1(n_1768),
.B2(n_1795),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1905),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1914),
.A2(n_1874),
.B(n_1892),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1916),
.B(n_1897),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1909),
.Y(n_1963)
);

AOI21xp33_ASAP7_75t_L g1964 ( 
.A1(n_1912),
.A2(n_1800),
.B(n_1852),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1909),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1913),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1904),
.B(n_1846),
.Y(n_1967)
);

NOR4xp25_ASAP7_75t_L g1968 ( 
.A(n_1912),
.B(n_1898),
.C(n_1897),
.D(n_1867),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1904),
.B(n_1871),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_SL g1970 ( 
.A1(n_1929),
.A2(n_1801),
.B(n_1764),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1929),
.A2(n_1848),
.B(n_1852),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1942),
.B(n_1927),
.Y(n_1972)
);

AND2x2_ASAP7_75t_SL g1973 ( 
.A(n_1941),
.B(n_1795),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1942),
.B(n_1898),
.Y(n_1974)
);

O2A1O1Ixp33_ASAP7_75t_L g1975 ( 
.A1(n_1941),
.A2(n_1757),
.B(n_1768),
.C(n_1732),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_SL g1976 ( 
.A1(n_1943),
.A2(n_1764),
.B(n_1778),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1938),
.B(n_1856),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1924),
.Y(n_1978)
);

NAND2x1_ASAP7_75t_L g1979 ( 
.A(n_1920),
.B(n_1737),
.Y(n_1979)
);

OAI21xp33_ASAP7_75t_L g1980 ( 
.A1(n_1927),
.A2(n_1732),
.B(n_1769),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1954),
.A2(n_1936),
.B(n_1901),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1944),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1953),
.B(n_1901),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1947),
.B(n_1946),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1949),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1952),
.A2(n_1757),
.B1(n_1921),
.B2(n_1768),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1948),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1945),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1976),
.B(n_1902),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1976),
.A2(n_1902),
.B1(n_1940),
.B2(n_1921),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1956),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1968),
.B(n_1911),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1958),
.B(n_1933),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1945),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_L g1995 ( 
.A(n_1964),
.B(n_1936),
.C(n_1939),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1978),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1955),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1972),
.B(n_1933),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1973),
.A2(n_1768),
.B1(n_1915),
.B2(n_1911),
.Y(n_1999)
);

AOI211xp5_ASAP7_75t_SL g2000 ( 
.A1(n_1961),
.A2(n_1943),
.B(n_1915),
.C(n_1922),
.Y(n_2000)
);

AOI31xp33_ASAP7_75t_L g2001 ( 
.A1(n_1962),
.A2(n_1943),
.A3(n_1922),
.B(n_1920),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1980),
.B(n_1934),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1955),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1960),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1950),
.B(n_1938),
.Y(n_2005)
);

NAND4xp25_ASAP7_75t_SL g2006 ( 
.A(n_1975),
.B(n_1959),
.C(n_1950),
.D(n_1971),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1980),
.B(n_1867),
.Y(n_2007)
);

NOR2x1_ASAP7_75t_L g2008 ( 
.A(n_2006),
.B(n_1951),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1985),
.B(n_1974),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1987),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1987),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_SL g2012 ( 
.A(n_1984),
.B(n_1970),
.C(n_1963),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1991),
.B(n_1973),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1992),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_2005),
.B(n_1969),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1995),
.B(n_1973),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2003),
.Y(n_2017)
);

XNOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_1990),
.B(n_1959),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1985),
.B(n_1957),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2003),
.Y(n_2020)
);

XNOR2x1_ASAP7_75t_L g2021 ( 
.A(n_1992),
.B(n_1979),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2004),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2005),
.B(n_1969),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1988),
.B(n_1994),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2004),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1996),
.B(n_1957),
.Y(n_2026)
);

INVxp33_ASAP7_75t_SL g2027 ( 
.A(n_1982),
.Y(n_2027)
);

NAND2xp33_ASAP7_75t_L g2028 ( 
.A(n_2012),
.B(n_1983),
.Y(n_2028)
);

NAND2x1_ASAP7_75t_L g2029 ( 
.A(n_2015),
.B(n_1951),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_SL g2030 ( 
.A(n_2014),
.B(n_2000),
.C(n_1981),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2008),
.A2(n_1970),
.B1(n_2007),
.B2(n_1989),
.Y(n_2031)
);

NOR3xp33_ASAP7_75t_L g2032 ( 
.A(n_2010),
.B(n_1993),
.C(n_2001),
.Y(n_2032)
);

NOR2x1_ASAP7_75t_L g2033 ( 
.A(n_2011),
.B(n_1997),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_2016),
.A2(n_1999),
.B1(n_1986),
.B2(n_1998),
.C(n_2002),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2024),
.B(n_1967),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2024),
.B(n_1967),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2019),
.Y(n_2037)
);

NAND4xp25_ASAP7_75t_L g2038 ( 
.A(n_2027),
.B(n_1963),
.C(n_1960),
.D(n_1965),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_2016),
.A2(n_1979),
.B(n_1966),
.C(n_1965),
.Y(n_2039)
);

NAND4xp25_ASAP7_75t_L g2040 ( 
.A(n_2027),
.B(n_1966),
.C(n_1977),
.D(n_1920),
.Y(n_2040)
);

NAND3xp33_ASAP7_75t_L g2041 ( 
.A(n_2033),
.B(n_2021),
.C(n_2018),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_2028),
.A2(n_2021),
.B(n_2013),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2030),
.A2(n_2026),
.B(n_2009),
.Y(n_2043)
);

AOI322xp5_ASAP7_75t_L g2044 ( 
.A1(n_2032),
.A2(n_2015),
.A3(n_2023),
.B1(n_2022),
.B2(n_2020),
.C1(n_2017),
.C2(n_2025),
.Y(n_2044)
);

XOR2xp5_ASAP7_75t_L g2045 ( 
.A(n_2031),
.B(n_2009),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2039),
.A2(n_2019),
.B(n_2023),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2037),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2034),
.A2(n_1922),
.B1(n_1930),
.B2(n_1977),
.Y(n_2048)
);

AOI211x1_ASAP7_75t_L g2049 ( 
.A1(n_2040),
.A2(n_1930),
.B(n_1913),
.C(n_1917),
.Y(n_2049)
);

O2A1O1Ixp33_ASAP7_75t_L g2050 ( 
.A1(n_2038),
.A2(n_1918),
.B(n_1923),
.C(n_1917),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2047),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2049),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_2035),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_2041),
.A2(n_2036),
.B1(n_2029),
.B2(n_1918),
.Y(n_2054)
);

AND2x2_ASAP7_75t_SL g2055 ( 
.A(n_2045),
.B(n_1930),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2050),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2055),
.A2(n_2042),
.B1(n_2043),
.B2(n_2056),
.Y(n_2057)
);

NOR3x1_ASAP7_75t_L g2058 ( 
.A(n_2054),
.B(n_2048),
.C(n_2044),
.Y(n_2058)
);

NOR3xp33_ASAP7_75t_L g2059 ( 
.A(n_2053),
.B(n_1910),
.C(n_1937),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2055),
.B(n_1934),
.Y(n_2060)
);

NOR2x1p5_ASAP7_75t_L g2061 ( 
.A(n_2052),
.B(n_1918),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2053),
.B(n_2052),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2051),
.A2(n_1925),
.B1(n_1923),
.B2(n_1931),
.Y(n_2063)
);

NOR4xp25_ASAP7_75t_L g2064 ( 
.A(n_2057),
.B(n_1900),
.C(n_1937),
.D(n_1935),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2060),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_2061),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_2062),
.B(n_1910),
.C(n_1937),
.Y(n_2067)
);

NAND4xp25_ASAP7_75t_L g2068 ( 
.A(n_2058),
.B(n_1908),
.C(n_1925),
.D(n_1931),
.Y(n_2068)
);

A2O1A1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_2059),
.A2(n_1925),
.B(n_1935),
.C(n_1900),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_2066),
.A2(n_2063),
.B(n_1900),
.C(n_1935),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_2065),
.Y(n_2071)
);

OR2x6_ASAP7_75t_L g2072 ( 
.A(n_2064),
.B(n_1770),
.Y(n_2072)
);

NAND4xp25_ASAP7_75t_L g2073 ( 
.A(n_2068),
.B(n_2067),
.C(n_2069),
.D(n_1908),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_2072),
.Y(n_2074)
);

OAI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_2074),
.A2(n_2071),
.B(n_2073),
.C(n_2070),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2075),
.B(n_1908),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2075),
.Y(n_2077)
);

OAI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2076),
.A2(n_1928),
.B(n_1932),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2077),
.Y(n_2079)
);

BUFx2_ASAP7_75t_L g2080 ( 
.A(n_2079),
.Y(n_2080)
);

AOI221xp5_ASAP7_75t_L g2081 ( 
.A1(n_2078),
.A2(n_1932),
.B1(n_1928),
.B2(n_1910),
.C(n_1931),
.Y(n_2081)
);

AOI322xp5_ASAP7_75t_L g2082 ( 
.A1(n_2080),
.A2(n_1932),
.A3(n_1928),
.B1(n_1910),
.B2(n_1919),
.C1(n_1906),
.C2(n_1938),
.Y(n_2082)
);

AOI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2082),
.A2(n_2081),
.B1(n_1910),
.B2(n_1896),
.C(n_1893),
.Y(n_2083)
);

AOI211xp5_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_1919),
.B(n_1906),
.C(n_1896),
.Y(n_2084)
);


endmodule