module fake_jpeg_4002_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_16),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_24),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_18),
.B(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_52),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_33),
.B1(n_29),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_56),
.B1(n_61),
.B2(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_25),
.B1(n_21),
.B2(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_33),
.B1(n_17),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_47),
.B1(n_22),
.B2(n_19),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_75),
.B(n_99),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_41),
.C(n_37),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_32),
.C(n_24),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_62),
.B1(n_47),
.B2(n_19),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_20),
.B1(n_39),
.B2(n_40),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_44),
.B1(n_39),
.B2(n_40),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_57),
.B1(n_26),
.B2(n_23),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_44),
.B1(n_39),
.B2(n_20),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_98),
.B1(n_68),
.B2(n_32),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_55),
.B(n_36),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_46),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_17),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_39),
.B1(n_26),
.B2(n_23),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_68),
.B1(n_36),
.B2(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_107),
.B1(n_112),
.B2(n_116),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_36),
.B1(n_38),
.B2(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_38),
.B1(n_36),
.B2(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_30),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_125),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_77),
.B1(n_75),
.B2(n_71),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_24),
.B1(n_28),
.B2(n_32),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_28),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_94),
.B1(n_92),
.B2(n_82),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_92),
.B(n_84),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_144),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_143),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_76),
.B(n_80),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_91),
.B(n_38),
.C(n_46),
.D(n_35),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_35),
.B(n_27),
.C(n_46),
.D(n_64),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_95),
.B(n_46),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_80),
.B1(n_84),
.B2(n_89),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_108),
.B1(n_90),
.B2(n_101),
.Y(n_171)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_106),
.B1(n_122),
.B2(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_123),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_174),
.A3(n_183),
.B1(n_139),
.B2(n_154),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_190),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_142),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_165),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_115),
.A3(n_127),
.B1(n_114),
.B2(n_116),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_110),
.C(n_124),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_178),
.C(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_104),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_14),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_191),
.B1(n_141),
.B2(n_147),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_30),
.B(n_34),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_153),
.B(n_130),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_140),
.B1(n_158),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_184),
.B1(n_192),
.B2(n_159),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_95),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_95),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_72),
.B1(n_87),
.B2(n_74),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_109),
.C(n_101),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_73),
.B1(n_100),
.B2(n_49),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_143),
.B1(n_138),
.B2(n_156),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_88),
.B(n_35),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_59),
.B1(n_52),
.B2(n_88),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_109),
.C(n_83),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_145),
.C(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_200),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_205),
.C(n_223),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_210),
.B1(n_208),
.B2(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_155),
.C(n_143),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_208),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_35),
.B1(n_27),
.B2(n_83),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_209),
.B1(n_214),
.B2(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_27),
.B1(n_15),
.B2(n_14),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_15),
.Y(n_211)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_162),
.B1(n_182),
.B2(n_189),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_215),
.B(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_3),
.B(n_4),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_3),
.B(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_170),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_236),
.Y(n_253)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_221),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_178),
.B1(n_185),
.B2(n_193),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_235),
.B1(n_199),
.B2(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_174),
.B1(n_169),
.B2(n_190),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_164),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_190),
.B1(n_175),
.B2(n_168),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_230),
.B1(n_225),
.B2(n_246),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_167),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_243),
.C(n_247),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_213),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_13),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_3),
.C(n_5),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_252),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_222),
.B(n_217),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_257),
.B(n_258),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_249),
.A2(n_219),
.B1(n_196),
.B2(n_197),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_249),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_215),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_264),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_207),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_206),
.C(n_209),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_231),
.C(n_234),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_12),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_5),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_12),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.C(n_285),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_238),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_251),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_258),
.A2(n_235),
.B1(n_229),
.B2(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_247),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_254),
.B(n_243),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_231),
.C(n_7),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_6),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_7),
.C(n_8),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_283),
.A2(n_255),
.B1(n_266),
.B2(n_260),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_292),
.B1(n_280),
.B2(n_278),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_259),
.B(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_256),
.B(n_7),
.Y(n_293)
);

NAND4xp25_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_6),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_276),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_305),
.B(n_314),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_277),
.B1(n_275),
.B2(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_287),
.B(n_274),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_313),
.B(n_295),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_290),
.B1(n_293),
.B2(n_294),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_294),
.B(n_274),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_317),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_289),
.C(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_322),
.Y(n_329)
);

INVx11_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_290),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_314),
.B(n_303),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_289),
.B(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_300),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_292),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_326),
.B(n_328),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_327),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_296),
.B(n_310),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_318),
.C(n_321),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_332),
.B(n_324),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_330),
.B(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_320),
.C(n_316),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_8),
.A3(n_9),
.B1(n_324),
.B2(n_326),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_8),
.Y(n_338)
);


endmodule