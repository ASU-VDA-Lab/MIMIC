module real_aes_11997_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_1840;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1800;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1802;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1280;
wire n_729;
wire n_394;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1410 ( .A1(n_0), .A2(n_410), .B1(n_1016), .B2(n_1411), .C(n_1416), .Y(n_1410) );
AOI21xp33_ASAP7_75t_L g1438 ( .A1(n_0), .A2(n_630), .B(n_1194), .Y(n_1438) );
INVxp67_ASAP7_75t_L g418 ( .A(n_1), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_1), .A2(n_189), .B1(n_480), .B2(n_509), .C(n_514), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_2), .A2(n_935), .B1(n_937), .B2(n_943), .C(n_949), .Y(n_934) );
INVx1_ASAP7_75t_L g973 ( .A(n_2), .Y(n_973) );
INVx1_ASAP7_75t_L g1339 ( .A(n_3), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_4), .Y(n_1271) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_5), .A2(n_239), .B1(n_360), .B2(n_371), .C(n_378), .Y(n_359) );
INVx1_ASAP7_75t_L g495 ( .A(n_5), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_6), .A2(n_96), .B1(n_374), .B2(n_926), .C(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g988 ( .A(n_6), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g1419 ( .A1(n_7), .A2(n_179), .B1(n_395), .B2(n_404), .C(n_407), .Y(n_1419) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_7), .Y(n_1443) );
AO22x1_ASAP7_75t_L g909 ( .A1(n_8), .A2(n_910), .B1(n_994), .B2(n_995), .Y(n_909) );
INVx1_ASAP7_75t_L g995 ( .A(n_8), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g1810 ( .A1(n_9), .A2(n_304), .B1(n_924), .B2(n_1379), .C(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1818 ( .A(n_9), .Y(n_1818) );
INVx1_ASAP7_75t_L g1151 ( .A(n_10), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_11), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_12), .A2(n_293), .B1(n_1085), .B2(n_1087), .Y(n_1084) );
INVx1_ASAP7_75t_L g1116 ( .A(n_12), .Y(n_1116) );
INVx1_ASAP7_75t_L g1796 ( .A(n_13), .Y(n_1796) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_14), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g1462 ( .A1(n_15), .A2(n_147), .B1(n_597), .B2(n_598), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_15), .A2(n_235), .B1(n_1196), .B2(n_1481), .C(n_1483), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_16), .A2(n_153), .B1(n_798), .B2(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g830 ( .A(n_16), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_17), .A2(n_104), .B1(n_393), .B2(n_402), .C(n_407), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_17), .A2(n_104), .B1(n_463), .B2(n_474), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g1045 ( .A1(n_18), .A2(n_70), .B1(n_474), .B2(n_1046), .C(n_1047), .Y(n_1045) );
INVx1_ASAP7_75t_L g1050 ( .A(n_18), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1318 ( .A(n_19), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_20), .A2(n_192), .B1(n_481), .B2(n_1082), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_20), .A2(n_192), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
AO221x2_ASAP7_75t_L g1572 ( .A1(n_21), .A2(n_254), .B1(n_1549), .B2(n_1571), .C(n_1573), .Y(n_1572) );
CKINVDCx16_ASAP7_75t_R g1593 ( .A(n_22), .Y(n_1593) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_23), .A2(n_212), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_23), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1798 ( .A1(n_24), .A2(n_41), .B1(n_1336), .B2(n_1799), .C(n_1800), .Y(n_1798) );
AOI22xp33_ASAP7_75t_L g1823 ( .A1(n_24), .A2(n_277), .B1(n_1824), .B2(n_1825), .Y(n_1823) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_25), .Y(n_1414) );
INVx1_ASAP7_75t_L g1802 ( .A(n_26), .Y(n_1802) );
AOI221xp5_ASAP7_75t_L g1820 ( .A1(n_26), .A2(n_41), .B1(n_1509), .B2(n_1821), .C(n_1822), .Y(n_1820) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_27), .A2(n_311), .B1(n_592), .B2(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g636 ( .A(n_27), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g1421 ( .A1(n_28), .A2(n_67), .B1(n_903), .B2(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1436 ( .A(n_28), .Y(n_1436) );
INVxp33_ASAP7_75t_L g1249 ( .A(n_29), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_29), .A2(n_86), .B1(n_1277), .B2(n_1278), .C(n_1280), .Y(n_1276) );
INVx1_ASAP7_75t_L g1813 ( .A(n_30), .Y(n_1813) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_31), .A2(n_226), .B1(n_515), .B2(n_647), .C(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g693 ( .A(n_31), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g1258 ( .A1(n_32), .A2(n_163), .B1(n_1259), .B2(n_1261), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_32), .A2(n_163), .B1(n_1291), .B2(n_1293), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_33), .A2(n_118), .B1(n_598), .B2(n_1108), .C(n_1110), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_33), .A2(n_151), .B1(n_1120), .B2(n_1122), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_34), .A2(n_38), .B1(n_746), .B2(n_924), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_34), .A2(n_96), .B1(n_990), .B2(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g335 ( .A(n_35), .Y(n_335) );
INVx1_ASAP7_75t_L g734 ( .A(n_36), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_36), .A2(n_267), .B1(n_777), .B2(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g1367 ( .A(n_37), .Y(n_1367) );
OAI221xp5_ASAP7_75t_L g1390 ( .A1(n_37), .A2(n_935), .B1(n_1102), .B2(n_1391), .C(n_1394), .Y(n_1390) );
INVx1_ASAP7_75t_L g986 ( .A(n_38), .Y(n_986) );
INVx1_ASAP7_75t_L g721 ( .A(n_39), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_40), .A2(n_102), .B1(n_582), .B2(n_585), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_40), .A2(n_203), .B1(n_628), .B2(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g1377 ( .A(n_42), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_42), .A2(n_223), .B1(n_1120), .B2(n_1122), .Y(n_1404) );
AOI22xp33_ASAP7_75t_SL g1263 ( .A1(n_43), .A2(n_288), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1285 ( .A1(n_43), .A2(n_288), .B1(n_660), .B2(n_1286), .C(n_1288), .Y(n_1285) );
INVx1_ASAP7_75t_L g601 ( .A(n_44), .Y(n_601) );
INVxp33_ASAP7_75t_L g724 ( .A(n_45), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_45), .A2(n_282), .B1(n_650), .B2(n_765), .C(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g1080 ( .A(n_46), .Y(n_1080) );
OAI211xp5_ASAP7_75t_SL g1103 ( .A1(n_46), .A2(n_913), .B(n_1104), .C(n_1111), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_47), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g1468 ( .A(n_48), .Y(n_1468) );
INVx1_ASAP7_75t_L g855 ( .A(n_49), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_49), .A2(n_274), .B1(n_882), .B2(n_883), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_50), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_51), .A2(n_93), .B1(n_929), .B2(n_933), .Y(n_928) );
OAI22xp5_ASAP7_75t_SL g958 ( .A1(n_51), .A2(n_93), .B1(n_959), .B2(n_963), .Y(n_958) );
XOR2x2_ASAP7_75t_L g1449 ( .A(n_52), .B(n_1450), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_53), .A2(n_327), .B1(n_518), .B2(n_1311), .Y(n_1313) );
OAI22xp33_ASAP7_75t_L g1347 ( .A1(n_53), .A2(n_307), .B1(n_935), .B2(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1175 ( .A(n_54), .Y(n_1175) );
OAI221xp5_ASAP7_75t_L g1180 ( .A1(n_54), .A2(n_270), .B1(n_1181), .B2(n_1182), .C(n_1184), .Y(n_1180) );
AOI22xp33_ASAP7_75t_SL g1266 ( .A1(n_55), .A2(n_122), .B1(n_1261), .B2(n_1264), .Y(n_1266) );
INVxp67_ASAP7_75t_SL g1274 ( .A(n_55), .Y(n_1274) );
INVx1_ASAP7_75t_L g753 ( .A(n_56), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g1459 ( .A(n_57), .Y(n_1459) );
AOI22xp5_ASAP7_75t_L g1599 ( .A1(n_58), .A2(n_303), .B1(n_1549), .B2(n_1571), .Y(n_1599) );
INVx1_ASAP7_75t_L g1795 ( .A(n_59), .Y(n_1795) );
INVxp33_ASAP7_75t_SL g1460 ( .A(n_60), .Y(n_1460) );
AOI221xp5_ASAP7_75t_L g1474 ( .A1(n_60), .A2(n_229), .B1(n_613), .B2(n_1475), .C(n_1477), .Y(n_1474) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_61), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_62), .A2(n_172), .B1(n_956), .B2(n_1385), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_62), .A2(n_172), .B1(n_533), .B2(n_792), .Y(n_1426) );
OAI22xp33_ASAP7_75t_L g1199 ( .A1(n_63), .A2(n_306), .B1(n_474), .B2(n_1200), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_63), .A2(n_306), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_1223) );
INVx1_ASAP7_75t_L g751 ( .A(n_64), .Y(n_751) );
INVx1_ASAP7_75t_L g951 ( .A(n_65), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g1463 ( .A1(n_66), .A2(n_235), .B1(n_1264), .B2(n_1464), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_66), .A2(n_147), .B1(n_633), .B2(n_1486), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_67), .A2(n_112), .B1(n_456), .B2(n_1434), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_68), .A2(n_292), .B1(n_545), .B2(n_902), .Y(n_1022) );
INVx1_ASAP7_75t_L g1048 ( .A(n_68), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1454 ( .A(n_69), .Y(n_1454) );
OAI22xp33_ASAP7_75t_L g1472 ( .A1(n_69), .A2(n_276), .B1(n_606), .B2(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1051 ( .A(n_70), .Y(n_1051) );
INVx1_ASAP7_75t_L g1212 ( .A(n_71), .Y(n_1212) );
XOR2xp5_ASAP7_75t_L g1302 ( .A(n_72), .B(n_1303), .Y(n_1302) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_73), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g1267 ( .A1(n_74), .A2(n_108), .B1(n_1259), .B2(n_1265), .Y(n_1267) );
INVxp67_ASAP7_75t_L g1284 ( .A(n_74), .Y(n_1284) );
INVx1_ASAP7_75t_L g1337 ( .A(n_75), .Y(n_1337) );
INVx1_ASAP7_75t_L g1457 ( .A(n_76), .Y(n_1457) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_77), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_78), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_79), .A2(n_289), .B1(n_1308), .B2(n_1309), .Y(n_1307) );
INVx1_ASAP7_75t_L g1326 ( .A(n_79), .Y(n_1326) );
INVx1_ASAP7_75t_L g560 ( .A(n_80), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_80), .A2(n_161), .B1(n_606), .B2(n_607), .Y(n_605) );
OAI222xp33_ASAP7_75t_L g1134 ( .A1(n_81), .A2(n_137), .B1(n_285), .B2(n_545), .C1(n_728), .C2(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1161 ( .A(n_81), .Y(n_1161) );
OAI211xp5_ASAP7_75t_SL g865 ( .A1(n_82), .A2(n_866), .B(n_867), .C(n_870), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_82), .A2(n_184), .B1(n_886), .B2(n_890), .Y(n_889) );
AOI221xp5_ASAP7_75t_L g1500 ( .A1(n_83), .A2(n_220), .B1(n_650), .B2(n_1501), .C(n_1502), .Y(n_1500) );
INVx1_ASAP7_75t_L g1520 ( .A(n_83), .Y(n_1520) );
INVx1_ASAP7_75t_L g756 ( .A(n_84), .Y(n_756) );
AO22x2_ASAP7_75t_L g996 ( .A1(n_85), .A2(n_997), .B1(n_1052), .B2(n_1053), .Y(n_996) );
CKINVDCx14_ASAP7_75t_R g1052 ( .A(n_85), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g1253 ( .A(n_86), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_87), .A2(n_320), .B1(n_656), .B2(n_810), .Y(n_809) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_87), .A2(n_320), .B1(n_393), .B2(n_403), .C(n_681), .Y(n_825) );
INVx1_ASAP7_75t_L g368 ( .A(n_88), .Y(n_368) );
OR2x2_ASAP7_75t_L g400 ( .A(n_88), .B(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g413 ( .A(n_88), .Y(n_413) );
BUFx2_ASAP7_75t_L g548 ( .A(n_88), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g1415 ( .A1(n_89), .A2(n_134), .B1(n_956), .B2(n_1385), .Y(n_1415) );
INVx1_ASAP7_75t_L g1432 ( .A(n_89), .Y(n_1432) );
INVx1_ASAP7_75t_L g1363 ( .A(n_90), .Y(n_1363) );
INVx1_ASAP7_75t_L g757 ( .A(n_91), .Y(n_757) );
INVx1_ASAP7_75t_L g942 ( .A(n_92), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_92), .A2(n_214), .B1(n_614), .B2(n_863), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_94), .Y(n_1198) );
AOI22xp33_ASAP7_75t_SL g1465 ( .A1(n_95), .A2(n_197), .B1(n_1264), .B2(n_1464), .Y(n_1465) );
INVxp33_ASAP7_75t_SL g1489 ( .A(n_95), .Y(n_1489) );
INVx1_ASAP7_75t_L g920 ( .A(n_97), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_97), .A2(n_248), .B1(n_455), .B2(n_614), .Y(n_975) );
CKINVDCx5p33_ASAP7_75t_R g1504 ( .A(n_98), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1400 ( .A(n_99), .Y(n_1400) );
INVx1_ASAP7_75t_L g723 ( .A(n_100), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_101), .A2(n_312), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_101), .A2(n_312), .B1(n_474), .B2(n_763), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_102), .A2(n_263), .B1(n_515), .B2(n_623), .C(n_625), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_103), .A2(n_186), .B1(n_647), .B2(n_767), .C(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_103), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g1466 ( .A1(n_105), .A2(n_246), .B1(n_597), .B2(n_598), .Y(n_1466) );
INVxp33_ASAP7_75t_L g1488 ( .A(n_105), .Y(n_1488) );
INVx1_ASAP7_75t_L g574 ( .A(n_106), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_106), .A2(n_114), .B1(n_610), .B2(n_613), .C(n_615), .Y(n_609) );
CKINVDCx16_ASAP7_75t_R g1595 ( .A(n_107), .Y(n_1595) );
INVxp33_ASAP7_75t_L g1295 ( .A(n_108), .Y(n_1295) );
INVx1_ASAP7_75t_L g1077 ( .A(n_109), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_109), .A2(n_935), .B1(n_1093), .B2(n_1096), .C(n_1102), .Y(n_1092) );
INVx1_ASAP7_75t_L g1812 ( .A(n_110), .Y(n_1812) );
OAI221xp5_ASAP7_75t_L g1816 ( .A1(n_110), .A2(n_304), .B1(n_808), .B2(n_1164), .C(n_1817), .Y(n_1816) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_111), .A2(n_125), .B1(n_650), .B2(n_1370), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_111), .A2(n_125), .B1(n_1323), .B2(n_1348), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_112), .A2(n_131), .B1(n_545), .B2(n_902), .Y(n_1423) );
INVx1_ASAP7_75t_L g552 ( .A(n_113), .Y(n_552) );
INVx1_ASAP7_75t_L g569 ( .A(n_114), .Y(n_569) );
INVx1_ASAP7_75t_L g1252 ( .A(n_115), .Y(n_1252) );
INVx1_ASAP7_75t_L g379 ( .A(n_116), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_117), .A2(n_155), .B1(n_519), .B2(n_647), .C(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g822 ( .A(n_117), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_118), .A2(n_195), .B1(n_990), .B2(n_992), .Y(n_1118) );
INVxp67_ASAP7_75t_L g743 ( .A(n_119), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_119), .A2(n_199), .B1(n_515), .B2(n_772), .C(n_774), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_120), .Y(n_1512) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_121), .Y(n_668) );
INVxp33_ASAP7_75t_L g1296 ( .A(n_122), .Y(n_1296) );
XOR2x2_ASAP7_75t_L g1355 ( .A(n_123), .B(n_1356), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1570 ( .A1(n_124), .A2(n_298), .B1(n_1549), .B2(n_1571), .Y(n_1570) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_126), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_127), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g1507 ( .A1(n_128), .A2(n_242), .B1(n_767), .B2(n_1508), .C(n_1509), .Y(n_1507) );
INVx1_ASAP7_75t_L g1529 ( .A(n_128), .Y(n_1529) );
CKINVDCx5p33_ASAP7_75t_R g1497 ( .A(n_129), .Y(n_1497) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_130), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g1275 ( .A1(n_130), .A2(n_168), .B1(n_463), .B2(n_474), .Y(n_1275) );
INVx1_ASAP7_75t_L g1440 ( .A(n_131), .Y(n_1440) );
INVx1_ASAP7_75t_L g793 ( .A(n_132), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g1492 ( .A(n_133), .B(n_1493), .Y(n_1492) );
AOI22xp5_ASAP7_75t_L g1609 ( .A1(n_133), .A2(n_138), .B1(n_1565), .B2(n_1568), .Y(n_1609) );
INVx1_ASAP7_75t_L g1429 ( .A(n_134), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_135), .Y(n_1058) );
AOI21xp33_ASAP7_75t_L g862 ( .A1(n_136), .A2(n_515), .B(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_136), .A2(n_167), .B1(n_886), .B2(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g1172 ( .A(n_137), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_139), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1610 ( .A1(n_140), .A2(n_310), .B1(n_1543), .B2(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1381 ( .A(n_141), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_141), .A2(n_209), .B1(n_992), .B2(n_1403), .Y(n_1402) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_142), .A2(n_184), .B1(n_533), .B2(n_535), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_142), .A2(n_252), .B1(n_883), .B2(n_894), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_143), .Y(n_662) );
AO221x2_ASAP7_75t_L g1542 ( .A1(n_144), .A2(n_205), .B1(n_1543), .B2(n_1549), .C(n_1550), .Y(n_1542) );
OAI22xp33_ASAP7_75t_SL g1498 ( .A1(n_145), .A2(n_296), .B1(n_1159), .B2(n_1499), .Y(n_1498) );
OAI221xp5_ASAP7_75t_L g1521 ( .A1(n_145), .A2(n_296), .B1(n_393), .B2(n_403), .C(n_1522), .Y(n_1521) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_146), .Y(n_868) );
INVx1_ASAP7_75t_L g1548 ( .A(n_148), .Y(n_1548) );
INVx1_ASAP7_75t_L g1694 ( .A(n_149), .Y(n_1694) );
INVx1_ASAP7_75t_L g1005 ( .A(n_150), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_150), .A2(n_291), .B1(n_614), .B2(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1105 ( .A(n_151), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1598 ( .A1(n_152), .A2(n_317), .B1(n_1565), .B2(n_1568), .Y(n_1598) );
INVx1_ASAP7_75t_L g836 ( .A(n_153), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_154), .A2(n_784), .B1(n_846), .B2(n_847), .Y(n_783) );
INVx1_ASAP7_75t_L g847 ( .A(n_154), .Y(n_847) );
INVx1_ASAP7_75t_L g819 ( .A(n_155), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g1506 ( .A(n_156), .Y(n_1506) );
INVx1_ASAP7_75t_L g1361 ( .A(n_157), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_158), .A2(n_204), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g817 ( .A(n_158), .Y(n_817) );
INVx1_ASAP7_75t_L g1546 ( .A(n_159), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_159), .B(n_1556), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_160), .A2(n_191), .B1(n_612), .B2(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g673 ( .A(n_160), .Y(n_673) );
INVx1_ASAP7_75t_L g565 ( .A(n_161), .Y(n_565) );
INVx1_ASAP7_75t_L g1143 ( .A(n_162), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_164), .Y(n_1503) );
INVx1_ASAP7_75t_L g781 ( .A(n_165), .Y(n_781) );
INVx2_ASAP7_75t_L g347 ( .A(n_166), .Y(n_347) );
INVx1_ASAP7_75t_L g857 ( .A(n_167), .Y(n_857) );
INVxp67_ASAP7_75t_SL g1247 ( .A(n_168), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1145 ( .A(n_169), .Y(n_1145) );
OAI222xp33_ASAP7_75t_L g1163 ( .A1(n_169), .A2(n_176), .B1(n_262), .B2(n_611), .C1(n_1164), .C2(n_1166), .Y(n_1163) );
INVx1_ASAP7_75t_L g1514 ( .A(n_170), .Y(n_1514) );
CKINVDCx5p33_ASAP7_75t_R g1210 ( .A(n_171), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_173), .Y(n_571) );
BUFx3_ASAP7_75t_L g458 ( .A(n_174), .Y(n_458) );
INVx1_ASAP7_75t_L g488 ( .A(n_174), .Y(n_488) );
XNOR2x2_ASAP7_75t_L g356 ( .A(n_175), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g1551 ( .A(n_175), .Y(n_1551) );
INVxp67_ASAP7_75t_L g1150 ( .A(n_176), .Y(n_1150) );
INVxp67_ASAP7_75t_L g432 ( .A(n_177), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_177), .A2(n_244), .B1(n_518), .B2(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g1334 ( .A(n_178), .Y(n_1334) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_179), .Y(n_1444) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_180), .A2(n_280), .B1(n_1192), .B2(n_1193), .C(n_1194), .Y(n_1191) );
INVx1_ASAP7_75t_L g1219 ( .A(n_180), .Y(n_1219) );
INVx1_ASAP7_75t_L g1000 ( .A(n_181), .Y(n_1000) );
AOI21xp33_ASAP7_75t_L g1043 ( .A1(n_181), .A2(n_455), .B(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1692 ( .A(n_182), .Y(n_1692) );
INVx1_ASAP7_75t_L g1803 ( .A(n_183), .Y(n_1803) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_185), .A2(n_305), .B1(n_1278), .B2(n_1365), .Y(n_1364) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_185), .Y(n_1396) );
INVxp67_ASAP7_75t_SL g831 ( .A(n_186), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_187), .A2(n_307), .B1(n_1196), .B2(n_1197), .Y(n_1314) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_187), .A2(n_327), .B1(n_913), .B2(n_1323), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_188), .Y(n_1320) );
INVxp67_ASAP7_75t_L g426 ( .A(n_189), .Y(n_426) );
INVx1_ASAP7_75t_L g1557 ( .A(n_190), .Y(n_1557) );
INVx1_ASAP7_75t_L g677 ( .A(n_191), .Y(n_677) );
INVx1_ASAP7_75t_L g461 ( .A(n_193), .Y(n_461) );
INVx1_ASAP7_75t_L g500 ( .A(n_193), .Y(n_500) );
INVx1_ASAP7_75t_L g789 ( .A(n_194), .Y(n_789) );
INVx1_ASAP7_75t_L g1106 ( .A(n_195), .Y(n_1106) );
INVx1_ASAP7_75t_L g1250 ( .A(n_196), .Y(n_1250) );
INVxp67_ASAP7_75t_SL g1471 ( .A(n_197), .Y(n_1471) );
XNOR2xp5_ASAP7_75t_L g1131 ( .A(n_198), .B(n_1132), .Y(n_1131) );
INVxp67_ASAP7_75t_L g738 ( .A(n_199), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_200), .Y(n_666) );
INVxp67_ASAP7_75t_L g1138 ( .A(n_201), .Y(n_1138) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_201), .A2(n_294), .B1(n_767), .B2(n_795), .C(n_1028), .Y(n_1168) );
INVx1_ASAP7_75t_L g1582 ( .A(n_202), .Y(n_1582) );
OAI21xp33_ASAP7_75t_L g1792 ( .A1(n_202), .A2(n_1793), .B(n_1814), .Y(n_1792) );
INVx1_ASAP7_75t_L g1832 ( .A(n_202), .Y(n_1832) );
AOI22xp5_ASAP7_75t_L g1839 ( .A1(n_202), .A2(n_1840), .B1(n_1845), .B2(n_1849), .Y(n_1839) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_203), .A2(n_263), .B1(n_589), .B2(n_592), .Y(n_588) );
INVx1_ASAP7_75t_L g823 ( .A(n_204), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_206), .Y(n_1008) );
OA22x2_ASAP7_75t_L g639 ( .A1(n_207), .A2(n_640), .B1(n_706), .B2(n_707), .Y(n_639) );
INVx1_ASAP7_75t_L g707 ( .A(n_207), .Y(n_707) );
XOR2xp5_ASAP7_75t_L g1407 ( .A(n_208), .B(n_1408), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_209), .A2(n_223), .B1(n_1383), .B2(n_1384), .C(n_1386), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_210), .A2(n_259), .B1(n_455), .B2(n_614), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_210), .A2(n_323), .B1(n_902), .B2(n_903), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g1564 ( .A1(n_211), .A2(n_271), .B1(n_1565), .B2(n_1568), .Y(n_1564) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_212), .Y(n_1101) );
INVx1_ASAP7_75t_L g1809 ( .A(n_213), .Y(n_1809) );
AOI221xp5_ASAP7_75t_L g1827 ( .A1(n_213), .A2(n_278), .B1(n_775), .B2(n_778), .C(n_1194), .Y(n_1827) );
INVx1_ASAP7_75t_L g940 ( .A(n_214), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g1340 ( .A(n_215), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_216), .A2(n_258), .B1(n_795), .B2(n_1203), .C(n_1205), .Y(n_1202) );
INVx1_ASAP7_75t_L g1230 ( .A(n_216), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_217), .A2(n_221), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx1_ASAP7_75t_L g1032 ( .A(n_217), .Y(n_1032) );
OA332x1_ASAP7_75t_L g998 ( .A1(n_218), .A2(n_410), .A3(n_999), .B1(n_1004), .B2(n_1007), .B3(n_1010), .C1(n_1015), .C2(n_1016), .Y(n_998) );
AOI21xp5_ASAP7_75t_L g1037 ( .A1(n_218), .A2(n_804), .B(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g813 ( .A(n_219), .Y(n_813) );
INVx1_ASAP7_75t_L g1518 ( .A(n_220), .Y(n_1518) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_221), .A2(n_292), .B1(n_455), .B2(n_614), .Y(n_1036) );
CKINVDCx16_ASAP7_75t_R g1578 ( .A(n_222), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_224), .A2(n_232), .B1(n_518), .B2(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1332 ( .A(n_224), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1841 ( .A1(n_225), .A2(n_1842), .B1(n_1843), .B2(n_1844), .Y(n_1841) );
CKINVDCx5p33_ASAP7_75t_R g1844 ( .A(n_225), .Y(n_1844) );
INVx1_ASAP7_75t_L g688 ( .A(n_226), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_227), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_228), .A2(n_231), .B1(n_654), .B2(n_656), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_228), .A2(n_231), .B1(n_403), .B2(n_680), .C(n_681), .Y(n_679) );
INVxp33_ASAP7_75t_SL g1456 ( .A(n_229), .Y(n_1456) );
INVx1_ASAP7_75t_L g1160 ( .A(n_230), .Y(n_1160) );
INVx1_ASAP7_75t_L g1330 ( .A(n_232), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_233), .A2(n_250), .B1(n_798), .B2(n_1174), .Y(n_1510) );
INVx1_ASAP7_75t_L g1525 ( .A(n_233), .Y(n_1525) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_234), .Y(n_947) );
INVx1_ASAP7_75t_L g1240 ( .A(n_236), .Y(n_1240) );
INVx1_ASAP7_75t_L g1368 ( .A(n_237), .Y(n_1368) );
OAI211xp5_ASAP7_75t_SL g1374 ( .A1(n_237), .A2(n_913), .B(n_1375), .C(n_1387), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_238), .A2(n_251), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g674 ( .A(n_238), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_239), .A2(n_325), .B1(n_480), .B2(n_483), .C(n_489), .Y(n_479) );
INVx1_ASAP7_75t_L g1071 ( .A(n_240), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g1297 ( .A(n_241), .Y(n_1297) );
INVx1_ASAP7_75t_L g1527 ( .A(n_242), .Y(n_1527) );
INVx1_ASAP7_75t_L g457 ( .A(n_243), .Y(n_457) );
BUFx3_ASAP7_75t_L g473 ( .A(n_243), .Y(n_473) );
INVxp67_ASAP7_75t_L g415 ( .A(n_244), .Y(n_415) );
AOI21xp33_ASAP7_75t_L g874 ( .A1(n_245), .A2(n_519), .B(n_804), .Y(n_874) );
INVx1_ASAP7_75t_L g899 ( .A(n_245), .Y(n_899) );
INVxp67_ASAP7_75t_SL g1479 ( .A(n_246), .Y(n_1479) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_247), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_247), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_247), .B(n_308), .Y(n_401) );
INVx1_ASAP7_75t_L g449 ( .A(n_247), .Y(n_449) );
INVx1_ASAP7_75t_L g918 ( .A(n_248), .Y(n_918) );
INVx1_ASAP7_75t_L g1698 ( .A(n_249), .Y(n_1698) );
INVx1_ASAP7_75t_L g1530 ( .A(n_250), .Y(n_1530) );
INVx1_ASAP7_75t_L g676 ( .A(n_251), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_252), .A2(n_792), .B1(n_853), .B2(n_858), .C(n_864), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_253), .Y(n_944) );
INVx1_ASAP7_75t_L g1583 ( .A(n_255), .Y(n_1583) );
OR2x2_ASAP7_75t_L g460 ( .A(n_256), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g468 ( .A(n_256), .Y(n_468) );
INVx1_ASAP7_75t_L g1696 ( .A(n_257), .Y(n_1696) );
INVx1_ASAP7_75t_L g1228 ( .A(n_258), .Y(n_1228) );
INVx1_ASAP7_75t_L g900 ( .A(n_259), .Y(n_900) );
INVx1_ASAP7_75t_L g1140 ( .A(n_260), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_261), .A2(n_275), .B1(n_363), .B2(n_841), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_261), .A2(n_275), .B1(n_535), .B2(n_866), .Y(n_1425) );
INVxp67_ASAP7_75t_L g1148 ( .A(n_262), .Y(n_1148) );
CKINVDCx16_ASAP7_75t_R g1580 ( .A(n_264), .Y(n_1580) );
INVx1_ASAP7_75t_L g1412 ( .A(n_265), .Y(n_1412) );
AOI21xp33_ASAP7_75t_L g1430 ( .A1(n_265), .A2(n_515), .B(n_767), .Y(n_1430) );
INVx1_ASAP7_75t_L g1588 ( .A(n_266), .Y(n_1588) );
INVxp67_ASAP7_75t_L g748 ( .A(n_267), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_268), .A2(n_302), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
INVx1_ASAP7_75t_L g1217 ( .A(n_268), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_269), .A2(n_273), .B1(n_597), .B2(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g621 ( .A(n_269), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_270), .A2(n_290), .B1(n_646), .B2(n_648), .C(n_1177), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_272), .Y(n_1208) );
INVx1_ASAP7_75t_L g635 ( .A(n_273), .Y(n_635) );
INVx1_ASAP7_75t_L g859 ( .A(n_274), .Y(n_859) );
INVxp67_ASAP7_75t_SL g1453 ( .A(n_276), .Y(n_1453) );
INVxp67_ASAP7_75t_SL g1801 ( .A(n_277), .Y(n_1801) );
INVx1_ASAP7_75t_L g1808 ( .A(n_278), .Y(n_1808) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_279), .A2(n_849), .B1(n_904), .B2(n_905), .Y(n_848) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_279), .Y(n_904) );
INVx1_ASAP7_75t_L g1221 ( .A(n_280), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_281), .Y(n_540) );
INVxp33_ASAP7_75t_L g719 ( .A(n_282), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g1371 ( .A1(n_283), .A2(n_319), .B1(n_963), .B2(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1389 ( .A(n_283), .Y(n_1389) );
OAI221xp5_ASAP7_75t_SL g1806 ( .A1(n_284), .A2(n_318), .B1(n_742), .B2(n_835), .C(n_1807), .Y(n_1806) );
AOI22xp33_ASAP7_75t_L g1828 ( .A1(n_284), .A2(n_318), .B1(n_633), .B2(n_863), .Y(n_1828) );
INVx1_ASAP7_75t_L g1157 ( .A(n_285), .Y(n_1157) );
INVx1_ASAP7_75t_L g1574 ( .A(n_286), .Y(n_1574) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_287), .Y(n_1013) );
INVx1_ASAP7_75t_L g1327 ( .A(n_289), .Y(n_1327) );
OAI332xp33_ASAP7_75t_L g1136 ( .A1(n_290), .A2(n_410), .A3(n_845), .B1(n_1021), .B2(n_1137), .B3(n_1141), .C1(n_1144), .C2(n_1149), .Y(n_1136) );
INVx1_ASAP7_75t_L g1001 ( .A(n_291), .Y(n_1001) );
INVx1_ASAP7_75t_L g1114 ( .A(n_293), .Y(n_1114) );
INVx1_ASAP7_75t_L g1142 ( .A(n_294), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
AND3x2_ASAP7_75t_L g1547 ( .A(n_295), .B(n_335), .C(n_1548), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1554 ( .A(n_295), .B(n_335), .Y(n_1554) );
INVx2_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_299), .A2(n_321), .B1(n_483), .B2(n_646), .Y(n_661) );
INVx1_ASAP7_75t_L g687 ( .A(n_299), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_300), .A2(n_913), .B(n_917), .C(n_922), .Y(n_912) );
INVx1_ASAP7_75t_L g974 ( .A(n_300), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_301), .A2(n_314), .B1(n_777), .B2(n_1026), .Y(n_1207) );
INVx1_ASAP7_75t_L g1226 ( .A(n_301), .Y(n_1226) );
INVx1_ASAP7_75t_L g1222 ( .A(n_302), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_305), .Y(n_1395) );
INVx1_ASAP7_75t_L g350 ( .A(n_308), .Y(n_350) );
INVx2_ASAP7_75t_L g370 ( .A(n_308), .Y(n_370) );
OR2x2_ASAP7_75t_L g850 ( .A(n_309), .B(n_544), .Y(n_850) );
INVx1_ASAP7_75t_L g604 ( .A(n_311), .Y(n_604) );
INVx1_ASAP7_75t_L g1344 ( .A(n_313), .Y(n_1344) );
INVx1_ASAP7_75t_L g1231 ( .A(n_314), .Y(n_1231) );
INVx1_ASAP7_75t_L g1589 ( .A(n_315), .Y(n_1589) );
INVx1_ASAP7_75t_L g802 ( .A(n_316), .Y(n_802) );
INVx1_ASAP7_75t_L g1055 ( .A(n_317), .Y(n_1055) );
INVx1_ASAP7_75t_L g1388 ( .A(n_319), .Y(n_1388) );
INVx1_ASAP7_75t_L g696 ( .A(n_321), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_322), .Y(n_1211) );
INVx1_ASAP7_75t_L g871 ( .A(n_323), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_324), .Y(n_1006) );
INVxp33_ASAP7_75t_SL g385 ( .A(n_325), .Y(n_385) );
INVx1_ASAP7_75t_L g1067 ( .A(n_326), .Y(n_1067) );
INVx1_ASAP7_75t_L g788 ( .A(n_328), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_351), .B(n_1535), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_338), .Y(n_332) );
AND2x4_ASAP7_75t_L g1838 ( .A(n_333), .B(n_339), .Y(n_1838) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_SL g1848 ( .A(n_334), .Y(n_1848) );
NAND2xp5_ASAP7_75t_L g1851 ( .A(n_334), .B(n_336), .Y(n_1851) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g1847 ( .A(n_336), .B(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g580 ( .A(n_342), .B(n_350), .Y(n_580) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g411 ( .A(n_343), .B(n_412), .Y(n_411) );
OR2x6_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g417 ( .A(n_345), .Y(n_417) );
OR2x2_ASAP7_75t_L g545 ( .A(n_345), .B(n_400), .Y(n_545) );
BUFx2_ASAP7_75t_L g686 ( .A(n_345), .Y(n_686) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_345), .Y(n_733) );
INVx2_ASAP7_75t_SL g829 ( .A(n_345), .Y(n_829) );
INVx2_ASAP7_75t_SL g946 ( .A(n_345), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g1800 ( .A1(n_345), .A2(n_421), .B1(n_1801), .B2(n_1802), .Y(n_1800) );
OAI22xp33_ASAP7_75t_L g1811 ( .A1(n_345), .A2(n_421), .B1(n_1812), .B2(n_1813), .Y(n_1811) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g364 ( .A(n_347), .Y(n_364) );
INVx1_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
AND2x2_ASAP7_75t_L g384 ( .A(n_347), .B(n_348), .Y(n_384) );
AND2x4_ASAP7_75t_L g391 ( .A(n_347), .B(n_377), .Y(n_391) );
INVx1_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
INVx1_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
INVx2_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx1_ASAP7_75t_L g398 ( .A(n_348), .Y(n_398) );
INVx1_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_348), .B(n_364), .Y(n_431) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_1125), .B2(n_1126), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
XNOR2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_710), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
XNOR2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_550), .Y(n_355) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_450), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g358 ( .A(n_359), .B(n_392), .C(n_408), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_361), .A2(n_381), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_361), .A2(n_372), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
AND2x2_ASAP7_75t_L g575 ( .A(n_362), .B(n_367), .Y(n_575) );
INVx2_ASAP7_75t_SL g593 ( .A(n_362), .Y(n_593) );
AND2x2_ASAP7_75t_L g678 ( .A(n_362), .B(n_367), .Y(n_678) );
AND2x2_ASAP7_75t_L g725 ( .A(n_362), .B(n_367), .Y(n_725) );
AND2x2_ASAP7_75t_L g824 ( .A(n_362), .B(n_367), .Y(n_824) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g887 ( .A(n_363), .Y(n_887) );
AND2x2_ASAP7_75t_L g919 ( .A(n_363), .B(n_369), .Y(n_919) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_363), .Y(n_924) );
BUFx6f_ASAP7_75t_L g1799 ( .A(n_363), .Y(n_1799) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g406 ( .A(n_364), .Y(n_406) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x6_ASAP7_75t_L g373 ( .A(n_367), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g381 ( .A(n_367), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g388 ( .A(n_367), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g818 ( .A(n_367), .B(n_695), .Y(n_818) );
AND2x2_ASAP7_75t_L g820 ( .A(n_367), .B(n_587), .Y(n_820) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_367), .B(n_956), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1805 ( .A1(n_367), .A2(n_895), .B1(n_1806), .B2(n_1810), .Y(n_1805) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g446 ( .A(n_368), .Y(n_446) );
OR2x2_ASAP7_75t_L g985 ( .A(n_368), .B(n_460), .Y(n_985) );
INVx2_ASAP7_75t_L g916 ( .A(n_369), .Y(n_916) );
AND2x4_ASAP7_75t_L g936 ( .A(n_369), .B(n_591), .Y(n_936) );
INVx1_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
INVx1_ASAP7_75t_L g448 ( .A(n_370), .Y(n_448) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_373), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_373), .A2(n_388), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_373), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_373), .A2(n_1217), .B1(n_1218), .B2(n_1219), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_373), .A2(n_570), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_373), .A2(n_570), .B1(n_1503), .B2(n_1518), .Y(n_1517) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_374), .B(n_399), .Y(n_407) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g567 ( .A(n_375), .Y(n_567) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_375), .Y(n_587) );
BUFx3_ASAP7_75t_L g884 ( .A(n_375), .Y(n_884) );
BUFx6f_ASAP7_75t_L g1385 ( .A(n_375), .Y(n_1385) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_385), .B2(n_386), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_379), .A2(n_490), .B1(n_495), .B2(n_496), .C(n_499), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_380), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1251) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_381), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_381), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_381), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_381), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_381), .A2(n_725), .B1(n_899), .B2(n_900), .C(n_901), .Y(n_898) );
INVx1_ASAP7_75t_L g1181 ( .A(n_381), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_381), .A2(n_678), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_381), .A2(n_678), .B1(n_1504), .B2(n_1520), .Y(n_1519) );
BUFx3_ASAP7_75t_L g597 ( .A(n_382), .Y(n_597) );
BUFx2_ASAP7_75t_L g882 ( .A(n_382), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g1807 ( .A1(n_382), .A2(n_567), .B1(n_1808), .B2(n_1809), .Y(n_1807) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g956 ( .A(n_383), .Y(n_956) );
INVx2_ASAP7_75t_L g1260 ( .A(n_383), .Y(n_1260) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_384), .Y(n_591) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g570 ( .A(n_388), .Y(n_570) );
BUFx2_ASAP7_75t_L g720 ( .A(n_388), .Y(n_720) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_388), .Y(n_1183) );
BUFx2_ASAP7_75t_L g1218 ( .A(n_388), .Y(n_1218) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_388), .Y(n_1254) );
BUFx3_ASAP7_75t_L g434 ( .A(n_389), .Y(n_434) );
INVx2_ASAP7_75t_L g835 ( .A(n_389), .Y(n_835) );
INVx1_ASAP7_75t_L g941 ( .A(n_389), .Y(n_941) );
INVx1_ASAP7_75t_SL g1413 ( .A(n_389), .Y(n_1413) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g695 ( .A(n_390), .Y(n_695) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_390), .Y(n_747) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_391), .Y(n_584) );
INVx1_ASAP7_75t_L g842 ( .A(n_391), .Y(n_842) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g727 ( .A(n_394), .Y(n_727) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_395), .Y(n_680) );
NAND2x1_ASAP7_75t_SL g395 ( .A(n_396), .B(n_399), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g929 ( .A(n_396), .B(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_396), .A2(n_405), .B1(n_1318), .B2(n_1320), .Y(n_1346) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_398), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_399), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g557 ( .A(n_399), .B(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g563 ( .A(n_399), .B(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g566 ( .A(n_399), .B(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g932 ( .A(n_401), .Y(n_932) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx4f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_404), .Y(n_728) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x6_ASAP7_75t_L g933 ( .A(n_406), .B(n_931), .Y(n_933) );
BUFx3_ASAP7_75t_L g681 ( .A(n_407), .Y(n_681) );
BUFx2_ASAP7_75t_L g729 ( .A(n_407), .Y(n_729) );
BUFx2_ASAP7_75t_L g1522 ( .A(n_407), .Y(n_1522) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_414), .A3(n_425), .B1(n_435), .B2(n_438), .B3(n_443), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI33xp33_ASAP7_75t_L g682 ( .A1(n_410), .A2(n_443), .A3(n_683), .B1(n_689), .B2(n_697), .B3(n_701), .Y(n_682) );
OAI33xp33_ASAP7_75t_L g730 ( .A1(n_410), .A2(n_443), .A3(n_731), .B1(n_739), .B2(n_749), .B3(n_754), .Y(n_730) );
OAI33xp33_ASAP7_75t_L g826 ( .A1(n_410), .A2(n_827), .A3(n_832), .B1(n_837), .B2(n_843), .B3(n_845), .Y(n_826) );
OAI33xp33_ASAP7_75t_L g1224 ( .A1(n_410), .A2(n_845), .A3(n_1225), .B1(n_1229), .B2(n_1233), .B3(n_1239), .Y(n_1224) );
OAI33xp33_ASAP7_75t_L g1523 ( .A1(n_410), .A2(n_443), .A3(n_1524), .B1(n_1528), .B2(n_1531), .B3(n_1533), .Y(n_1523) );
OR2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
BUFx2_ASAP7_75t_L g539 ( .A(n_413), .Y(n_539) );
INVx2_ASAP7_75t_L g579 ( .A(n_413), .Y(n_579) );
OAI22xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B1(n_418), .B2(n_419), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_416), .A2(n_427), .B1(n_436), .B2(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g755 ( .A(n_417), .Y(n_755) );
INVx1_ASAP7_75t_L g1227 ( .A(n_417), .Y(n_1227) );
OAI22xp5_ASAP7_75t_SL g1149 ( .A1(n_419), .A2(n_755), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
BUFx3_ASAP7_75t_L g844 ( .A(n_421), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_421), .A2(n_733), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_421), .A2(n_755), .B1(n_1339), .B2(n_1340), .C(n_1341), .Y(n_1338) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x2_ASAP7_75t_L g705 ( .A(n_423), .B(n_424), .Y(n_705) );
INVx1_ASAP7_75t_L g559 ( .A(n_424), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_432), .B2(n_433), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_427), .A2(n_1097), .B1(n_1098), .B2(n_1101), .Y(n_1096) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g1333 ( .A1(n_428), .A2(n_1334), .B1(n_1335), .B2(n_1337), .Y(n_1333) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g833 ( .A(n_429), .Y(n_833) );
INVx2_ASAP7_75t_L g1139 ( .A(n_429), .Y(n_1139) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g742 ( .A(n_430), .Y(n_742) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g692 ( .A(n_431), .Y(n_692) );
BUFx2_ASAP7_75t_L g939 ( .A(n_431), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_433), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g1262 ( .A(n_434), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_436), .A2(n_439), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_437), .A2(n_453), .B(n_462), .C(n_479), .Y(n_452) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_441), .A2(n_684), .B1(n_687), .B2(n_688), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_441), .A2(n_945), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1524 ( .A1(n_441), .A2(n_1525), .B1(n_1526), .B2(n_1527), .Y(n_1524) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_442), .A2(n_502), .B1(n_508), .B2(n_517), .C(n_525), .Y(n_501) );
INVx1_ASAP7_75t_L g1268 ( .A(n_443), .Y(n_1268) );
CKINVDCx8_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx6_ASAP7_75t_L g599 ( .A(n_445), .Y(n_599) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g962 ( .A(n_446), .B(n_465), .Y(n_962) );
INVx2_ASAP7_75t_L g896 ( .A(n_447), .Y(n_896) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_447), .Y(n_1386) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_536), .B1(n_540), .B2(n_541), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_501), .C(n_531), .Y(n_451) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI211xp5_ASAP7_75t_SL g603 ( .A1(n_454), .A2(n_604), .B(n_605), .C(n_609), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g761 ( .A1(n_454), .A2(n_751), .B(n_762), .C(n_764), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_454), .A2(n_1191), .B1(n_1195), .B2(n_1198), .C(n_1199), .Y(n_1190) );
AOI211xp5_ASAP7_75t_L g1273 ( .A1(n_454), .A2(n_1274), .B(n_1275), .C(n_1276), .Y(n_1273) );
AOI211xp5_ASAP7_75t_L g1470 ( .A1(n_454), .A2(n_1471), .B(n_1472), .C(n_1474), .Y(n_1470) );
AOI211xp5_ASAP7_75t_SL g1496 ( .A1(n_454), .A2(n_1497), .B(n_1498), .C(n_1500), .Y(n_1496) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
INVx2_ASAP7_75t_SL g773 ( .A(n_455), .Y(n_773) );
BUFx3_ASAP7_75t_L g1370 ( .A(n_455), .Y(n_1370) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx3_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_456), .Y(n_612) );
BUFx2_ASAP7_75t_L g660 ( .A(n_456), .Y(n_660) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_456), .Y(n_767) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_456), .Y(n_806) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_456), .Y(n_863) );
INVx2_ASAP7_75t_SL g983 ( .A(n_456), .Y(n_983) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_456), .Y(n_1501) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g494 ( .A(n_457), .Y(n_494) );
INVx2_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
AND2x2_ASAP7_75t_L g507 ( .A(n_458), .B(n_473), .Y(n_507) );
AND2x4_ASAP7_75t_L g505 ( .A(n_459), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g651 ( .A(n_459), .B(n_612), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_459), .A2(n_505), .B1(n_663), .B2(n_1151), .C(n_1163), .Y(n_1162) );
AOI222xp33_ASAP7_75t_L g1815 ( .A1(n_459), .A2(n_655), .B1(n_657), .B2(n_1795), .C1(n_1796), .C2(n_1816), .Y(n_1815) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g533 ( .A(n_460), .B(n_498), .Y(n_533) );
OR2x2_ASAP7_75t_L g535 ( .A(n_460), .B(n_486), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g1024 ( .A1(n_460), .A2(n_1025), .B(n_1027), .C(n_1029), .Y(n_1024) );
INVx1_ASAP7_75t_L g466 ( .A(n_461), .Y(n_466) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g606 ( .A(n_464), .Y(n_606) );
INVx1_ASAP7_75t_L g763 ( .A(n_464), .Y(n_763) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_464), .Y(n_1046) );
INVx1_ASAP7_75t_L g1200 ( .A(n_464), .Y(n_1200) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
AND2x2_ASAP7_75t_L g475 ( .A(n_465), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
AND2x2_ASAP7_75t_L g549 ( .A(n_465), .B(n_521), .Y(n_549) );
AND2x2_ASAP7_75t_L g608 ( .A(n_465), .B(n_476), .Y(n_608) );
AND2x4_ASAP7_75t_L g655 ( .A(n_465), .B(n_469), .Y(n_655) );
AND2x4_ASAP7_75t_L g657 ( .A(n_465), .B(n_476), .Y(n_657) );
BUFx2_ASAP7_75t_L g664 ( .A(n_465), .Y(n_664) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x4_ASAP7_75t_L g499 ( .A(n_467), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g516 ( .A(n_468), .B(n_500), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_469), .A2(n_476), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g960 ( .A(n_470), .Y(n_960) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g521 ( .A(n_472), .B(n_478), .Y(n_521) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g487 ( .A(n_473), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g964 ( .A(n_476), .Y(n_964) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g1174 ( .A(n_484), .Y(n_1174) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g779 ( .A(n_485), .Y(n_779) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1434 ( .A(n_486), .Y(n_1434) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_487), .Y(n_524) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_487), .Y(n_614) );
INVx1_ASAP7_75t_L g991 ( .A(n_487), .Y(n_991) );
INVx1_ASAP7_75t_L g1279 ( .A(n_487), .Y(n_1279) );
INVx1_ASAP7_75t_L g493 ( .A(n_488), .Y(n_493) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g616 ( .A(n_492), .Y(n_616) );
BUFx4f_ASAP7_75t_L g861 ( .A(n_492), .Y(n_861) );
INVx2_ASAP7_75t_L g993 ( .A(n_492), .Y(n_993) );
INVx1_ASAP7_75t_L g1035 ( .A(n_492), .Y(n_1035) );
INVx1_ASAP7_75t_L g1070 ( .A(n_492), .Y(n_1070) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
OR2x2_ASAP7_75t_L g498 ( .A(n_493), .B(n_494), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g1076 ( .A1(n_496), .A2(n_1077), .B1(n_1078), .B2(n_1080), .C(n_1081), .Y(n_1076) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g769 ( .A(n_497), .Y(n_769) );
INVx2_ASAP7_75t_L g854 ( .A(n_497), .Y(n_854) );
INVx1_ASAP7_75t_L g1121 ( .A(n_497), .Y(n_1121) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g618 ( .A(n_498), .Y(n_618) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_498), .Y(n_1066) );
INVx1_ASAP7_75t_L g1165 ( .A(n_498), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_499), .Y(n_619) );
INVx1_ASAP7_75t_L g648 ( .A(n_499), .Y(n_648) );
INVx2_ASAP7_75t_SL g804 ( .A(n_499), .Y(n_804) );
AND2x4_ASAP7_75t_L g971 ( .A(n_499), .B(n_548), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_499), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1502 ( .A1(n_499), .A2(n_1035), .B1(n_1121), .B2(n_1503), .C(n_1504), .Y(n_1502) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_504), .A2(n_527), .B1(n_621), .B2(n_622), .C(n_627), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_504), .A2(n_527), .B1(n_753), .B2(n_771), .C(n_776), .Y(n_770) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_504), .A2(n_663), .B1(n_1202), .B2(n_1207), .C(n_1208), .Y(n_1201) );
AOI221xp5_ASAP7_75t_L g1478 ( .A1(n_504), .A2(n_527), .B1(n_1479), .B2(n_1480), .C(n_1485), .Y(n_1478) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_505), .A2(n_659), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_658) );
INVx2_ASAP7_75t_SL g792 ( .A(n_505), .Y(n_792) );
HB1xp67_ASAP7_75t_L g1283 ( .A(n_505), .Y(n_1283) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_505), .A2(n_663), .B1(n_1506), .B2(n_1507), .C(n_1510), .Y(n_1505) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_506), .Y(n_626) );
AND2x4_ASAP7_75t_L g663 ( .A(n_506), .B(n_664), .Y(n_663) );
BUFx4f_ASAP7_75t_L g1028 ( .A(n_506), .Y(n_1028) );
INVx1_ASAP7_75t_L g1178 ( .A(n_506), .Y(n_1178) );
BUFx3_ASAP7_75t_L g1192 ( .A(n_506), .Y(n_1192) );
INVx2_ASAP7_75t_SL g1206 ( .A(n_506), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g1817 ( .A1(n_506), .A2(n_612), .B1(n_1813), .B2(n_1818), .Y(n_1817) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_507), .Y(n_513) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g647 ( .A(n_512), .Y(n_647) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_513), .Y(n_530) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_513), .Y(n_775) );
INVx1_ASAP7_75t_L g978 ( .A(n_513), .Y(n_978) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g1484 ( .A(n_515), .Y(n_1484) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g796 ( .A(n_516), .Y(n_796) );
INVx1_ASAP7_75t_L g967 ( .A(n_516), .Y(n_967) );
INVx1_ASAP7_75t_L g1044 ( .A(n_516), .Y(n_1044) );
INVx2_ASAP7_75t_L g1064 ( .A(n_516), .Y(n_1064) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g987 ( .A(n_519), .B(n_984), .Y(n_987) );
A2O1A1Ixp33_ASAP7_75t_L g1439 ( .A1(n_519), .A2(n_1440), .B(n_1441), .C(n_1445), .Y(n_1439) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g1038 ( .A(n_520), .Y(n_1038) );
INVx1_ASAP7_75t_L g1486 ( .A(n_520), .Y(n_1486) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx6_ASAP7_75t_L g631 ( .A(n_521), .Y(n_631) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_521), .Y(n_1292) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI221xp5_ASAP7_75t_SL g1167 ( .A1(n_523), .A2(n_1140), .B1(n_1143), .B2(n_1164), .C(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_524), .Y(n_633) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_524), .Y(n_800) );
INVx1_ASAP7_75t_L g808 ( .A(n_524), .Y(n_808) );
BUFx6f_ASAP7_75t_L g1026 ( .A(n_524), .Y(n_1026) );
INVx2_ASAP7_75t_L g1166 ( .A(n_524), .Y(n_1166) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_527), .A2(n_1283), .B1(n_1284), .B2(n_1285), .C(n_1290), .Y(n_1282) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_529), .B(n_964), .Y(n_1473) );
INVx1_ASAP7_75t_L g1312 ( .A(n_530), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_532), .A2(n_534), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_532), .A2(n_534), .B1(n_666), .B2(n_667), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_532), .A2(n_534), .B1(n_756), .B2(n_757), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_532), .A2(n_534), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_532), .A2(n_534), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_532), .A2(n_534), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_532), .A2(n_534), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_532), .A2(n_534), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
INVx6_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx5_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g911 ( .A1(n_537), .A2(n_912), .B(n_934), .Y(n_911) );
BUFx8_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g1188 ( .A(n_538), .Y(n_1188) );
AOI31xp33_ASAP7_75t_L g1272 ( .A1(n_538), .A2(n_1273), .A3(n_1282), .B(n_1294), .Y(n_1272) );
OAI31xp33_ASAP7_75t_L g1321 ( .A1(n_538), .A2(n_1322), .A3(n_1324), .B(n_1347), .Y(n_1321) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g638 ( .A(n_539), .Y(n_638) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_543), .A2(n_601), .B(n_602), .Y(n_600) );
AOI21xp33_ASAP7_75t_SL g758 ( .A1(n_543), .A2(n_759), .B(n_760), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g1467 ( .A1(n_543), .A2(n_1468), .B(n_1469), .Y(n_1467) );
INVx5_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g669 ( .A(n_544), .Y(n_669) );
INVx1_ASAP7_75t_L g1213 ( .A(n_544), .Y(n_1213) );
INVx2_ASAP7_75t_L g1270 ( .A(n_544), .Y(n_1270) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g1804 ( .A(n_545), .Y(n_1804) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x6_ASAP7_75t_L g952 ( .A(n_547), .B(n_953), .Y(n_952) );
AOI222xp33_ASAP7_75t_L g1349 ( .A1(n_547), .A2(n_987), .B1(n_1337), .B2(n_1340), .C1(n_1344), .C2(n_1350), .Y(n_1349) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_549), .B(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1156 ( .A(n_549), .Y(n_1156) );
AO22x2_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_639), .B1(n_708), .B2(n_709), .Y(n_550) );
INVx1_ASAP7_75t_L g709 ( .A(n_551), .Y(n_709) );
XNOR2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_600), .Y(n_553) );
AND4x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_568), .C(n_572), .D(n_576), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B1(n_561), .B2(n_565), .C(n_566), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g1452 ( .A1(n_556), .A2(n_561), .B1(n_566), .B2(n_1453), .C(n_1454), .Y(n_1452) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_557), .A2(n_563), .B1(n_566), .B2(n_868), .C(n_869), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_557), .A2(n_563), .B1(n_566), .B2(n_1050), .C(n_1051), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g1245 ( .A1(n_557), .A2(n_563), .B1(n_566), .B2(n_1246), .C(n_1247), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1794 ( .A1(n_557), .A2(n_563), .B1(n_566), .B2(n_1795), .C(n_1796), .Y(n_1794) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g1184 ( .A1(n_563), .A2(n_566), .B(n_1160), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_564), .B(n_955), .Y(n_1113) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_567), .Y(n_1265) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_571), .A2(n_573), .B1(n_616), .B2(n_617), .C(n_619), .Y(n_615) );
AOI33xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .A3(n_588), .B1(n_594), .B2(n_596), .B3(n_599), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g1257 ( .A(n_578), .Y(n_1257) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g642 ( .A(n_579), .Y(n_642) );
BUFx2_ASAP7_75t_L g812 ( .A(n_579), .Y(n_812) );
AND2x4_ASAP7_75t_L g880 ( .A(n_579), .B(n_580), .Y(n_880) );
AND2x2_ASAP7_75t_L g895 ( .A(n_579), .B(n_896), .Y(n_895) );
OR2x2_ASAP7_75t_L g966 ( .A(n_579), .B(n_967), .Y(n_966) );
OR2x6_ASAP7_75t_L g1063 ( .A(n_579), .B(n_1064), .Y(n_1063) );
BUFx2_ASAP7_75t_SL g948 ( .A(n_580), .Y(n_948) );
INVx1_ASAP7_75t_L g1095 ( .A(n_580), .Y(n_1095) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_583), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g1137 ( .A1(n_583), .A2(n_1138), .B1(n_1139), .B2(n_1140), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1531 ( .A1(n_583), .A2(n_1497), .B1(n_1513), .B2(n_1532), .Y(n_1531) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g595 ( .A(n_584), .Y(n_595) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_584), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1397 ( .A(n_584), .Y(n_1397) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
INVx2_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g894 ( .A(n_590), .Y(n_894) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_591), .Y(n_926) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g1232 ( .A(n_595), .Y(n_1232) );
INVx2_ASAP7_75t_L g845 ( .A(n_599), .Y(n_845) );
INVx1_ASAP7_75t_L g1015 ( .A(n_599), .Y(n_1015) );
AOI33xp33_ASAP7_75t_L g1461 ( .A1(n_599), .A2(n_1256), .A3(n_1462), .B1(n_1463), .B2(n_1465), .B3(n_1466), .Y(n_1461) );
AOI31xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_620), .A3(n_634), .B(n_637), .Y(n_602) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_611), .B(n_985), .Y(n_1122) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g624 ( .A(n_612), .Y(n_624) );
BUFx2_ASAP7_75t_L g1365 ( .A(n_612), .Y(n_1365) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_614), .Y(n_650) );
INVx1_ASAP7_75t_L g856 ( .A(n_614), .Y(n_856) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_616), .A2(n_619), .B1(n_721), .B2(n_723), .C(n_769), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g1435 ( .A1(n_616), .A2(n_1436), .B(n_1437), .C(n_1438), .Y(n_1435) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_617), .A2(n_860), .B1(n_973), .B2(n_974), .C(n_975), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_617), .A2(n_1414), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g1477 ( .A1(n_619), .A2(n_769), .B1(n_993), .B2(n_1457), .C(n_1459), .Y(n_1477) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g1482 ( .A(n_626), .Y(n_1482) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx6f_ASAP7_75t_L g1824 ( .A(n_630), .Y(n_1824) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g646 ( .A(n_631), .Y(n_646) );
INVx2_ASAP7_75t_L g778 ( .A(n_631), .Y(n_778) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_631), .Y(n_799) );
INVx1_ASAP7_75t_L g1042 ( .A(n_631), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g1075 ( .A(n_633), .Y(n_1075) );
AOI31xp33_ASAP7_75t_L g760 ( .A1(n_637), .A2(n_761), .A3(n_770), .B(n_780), .Y(n_760) );
INVx1_ASAP7_75t_L g1179 ( .A(n_637), .Y(n_1179) );
AOI31xp33_ASAP7_75t_L g1469 ( .A1(n_637), .A2(n_1470), .A3(n_1478), .B(n_1487), .Y(n_1469) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI31xp33_ASAP7_75t_L g1023 ( .A1(n_638), .A2(n_1024), .A3(n_1030), .B(n_1045), .Y(n_1023) );
INVx3_ASAP7_75t_L g708 ( .A(n_639), .Y(n_708) );
INVx1_ASAP7_75t_L g706 ( .A(n_640), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_670), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_668), .B2(n_669), .Y(n_641) );
INVx2_ASAP7_75t_L g877 ( .A(n_642), .Y(n_877) );
NOR2xp67_ASAP7_75t_L g953 ( .A(n_642), .B(n_954), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1494 ( .A1(n_642), .A2(n_1270), .B1(n_1495), .B2(n_1514), .Y(n_1494) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_658), .C(n_665), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_651), .B2(n_652), .C(n_653), .Y(n_644) );
INVx1_ASAP7_75t_L g1287 ( .A(n_647), .Y(n_1287) );
INVx1_ASAP7_75t_L g1281 ( .A(n_648), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_651), .A2(n_802), .B1(n_803), .B2(n_805), .C(n_809), .Y(n_801) );
INVx1_ASAP7_75t_L g866 ( .A(n_651), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_652), .A2(n_667), .B1(n_690), .B2(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g810 ( .A(n_655), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_655), .A2(n_657), .B1(n_868), .B2(n_869), .Y(n_867) );
INVx4_ASAP7_75t_L g1159 ( .A(n_655), .Y(n_1159) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AOI222xp33_ASAP7_75t_SL g1154 ( .A1(n_657), .A2(n_1155), .B1(n_1157), .B2(n_1158), .C1(n_1160), .C2(n_1161), .Y(n_1154) );
INVx2_ASAP7_75t_L g1499 ( .A(n_657), .Y(n_1499) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_662), .A2(n_666), .B1(n_684), .B2(n_702), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_663), .A2(n_791), .B1(n_793), .B2(n_794), .C(n_797), .Y(n_790) );
INVx1_ASAP7_75t_L g864 ( .A(n_663), .Y(n_864) );
INVx1_ASAP7_75t_L g1029 ( .A(n_663), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1819 ( .A1(n_663), .A2(n_1820), .B(n_1823), .Y(n_1819) );
BUFx3_ASAP7_75t_L g1445 ( .A(n_664), .Y(n_1445) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_669), .A2(n_786), .B1(n_811), .B2(n_813), .Y(n_785) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_679), .C(n_682), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .Y(n_671) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g1331 ( .A(n_685), .Y(n_1331) );
INVx1_ASAP7_75t_L g1526 ( .A(n_685), .Y(n_1526) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B1(n_694), .B2(n_696), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g1528 ( .A1(n_690), .A2(n_1335), .B1(n_1529), .B2(n_1530), .Y(n_1528) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_691), .Y(n_1012) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_692), .Y(n_839) );
INVx1_ASAP7_75t_L g1236 ( .A(n_692), .Y(n_1236) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g700 ( .A(n_695), .Y(n_700) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_695), .Y(n_1003) );
INVx1_ASAP7_75t_L g1100 ( .A(n_695), .Y(n_1100) );
INVx2_ASAP7_75t_L g1380 ( .A(n_695), .Y(n_1380) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g888 ( .A(n_700), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_702), .A2(n_828), .B1(n_830), .B2(n_831), .Y(n_827) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x6_ASAP7_75t_L g949 ( .A(n_704), .B(n_931), .Y(n_949) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_704), .B(n_931), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_704), .A2(n_945), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g737 ( .A(n_705), .Y(n_737) );
INVx2_ASAP7_75t_L g1329 ( .A(n_705), .Y(n_1329) );
BUFx2_ASAP7_75t_L g1393 ( .A(n_705), .Y(n_1393) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_907), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_782), .B2(n_906), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
XNOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_781), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_758), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_726), .C(n_730), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_722), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_735), .B2(n_738), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_732), .A2(n_844), .B1(n_1208), .B2(n_1210), .Y(n_1239) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_733), .A2(n_788), .B1(n_793), .B2(n_844), .Y(n_843) );
OAI22xp33_ASAP7_75t_L g1533 ( .A1(n_733), .A2(n_1329), .B1(n_1506), .B2(n_1512), .Y(n_1533) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g752 ( .A(n_737), .Y(n_752) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_737), .A2(n_944), .B1(n_945), .B2(n_947), .C(n_948), .Y(n_943) );
AOI21xp33_ASAP7_75t_L g1345 ( .A1(n_737), .A2(n_931), .B(n_1346), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_744), .B2(n_748), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_740), .A2(n_1014), .B1(n_1105), .B2(n_1106), .C(n_1107), .Y(n_1104) );
OAI22xp5_ASAP7_75t_SL g1229 ( .A1(n_740), .A2(n_1230), .B1(n_1231), .B2(n_1232), .Y(n_1229) );
OAI22xp5_ASAP7_75t_SL g1394 ( .A1(n_740), .A2(n_1395), .B1(n_1396), .B2(n_1397), .Y(n_1394) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g750 ( .A(n_741), .Y(n_750) );
INVx1_ASAP7_75t_L g1376 ( .A(n_741), .Y(n_1376) );
INVx2_ASAP7_75t_L g1532 ( .A(n_741), .Y(n_1532) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g1238 ( .A(n_747), .Y(n_1238) );
INVx2_ASAP7_75t_L g1336 ( .A(n_747), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_752), .A2(n_945), .B1(n_1067), .B2(n_1071), .C(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
BUFx3_ASAP7_75t_L g1171 ( .A(n_767), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_769), .A2(n_860), .B1(n_944), .B2(n_947), .C(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g1073 ( .A(n_773), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_778), .A2(n_1008), .B1(n_1013), .B2(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g906 ( .A(n_782), .Y(n_906) );
XOR2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_848), .Y(n_782) );
INVx1_ASAP7_75t_L g846 ( .A(n_784), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_814), .Y(n_784) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_790), .C(n_801), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_789), .A2(n_802), .B1(n_838), .B2(n_840), .Y(n_837) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g1509 ( .A(n_796), .Y(n_1509) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx4_ASAP7_75t_L g1193 ( .A(n_799), .Y(n_1193) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g1825 ( .A(n_808), .Y(n_1825) );
CKINVDCx8_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_825), .C(n_826), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_816), .B(n_821), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_816) );
INVx2_ASAP7_75t_L g902 ( .A(n_818), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_820), .Y(n_903) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_820), .Y(n_1021) );
INVx1_ASAP7_75t_L g1020 ( .A(n_824), .Y(n_1020) );
INVx1_ASAP7_75t_L g1135 ( .A(n_824), .Y(n_1135) );
INVx1_ASAP7_75t_L g1422 ( .A(n_824), .Y(n_1422) );
OAI221xp5_ASAP7_75t_L g1391 ( .A1(n_828), .A2(n_948), .B1(n_1361), .B2(n_1363), .C(n_1392), .Y(n_1391) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_835), .B2(n_836), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_833), .A2(n_1014), .B1(n_1326), .B2(n_1327), .Y(n_1325) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g892 ( .A(n_842), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_844), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1225) );
INVx1_ASAP7_75t_L g905 ( .A(n_849), .Y(n_905) );
NAND4xp75_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .C(n_878), .D(n_898), .Y(n_849) );
OAI31xp33_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_865), .A3(n_875), .B(n_876), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g1366 ( .A1(n_854), .A2(n_872), .B1(n_1367), .B2(n_1368), .C(n_1369), .Y(n_1366) );
OAI21xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B(n_862), .Y(n_858) );
INVx2_ASAP7_75t_SL g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g872 ( .A(n_861), .Y(n_872) );
INVx1_ASAP7_75t_L g1040 ( .A(n_861), .Y(n_1040) );
BUFx3_ASAP7_75t_L g1196 ( .A(n_863), .Y(n_1196) );
INVx2_ASAP7_75t_L g1204 ( .A(n_863), .Y(n_1204) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_863), .Y(n_1308) );
INVx1_ASAP7_75t_L g1476 ( .A(n_863), .Y(n_1476) );
OAI211xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_873), .C(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI31xp33_ASAP7_75t_SL g1088 ( .A1(n_877), .A2(n_1089), .A3(n_1092), .B(n_1103), .Y(n_1088) );
OAI31xp33_ASAP7_75t_L g1373 ( .A1(n_877), .A2(n_1374), .A3(n_1390), .B(n_1398), .Y(n_1373) );
AOI31xp33_ASAP7_75t_SL g1814 ( .A1(n_877), .A2(n_1815), .A3(n_1819), .B(n_1826), .Y(n_1814) );
AND2x2_ASAP7_75t_SL g878 ( .A(n_879), .B(n_897), .Y(n_878) );
AOI33xp33_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .A3(n_885), .B1(n_889), .B2(n_893), .B3(n_895), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g1797 ( .A1(n_880), .A2(n_1798), .B1(n_1803), .B2(n_1804), .Y(n_1797) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AND2x4_ASAP7_75t_L g914 ( .A(n_884), .B(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AND2x4_ASAP7_75t_L g921 ( .A(n_892), .B(n_915), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g1416 ( .A(n_895), .B(n_1417), .C(n_1418), .Y(n_1416) );
INVx2_ASAP7_75t_SL g927 ( .A(n_896), .Y(n_927) );
INVx1_ASAP7_75t_L g1110 ( .A(n_896), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_1054), .B1(n_1123), .B2(n_1124), .Y(n_907) );
INVx1_ASAP7_75t_L g1123 ( .A(n_908), .Y(n_1123) );
XNOR2x1_ASAP7_75t_L g908 ( .A(n_909), .B(n_996), .Y(n_908) );
INVx1_ASAP7_75t_L g994 ( .A(n_910), .Y(n_994) );
NAND4xp25_ASAP7_75t_L g910 ( .A(n_911), .B(n_950), .C(n_957), .D(n_980), .Y(n_910) );
INVx8_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_917) );
INVx3_ASAP7_75t_L g1090 ( .A(n_919), .Y(n_1090) );
INVx3_ASAP7_75t_L g1348 ( .A(n_919), .Y(n_1348) );
INVx3_ASAP7_75t_L g1091 ( .A(n_921), .Y(n_1091) );
INVx3_ASAP7_75t_L g1323 ( .A(n_921), .Y(n_1323) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_925), .B(n_928), .Y(n_922) );
BUFx3_ASAP7_75t_L g1264 ( .A(n_924), .Y(n_1264) );
INVx1_ASAP7_75t_L g1109 ( .A(n_926), .Y(n_1109) );
INVx1_ASAP7_75t_L g1341 ( .A(n_927), .Y(n_1341) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g955 ( .A(n_931), .Y(n_955) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
CKINVDCx11_ASAP7_75t_R g1115 ( .A(n_933), .Y(n_1115) );
CKINVDCx6p67_ASAP7_75t_R g935 ( .A(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_940), .B1(n_941), .B2(n_942), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_938), .A2(n_1000), .B1(n_1001), .B2(n_1002), .Y(n_999) );
BUFx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx2_ASAP7_75t_L g1147 ( .A(n_939), .Y(n_1147) );
INVx3_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_952), .B(n_1058), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_952), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1343 ( .A(n_954), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .Y(n_954) );
BUFx2_ASAP7_75t_L g1383 ( .A(n_956), .Y(n_1383) );
NOR3xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_965), .C(n_976), .Y(n_957) );
INVx2_ASAP7_75t_L g1086 ( .A(n_959), .Y(n_1086) );
INVx1_ASAP7_75t_L g1319 ( .A(n_959), .Y(n_1319) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_959), .Y(n_1372) );
NAND2x1p5_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
INVx2_ASAP7_75t_SL g961 ( .A(n_962), .Y(n_961) );
OR2x6_ASAP7_75t_L g963 ( .A(n_962), .B(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g979 ( .A(n_962), .Y(n_979) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_962), .B(n_964), .Y(n_1087) );
INVx2_ASAP7_75t_L g1317 ( .A(n_963), .Y(n_1317) );
OAI22xp5_ASAP7_75t_SL g965 ( .A1(n_966), .A2(n_968), .B1(n_970), .B2(n_972), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_970), .A2(n_1061), .B1(n_1065), .B2(n_1076), .Y(n_1060) );
INVx1_ASAP7_75t_L g1315 ( .A(n_970), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_970), .A2(n_1063), .B1(n_1359), .B2(n_1366), .Y(n_1358) );
INVx4_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_976), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1316 ( .A1(n_976), .A2(n_1317), .B1(n_1318), .B2(n_1319), .C(n_1320), .Y(n_1316) );
AND2x2_ASAP7_75t_L g976 ( .A(n_977), .B(n_979), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_986), .B1(n_987), .B2(n_988), .C(n_989), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_981), .A2(n_1334), .B1(n_1339), .B2(n_1352), .Y(n_1351) );
AND2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_982), .A2(n_1009), .B1(n_1011), .B2(n_1028), .Y(n_1027) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx2_ASAP7_75t_SL g1277 ( .A(n_983), .Y(n_1277) );
INVx1_ASAP7_75t_L g1821 ( .A(n_983), .Y(n_1821) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
OR2x6_ASAP7_75t_L g990 ( .A(n_985), .B(n_991), .Y(n_990) );
OR2x6_ASAP7_75t_L g992 ( .A(n_985), .B(n_993), .Y(n_992) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_985), .B(n_1121), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1403 ( .A(n_985), .B(n_991), .Y(n_1403) );
CKINVDCx6p67_ASAP7_75t_R g1350 ( .A(n_990), .Y(n_1350) );
INVx2_ASAP7_75t_L g1082 ( .A(n_991), .Y(n_1082) );
CKINVDCx6p67_ASAP7_75t_R g1352 ( .A(n_992), .Y(n_1352) );
INVx1_ASAP7_75t_L g1079 ( .A(n_993), .Y(n_1079) );
OAI21xp33_ASAP7_75t_L g1428 ( .A1(n_993), .A2(n_1429), .B(n_1430), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1573 ( .A1(n_995), .A2(n_1553), .B1(n_1558), .B2(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_SL g1053 ( .A(n_997), .Y(n_1053) );
NAND4xp75_ASAP7_75t_L g997 ( .A(n_998), .B(n_1018), .C(n_1023), .D(n_1049), .Y(n_997) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_1006), .A2(n_1040), .B(n_1041), .C(n_1043), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1012), .B1(n_1013), .B2(n_1014), .Y(n_1010) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
NOR2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1022), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1039), .Y(n_1030) );
OAI211xp5_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1033), .B(n_1036), .C(n_1037), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1033), .A2(n_1066), .B1(n_1250), .B2(n_1252), .C(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
NAND2xp33_ASAP7_75t_L g1441 ( .A(n_1035), .B(n_1442), .Y(n_1441) );
BUFx2_ASAP7_75t_L g1362 ( .A(n_1040), .Y(n_1362) );
INVxp67_ASAP7_75t_SL g1124 ( .A(n_1054), .Y(n_1124) );
XNOR2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
AND4x1_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1059), .C(n_1088), .D(n_1117), .Y(n_1056) );
NOR3xp33_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1083), .C(n_1084), .Y(n_1059) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g1306 ( .A(n_1063), .Y(n_1306) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1064), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B1(n_1068), .B2(n_1071), .C(n_1072), .Y(n_1065) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1309 ( .A(n_1082), .Y(n_1309) );
NOR3xp33_ASAP7_75t_L g1357 ( .A(n_1083), .B(n_1358), .C(n_1371), .Y(n_1357) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_1094), .A2(n_1329), .B1(n_1330), .B2(n_1331), .C(n_1332), .Y(n_1328) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_1100), .A2(n_1145), .B1(n_1146), .B2(n_1148), .Y(n_1144) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_1113), .A2(n_1115), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .Y(n_1117) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
XNOR2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1298), .Y(n_1126) );
AO22x2_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1129), .B1(n_1241), .B2(n_1242), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
XNOR2xp5_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1185), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1152), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1136), .Y(n_1133) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
AOI21xp5_ASAP7_75t_SL g1152 ( .A1(n_1153), .A2(n_1179), .B(n_1180), .Y(n_1152) );
NAND4xp25_ASAP7_75t_SL g1153 ( .A(n_1154), .B(n_1162), .C(n_1167), .D(n_1169), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1826 ( .A1(n_1155), .A2(n_1803), .B1(n_1827), .B2(n_1828), .Y(n_1826) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1360 ( .A(n_1164), .Y(n_1360) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1166), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1172), .B1(n_1173), .B2(n_1175), .C(n_1176), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
XNOR2x1_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1240), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1214), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1189), .B1(n_1212), .B2(n_1213), .Y(n_1187) );
OAI31xp33_ASAP7_75t_SL g1424 ( .A1(n_1188), .A2(n_1425), .A3(n_1426), .B(n_1427), .Y(n_1424) );
NAND3xp33_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1201), .C(n_1209), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_1198), .A2(n_1211), .B1(n_1234), .B2(n_1237), .Y(n_1233) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1206), .Y(n_1508) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1206), .Y(n_1822) );
NOR3xp33_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1223), .C(n_1224), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1220), .Y(n_1215) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_1236), .A2(n_1412), .B1(n_1413), .B2(n_1414), .C(n_1415), .Y(n_1411) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
XOR2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1297), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1269), .Y(n_1243) );
AND4x1_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1248), .C(n_1251), .D(n_1255), .Y(n_1244) );
AOI33xp33_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1258), .A3(n_1263), .B1(n_1266), .B2(n_1267), .B3(n_1268), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
BUFx3_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AOI21xp5_ASAP7_75t_L g1269 ( .A1(n_1270), .A2(n_1271), .B(n_1272), .Y(n_1269) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1279), .Y(n_1293) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
HB1xp67_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1446), .B2(n_1447), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
XNOR2x1_ASAP7_75t_SL g1300 ( .A(n_1301), .B(n_1353), .Y(n_1300) );
BUFx2_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
NAND4xp75_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1321), .C(n_1349), .D(n_1351), .Y(n_1303) );
AND2x2_ASAP7_75t_SL g1304 ( .A(n_1305), .B(n_1316), .Y(n_1304) );
AOI33xp33_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .A3(n_1310), .B1(n_1313), .B2(n_1314), .B3(n_1315), .Y(n_1305) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
OAI221xp5_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1328), .B1(n_1333), .B2(n_1338), .C(n_1342), .Y(n_1324) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
AOI21xp5_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1344), .B(n_1345), .Y(n_1342) );
AO22x2_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1355), .B1(n_1405), .B2(n_1406), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
AND4x1_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1373), .C(n_1399), .D(n_1401), .Y(n_1356) );
OAI221xp5_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1361), .B1(n_1362), .B2(n_1363), .C(n_1364), .Y(n_1359) );
OAI221xp5_ASAP7_75t_L g1375 ( .A1(n_1376), .A2(n_1377), .B1(n_1378), .B2(n_1381), .C(n_1382), .Y(n_1375) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx2_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1397), .Y(n_1464) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1404), .Y(n_1401) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
NAND3xp33_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1420), .C(n_1424), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1419), .Y(n_1409) );
NOR2xp33_ASAP7_75t_SL g1420 ( .A(n_1421), .B(n_1423), .Y(n_1420) );
OAI211xp5_ASAP7_75t_SL g1427 ( .A1(n_1428), .A2(n_1431), .B(n_1435), .C(n_1439), .Y(n_1427) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVxp67_ASAP7_75t_SL g1446 ( .A(n_1447), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1449), .B1(n_1490), .B2(n_1534), .Y(n_1447) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1467), .Y(n_1450) );
AND4x1_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1455), .C(n_1458), .D(n_1461), .Y(n_1451) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1490), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1515), .Y(n_1493) );
NAND3xp33_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1505), .C(n_1511), .Y(n_1495) );
NOR3xp33_ASAP7_75t_SL g1515 ( .A(n_1516), .B(n_1521), .C(n_1523), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1519), .Y(n_1516) );
OAI221xp5_ASAP7_75t_SL g1535 ( .A1(n_1536), .A2(n_1697), .B1(n_1789), .B2(n_1833), .C(n_1839), .Y(n_1535) );
NOR3xp33_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1700), .C(n_1746), .Y(n_1536) );
AOI21xp5_ASAP7_75t_L g1537 ( .A1(n_1538), .A2(n_1651), .B(n_1690), .Y(n_1537) );
AOI221xp5_ASAP7_75t_L g1538 ( .A1(n_1539), .A2(n_1584), .B1(n_1600), .B2(n_1606), .C(n_1614), .Y(n_1538) );
INVxp67_ASAP7_75t_SL g1539 ( .A(n_1540), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1560), .Y(n_1540) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1541), .Y(n_1672) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1541), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1719 ( .A(n_1541), .B(n_1703), .Y(n_1719) );
HB1xp67_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
INVx2_ASAP7_75t_SL g1604 ( .A(n_1542), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1542), .B(n_1597), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1542), .B(n_1597), .Y(n_1656) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1543), .Y(n_1594) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1543), .Y(n_1693) );
AND2x4_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1547), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1544), .B(n_1547), .Y(n_1571) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
AND2x4_ASAP7_75t_L g1549 ( .A(n_1545), .B(n_1547), .Y(n_1549) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1546), .B(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1548), .Y(n_1556) );
INVx1_ASAP7_75t_SL g1579 ( .A(n_1549), .Y(n_1579) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1549), .Y(n_1612) );
OAI22xp33_ASAP7_75t_L g1550 ( .A1(n_1551), .A2(n_1552), .B1(n_1557), .B2(n_1558), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1581 ( .A1(n_1552), .A2(n_1558), .B1(n_1582), .B2(n_1583), .Y(n_1581) );
OAI22xp33_ASAP7_75t_L g1587 ( .A1(n_1552), .A2(n_1588), .B1(n_1589), .B2(n_1590), .Y(n_1587) );
BUFx3_ASAP7_75t_L g1697 ( .A(n_1552), .Y(n_1697) );
BUFx6f_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
OR2x2_ASAP7_75t_L g1558 ( .A(n_1554), .B(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1554), .Y(n_1567) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1555), .Y(n_1566) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1558), .Y(n_1591) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1559), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1575), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1561), .B(n_1607), .Y(n_1674) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_1561), .B(n_1641), .Y(n_1686) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
NOR2xp33_ASAP7_75t_L g1633 ( .A(n_1562), .B(n_1618), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1722 ( .A(n_1562), .B(n_1575), .Y(n_1722) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1562), .B(n_1608), .Y(n_1771) );
OR2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1572), .Y(n_1562) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1563), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1563), .B(n_1575), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1563), .B(n_1639), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1563), .B(n_1572), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1570), .Y(n_1563) );
AND2x4_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1567), .Y(n_1565) );
OAI21xp33_ASAP7_75t_SL g1850 ( .A1(n_1566), .A2(n_1848), .B(n_1851), .Y(n_1850) );
AND2x4_ASAP7_75t_L g1568 ( .A(n_1567), .B(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1571), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1572), .B(n_1607), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1572), .B(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1572), .Y(n_1639) );
NOR2xp33_ASAP7_75t_L g1752 ( .A(n_1572), .B(n_1613), .Y(n_1752) );
CKINVDCx6p67_ASAP7_75t_R g1613 ( .A(n_1575), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1575), .B(n_1633), .Y(n_1632) );
OAI331xp33_ASAP7_75t_L g1652 ( .A1(n_1575), .A2(n_1639), .A3(n_1653), .B1(n_1657), .B2(n_1660), .B3(n_1662), .C1(n_1664), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1575), .B(n_1638), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1575), .B(n_1620), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1575), .B(n_1621), .Y(n_1735) );
OR2x2_ASAP7_75t_L g1742 ( .A(n_1575), .B(n_1621), .Y(n_1742) );
OR2x6_ASAP7_75t_SL g1575 ( .A(n_1576), .B(n_1581), .Y(n_1575) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_1577), .A2(n_1578), .B1(n_1579), .B2(n_1580), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g1592 ( .A1(n_1579), .A2(n_1593), .B1(n_1594), .B2(n_1595), .Y(n_1592) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1584), .Y(n_1675) );
A2O1A1Ixp33_ASAP7_75t_SL g1778 ( .A1(n_1584), .A2(n_1761), .B(n_1779), .C(n_1780), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1585), .B(n_1596), .Y(n_1584) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1585), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1585), .B(n_1628), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1666 ( .A(n_1585), .B(n_1597), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1585), .B(n_1597), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1585), .B(n_1649), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1585), .B(n_1604), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_1585), .B(n_1690), .Y(n_1737) );
INVx3_ASAP7_75t_L g1766 ( .A(n_1585), .Y(n_1766) );
INVx3_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1586), .B(n_1597), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1586), .B(n_1608), .Y(n_1663) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1586), .B(n_1656), .Y(n_1787) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1592), .Y(n_1586) );
HB1xp67_ASAP7_75t_L g1699 ( .A(n_1590), .Y(n_1699) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
OAI211xp5_ASAP7_75t_SL g1614 ( .A1(n_1596), .A2(n_1615), .B(n_1622), .C(n_1644), .Y(n_1614) );
AOI22xp33_ASAP7_75t_SL g1755 ( .A1(n_1596), .A2(n_1721), .B1(n_1756), .B2(n_1760), .Y(n_1755) );
O2A1O1Ixp33_ASAP7_75t_L g1760 ( .A1(n_1596), .A2(n_1618), .B(n_1649), .C(n_1705), .Y(n_1760) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1597), .B(n_1604), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1597), .B(n_1604), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1706 ( .A1(n_1597), .A2(n_1642), .B1(n_1707), .B2(n_1709), .Y(n_1706) );
AND2x4_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1599), .Y(n_1597) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1605), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1602), .B(n_1704), .Y(n_1777) );
INVx2_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
OR2x2_ASAP7_75t_L g1768 ( .A(n_1603), .B(n_1704), .Y(n_1768) );
INVx2_ASAP7_75t_SL g1628 ( .A(n_1604), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1605), .B(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_1607), .B(n_1620), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1607), .B(n_1679), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1613), .Y(n_1607) );
INVx4_ASAP7_75t_L g1618 ( .A(n_1608), .Y(n_1618) );
INVx2_ASAP7_75t_L g1625 ( .A(n_1608), .Y(n_1625) );
NOR2xp33_ASAP7_75t_L g1641 ( .A(n_1608), .B(n_1613), .Y(n_1641) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1608), .B(n_1679), .Y(n_1711) );
OR2x2_ASAP7_75t_L g1721 ( .A(n_1608), .B(n_1722), .Y(n_1721) );
AOI322xp5_ASAP7_75t_L g1725 ( .A1(n_1608), .A2(n_1649), .A3(n_1655), .B1(n_1661), .B2(n_1726), .C1(n_1729), .C2(n_1731), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1608), .B(n_1661), .Y(n_1754) );
AND2x6_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1610), .Y(n_1608) );
INVx2_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
OAI22xp5_ASAP7_75t_L g1691 ( .A1(n_1612), .A2(n_1692), .B1(n_1693), .B2(n_1694), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1613), .B(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1613), .B(n_1638), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1613), .B(n_1678), .Y(n_1677) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_1613), .B(n_1711), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1613), .B(n_1639), .Y(n_1757) );
OR2x2_ASAP7_75t_L g1782 ( .A(n_1613), .B(n_1639), .Y(n_1782) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1619), .Y(n_1617) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1618), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1618), .B(n_1655), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1618), .B(n_1650), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1618), .B(n_1679), .Y(n_1678) );
NOR2xp33_ASAP7_75t_L g1758 ( .A(n_1618), .B(n_1759), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1619), .B(n_1646), .Y(n_1724) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1620), .Y(n_1659) );
OAI22xp5_ASAP7_75t_SL g1773 ( .A1(n_1621), .A2(n_1774), .B1(n_1775), .B2(n_1777), .Y(n_1773) );
AOI211xp5_ASAP7_75t_L g1622 ( .A1(n_1623), .A2(n_1627), .B(n_1630), .C(n_1634), .Y(n_1622) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1625), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1744 ( .A(n_1625), .B(n_1745), .Y(n_1744) );
OAI32xp33_ASAP7_75t_L g1756 ( .A1(n_1625), .A2(n_1649), .A3(n_1705), .B1(n_1757), .B2(n_1758), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1628), .Y(n_1631) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1628), .Y(n_1646) );
NOR2xp33_ASAP7_75t_L g1733 ( .A(n_1628), .B(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1628), .Y(n_1745) );
OAI22xp5_ASAP7_75t_L g1769 ( .A1(n_1628), .A2(n_1705), .B1(n_1770), .B2(n_1772), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1770 ( .A(n_1628), .B(n_1771), .Y(n_1770) );
OAI21xp33_ASAP7_75t_L g1717 ( .A1(n_1629), .A2(n_1718), .B(n_1720), .Y(n_1717) );
NOR2xp33_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1632), .Y(n_1630) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1632), .Y(n_1714) );
AOI21xp33_ASAP7_75t_SL g1634 ( .A1(n_1635), .A2(n_1636), .B(n_1642), .Y(n_1634) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1635), .Y(n_1772) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1636), .Y(n_1738) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1640), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1637), .B(n_1659), .Y(n_1658) );
NOR2xp33_ASAP7_75t_L g1680 ( .A(n_1637), .B(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NOR3xp33_ASAP7_75t_L g1784 ( .A(n_1639), .B(n_1704), .C(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
OAI21xp5_ASAP7_75t_L g1644 ( .A1(n_1645), .A2(n_1647), .B(n_1650), .Y(n_1644) );
AOI221xp5_ASAP7_75t_SL g1732 ( .A1(n_1645), .A2(n_1733), .B1(n_1736), .B2(n_1738), .C(n_1739), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1649), .Y(n_1647) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1650), .Y(n_1728) );
NOR5xp2_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1668), .C(n_1680), .D(n_1683), .E(n_1687), .Y(n_1651) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
A2O1A1Ixp33_ASAP7_75t_L g1788 ( .A1(n_1654), .A2(n_1687), .B(n_1752), .C(n_1766), .Y(n_1788) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
NOR2xp33_ASAP7_75t_L g1687 ( .A(n_1656), .B(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
NOR2x1_ASAP7_75t_R g1716 ( .A(n_1659), .B(n_1704), .Y(n_1716) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1661), .B(n_1685), .Y(n_1684) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1661), .B(n_1689), .Y(n_1749) );
INVxp67_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1667), .Y(n_1664) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
OAI22xp5_ASAP7_75t_SL g1668 ( .A1(n_1669), .A2(n_1671), .B1(n_1675), .B2(n_1676), .Y(n_1668) );
AOI21xp33_ASAP7_75t_L g1739 ( .A1(n_1669), .A2(n_1737), .B(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1670), .B(n_1781), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1673), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1672), .B(n_1730), .Y(n_1774) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1707 ( .A(n_1674), .B(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
AOI21xp33_ASAP7_75t_L g1712 ( .A1(n_1681), .A2(n_1713), .B(n_1715), .Y(n_1712) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1690), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1765 ( .A(n_1690), .B(n_1766), .Y(n_1765) );
CKINVDCx5p33_ASAP7_75t_R g1785 ( .A(n_1690), .Y(n_1785) );
OR2x6_ASAP7_75t_SL g1690 ( .A(n_1691), .B(n_1695), .Y(n_1690) );
OAI22xp5_ASAP7_75t_L g1695 ( .A1(n_1696), .A2(n_1697), .B1(n_1698), .B2(n_1699), .Y(n_1695) );
NAND4xp25_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1717), .C(n_1725), .D(n_1732), .Y(n_1700) );
AOI211xp5_ASAP7_75t_SL g1701 ( .A1(n_1702), .A2(n_1703), .B(n_1706), .C(n_1712), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1705), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1704), .B(n_1735), .Y(n_1734) );
NOR2x1_ASAP7_75t_L g1781 ( .A(n_1704), .B(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1705), .Y(n_1727) );
OAI31xp33_ASAP7_75t_L g1783 ( .A1(n_1705), .A2(n_1731), .A3(n_1784), .B(n_1786), .Y(n_1783) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1711), .Y(n_1779) );
INVxp67_ASAP7_75t_SL g1713 ( .A(n_1714), .Y(n_1713) );
INVxp33_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
NAND2xp33_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1723), .Y(n_1720) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1721), .Y(n_1731) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1722), .Y(n_1776) );
INVxp33_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1728), .Y(n_1726) );
NOR2xp33_ASAP7_75t_L g1775 ( .A(n_1729), .B(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
AOI22xp5_ASAP7_75t_L g1763 ( .A1(n_1736), .A2(n_1764), .B1(n_1767), .B2(n_1773), .Y(n_1763) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1743), .Y(n_1740) );
OAI21xp5_ASAP7_75t_SL g1767 ( .A1(n_1741), .A2(n_1768), .B(n_1769), .Y(n_1767) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
NAND5xp2_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1763), .C(n_1778), .D(n_1783), .E(n_1788), .Y(n_1746) );
OAI31xp33_ASAP7_75t_SL g1747 ( .A1(n_1748), .A2(n_1750), .A3(n_1755), .B(n_1761), .Y(n_1747) );
INVxp67_ASAP7_75t_SL g1748 ( .A(n_1749), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1750 ( .A(n_1751), .B(n_1753), .Y(n_1750) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1757), .Y(n_1759) );
CKINVDCx14_ASAP7_75t_R g1761 ( .A(n_1762), .Y(n_1761) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
NAND2xp5_ASAP7_75t_SL g1791 ( .A(n_1792), .B(n_1829), .Y(n_1791) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1793), .Y(n_1831) );
NAND3xp33_ASAP7_75t_SL g1793 ( .A(n_1794), .B(n_1797), .C(n_1805), .Y(n_1793) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1814), .Y(n_1830) );
NAND3xp33_ASAP7_75t_L g1829 ( .A(n_1830), .B(n_1831), .C(n_1832), .Y(n_1829) );
NAND2xp5_ASAP7_75t_L g1843 ( .A(n_1830), .B(n_1831), .Y(n_1843) );
CKINVDCx14_ASAP7_75t_R g1833 ( .A(n_1834), .Y(n_1833) );
INVx4_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
INVxp33_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
CKINVDCx5p33_ASAP7_75t_R g1846 ( .A(n_1847), .Y(n_1846) );
HB1xp67_ASAP7_75t_L g1849 ( .A(n_1850), .Y(n_1849) );
endmodule