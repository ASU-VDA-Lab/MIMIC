module fake_jpeg_25492_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_36),
.B(n_35),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_68),
.B1(n_24),
.B2(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_54),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_36),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_55),
.B(n_59),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_65),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_70),
.B1(n_81),
.B2(n_20),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_20),
.B(n_22),
.C(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_86),
.B1(n_97),
.B2(n_113),
.Y(n_134)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_63),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_29),
.B1(n_22),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_77),
.B1(n_80),
.B2(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_28),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_78),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_31),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_24),
.B1(n_32),
.B2(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_131),
.Y(n_143)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_80),
.B1(n_60),
.B2(n_66),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_139),
.B1(n_87),
.B2(n_104),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_13),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_106),
.B(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2x1_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_145),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_88),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_116),
.C(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_161),
.B1(n_135),
.B2(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_107),
.B1(n_97),
.B2(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_91),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_151),
.B(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_92),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_169),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_174),
.B(n_181),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_126),
.A3(n_118),
.B1(n_108),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_14),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_134),
.B1(n_125),
.B2(n_127),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_178),
.B1(n_186),
.B2(n_159),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_127),
.B1(n_138),
.B2(n_121),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_109),
.B(n_102),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_148),
.B(n_165),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_121),
.B(n_110),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_12),
.C(n_16),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_2),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_123),
.B1(n_115),
.B2(n_95),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_142),
.B1(n_153),
.B2(n_149),
.C(n_143),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_192),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_150),
.C(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_176),
.C(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_145),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_156),
.B(n_123),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_179),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_170),
.CI(n_173),
.CON(n_212),
.SN(n_212)
);

OAI321xp33_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_156),
.A3(n_115),
.B1(n_32),
.B2(n_17),
.C(n_8),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_203),
.A3(n_180),
.B1(n_4),
.B2(n_6),
.C(n_9),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_156),
.A3(n_32),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_169),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_195),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_193),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_203),
.A3(n_184),
.B(n_9),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_176),
.C(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_193),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_167),
.C(n_186),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_192),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_199),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_213),
.B1(n_189),
.B2(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_204),
.B1(n_4),
.B2(n_10),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_210),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_216),
.B(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

NAND4xp25_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_207),
.C(n_209),
.D(n_210),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_2),
.C(n_10),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_2),
.C(n_10),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_226),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_237),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_235),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_234),
.B(n_225),
.Y(n_241)
);


endmodule