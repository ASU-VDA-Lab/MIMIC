module real_jpeg_11486_n_16 (n_5, n_4, n_8, n_0, n_12, n_384, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_384;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_45),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_3),
.B(n_67),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_3),
.B(n_61),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_35),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_4),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_54),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_4),
.B(n_61),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_35),
.Y(n_166)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_7),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_28),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_45),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_61),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_35),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_8),
.B(n_69),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_54),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_12),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_67),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_12),
.B(n_45),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_69),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_13),
.B(n_61),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_45),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_13),
.B(n_67),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_13),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_13),
.B(n_35),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_13),
.B(n_54),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_13),
.B(n_40),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_40),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_67),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_14),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_14),
.B(n_28),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_14),
.B(n_61),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_14),
.B(n_54),
.Y(n_315)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_54),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_45),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_28),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_149),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_20),
.B(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_98),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_21),
.B(n_82),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_23),
.B(n_49),
.C(n_57),
.Y(n_147)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.C(n_43),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_25),
.A2(n_26),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.C(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_27),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_27),
.B(n_121),
.C(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_27),
.A2(n_113),
.B1(n_121),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_27),
.A2(n_113),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_27),
.B(n_194),
.Y(n_210)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_29),
.A2(n_30),
.B1(n_68),
.B2(n_71),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_29),
.B(n_68),
.C(n_304),
.Y(n_323)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_39),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_SL g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_32),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_32),
.B(n_79),
.Y(n_320)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_34),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_34),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_34),
.A2(n_111),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_37),
.A2(n_43),
.B1(n_44),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_39),
.B(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_39),
.B(n_233),
.Y(n_304)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_66),
.C(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_43),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_43),
.A2(n_44),
.B1(n_123),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_43),
.A2(n_44),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_120),
.C(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_44),
.B(n_214),
.Y(n_268)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_46),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_46),
.B(n_233),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_51),
.B(n_53),
.C(n_55),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_54),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_73),
.C(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_59),
.A2(n_60),
.B1(n_107),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_107),
.C(n_108),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_66),
.C(n_68),
.Y(n_129)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_65),
.A2(n_66),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_66),
.B(n_254),
.C(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_68),
.A2(n_71),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx5_ASAP7_75t_SL g202 ( 
.A(n_69),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_77),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_75),
.B(n_192),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_78),
.B(n_190),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_81),
.A2(n_87),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_81),
.B(n_142),
.C(n_316),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.C(n_93),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_88),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.C(n_92),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_90),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_91),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_91),
.B(n_202),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_93),
.A2(n_94),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_115),
.C(n_119),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_99),
.A2(n_100),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_109),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_102),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_107),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_108),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_121),
.A2(n_164),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_121),
.B(n_261),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_147),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_145),
.B2(n_146),
.Y(n_125)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_141),
.A2(n_142),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_176),
.B(n_380),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_174),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_151),
.B(n_174),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_167),
.C(n_171),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_152),
.B(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.C(n_161),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_153),
.A2(n_154),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_158),
.B(n_161),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_162),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_165),
.A2(n_166),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_165),
.Y(n_353)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_166),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_167),
.B(n_171),
.Y(n_373)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_360),
.A3(n_370),
.B1(n_374),
.B2(n_379),
.C(n_384),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_307),
.C(n_355),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_278),
.B(n_306),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_248),
.B(n_277),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_217),
.B(n_247),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_196),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_182),
.B(n_196),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_193),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_199),
.B1(n_200),
.B2(n_208),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_244),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.CI(n_186),
.CON(n_183),
.SN(n_183)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_209),
.B2(n_216),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_208),
.C(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_204),
.C(n_207),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_214),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_214),
.A2(n_215),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_214),
.B(n_328),
.C(n_331),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_241),
.B(n_246),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_230),
.B(n_240),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_228),
.C(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_235),
.B(n_239),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_250),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_263),
.B2(n_264),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_265),
.C(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_259),
.C(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_275),
.B2(n_276),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_274),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_279),
.B(n_280),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_296),
.B2(n_305),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_295),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_295),
.C(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_293),
.C(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_287),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.CI(n_290),
.CON(n_287),
.SN(n_287)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_296),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.CI(n_302),
.CON(n_296),
.SN(n_296)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_298),
.C(n_302),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B(n_301),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_301),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_308),
.A2(n_376),
.B(n_377),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_337),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_337),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_325),
.C(n_336),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_324),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_317),
.C(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_321),
.C(n_323),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_326),
.B1(n_336),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_332),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_333),
.C(n_335),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_330),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_354),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_346),
.C(n_354),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_344),
.C(n_345),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_349),
.C(n_350),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_375),
.B(n_378),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_362),
.B(n_363),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_366),
.C(n_369),
.Y(n_371)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_372),
.Y(n_379)
);


endmodule