module fake_jpeg_2737_n_83 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_24),
.Y(n_39)
);

NAND2x1p5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_28),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_26),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_32),
.B(n_28),
.Y(n_47)
);

XNOR2x1_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_35),
.B1(n_33),
.B2(n_26),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_51),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_35),
.C(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_41),
.C(n_42),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_66),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_10),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_8),
.B(n_18),
.C(n_17),
.D(n_16),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_20),
.B(n_12),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_70),
.A3(n_67),
.B1(n_68),
.B2(n_66),
.C1(n_65),
.C2(n_3),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_73),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_76),
.B(n_72),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_4),
.Y(n_80)
);

XOR2x2_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_5),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_6),
.C(n_7),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_6),
.Y(n_83)
);


endmodule