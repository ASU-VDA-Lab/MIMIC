module real_jpeg_24013_n_26 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_147, n_24, n_146, n_6, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_155, n_26);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_147;
input n_24;
input n_146;
input n_6;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_26;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_2),
.B(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_3),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_5),
.B(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_6),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_9),
.B(n_78),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_11),
.B(n_48),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_12),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_13),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.C(n_123),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_15),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_16),
.B(n_98),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_17),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_18),
.B(n_41),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_21),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_21),
.B(n_109),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_22),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_23),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_140),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_39),
.B(n_137),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_30),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_35),
.B(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_37),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_37),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_37),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_37),
.B(n_143),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_38),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_136),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_130),
.B(n_135),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_125),
.B(n_129),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_122),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_116),
.B(n_121),
.Y(n_50)
);

OAI321xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_108),
.A3(n_111),
.B1(n_114),
.B2(n_115),
.C(n_146),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_102),
.B(n_107),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_97),
.B(n_101),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_89),
.B(n_96),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_88),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_81),
.B(n_87),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_77),
.B(n_80),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_70),
.B(n_76),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_120),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_134),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_141),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_147),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_148),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_149),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_150),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_151),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_152),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_153),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_154),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_155),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_156),
.Y(n_113)
);


endmodule