module fake_netlist_1_11715_n_37 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g14 ( .A(n_1), .B(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_7), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_2), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_13), .B(n_11), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_8), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_17), .B(n_0), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_12), .B(n_9), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
OAI21xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_20), .B(n_14), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_19), .B(n_18), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AND3x1_ASAP7_75t_L g27 ( .A(n_26), .B(n_15), .C(n_24), .Y(n_27) );
OAI31xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_14), .A3(n_25), .B(n_2), .Y(n_28) );
NOR2xp33_ASAP7_75t_L g29 ( .A(n_27), .B(n_26), .Y(n_29) );
AOI321xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_14), .A3(n_1), .B1(n_3), .B2(n_4), .C(n_5), .Y(n_30) );
NOR2x1_ASAP7_75t_L g31 ( .A(n_28), .B(n_26), .Y(n_31) );
NOR3xp33_ASAP7_75t_L g32 ( .A(n_31), .B(n_16), .C(n_3), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_16), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
NAND3xp33_ASAP7_75t_L g35 ( .A(n_33), .B(n_17), .C(n_23), .Y(n_35) );
OAI221xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_17), .B1(n_23), .B2(n_0), .C(n_4), .Y(n_36) );
NAND2x1p5_ASAP7_75t_L g37 ( .A(n_36), .B(n_35), .Y(n_37) );
endmodule