module real_aes_6282_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_800;
wire n_1170;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_673;
wire n_1067;
wire n_518;
wire n_905;
wire n_792;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1123;
wire n_549;
wire n_571;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_448;
wire n_545;
wire n_556;
wire n_752;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_1160;
wire n_550;
wire n_966;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_994;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_1182;
wire n_872;
wire n_1053;
wire n_976;
wire n_636;
wire n_477;
wire n_906;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_817;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_1100;
wire n_1174;
wire n_1167;
wire n_1193;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_1142;
wire n_508;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_869;
wire n_613;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_1179;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_1187;
wire n_1028;
wire n_1000;
wire n_533;
wire n_1003;
wire n_727;
wire n_1083;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_968;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_926;
wire n_679;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_1071;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_1191;
wire n_705;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_1190;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_1045;
wire n_837;
wire n_871;
wire n_1159;
wire n_474;
wire n_1156;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_652;
wire n_703;
wire n_1040;
wire n_601;
wire n_500;
wire n_1185;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g1078 ( .A(n_0), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_1), .A2(n_179), .B1(n_545), .B2(n_548), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_2), .A2(n_183), .B1(n_609), .B2(n_682), .Y(n_1114) );
INVx1_ASAP7_75t_L g765 ( .A(n_3), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_4), .A2(n_365), .B1(n_469), .B2(n_830), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_5), .A2(n_144), .B1(n_548), .B2(n_827), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_6), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g1173 ( .A(n_7), .Y(n_1173) );
AOI222xp33_ASAP7_75t_L g876 ( .A1(n_8), .A2(n_209), .B1(n_316), .B2(n_489), .C1(n_496), .C2(n_560), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_9), .A2(n_110), .B1(n_547), .B2(n_848), .Y(n_1029) );
AO22x2_ASAP7_75t_L g430 ( .A1(n_10), .A2(n_239), .B1(n_422), .B2(n_427), .Y(n_430) );
INVx1_ASAP7_75t_L g1135 ( .A(n_10), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_11), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_12), .A2(n_167), .B1(n_442), .B2(n_473), .Y(n_822) );
AOI222xp33_ASAP7_75t_L g949 ( .A1(n_13), .A2(n_340), .B1(n_350), .B2(n_488), .C1(n_642), .C2(n_950), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_14), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_15), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_16), .Y(n_975) );
INVx1_ASAP7_75t_L g815 ( .A(n_17), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_18), .A2(n_59), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_19), .A2(n_138), .B1(n_553), .B2(n_628), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_20), .A2(n_127), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_21), .A2(n_218), .B1(n_527), .B2(n_932), .C(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g800 ( .A(n_22), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_23), .A2(n_299), .B1(n_488), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g804 ( .A(n_24), .Y(n_804) );
INVx1_ASAP7_75t_L g1061 ( .A(n_25), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_26), .A2(n_333), .B1(n_468), .B2(n_471), .Y(n_467) );
AOI22xp5_ASAP7_75t_SL g838 ( .A1(n_27), .A2(n_212), .B1(n_682), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_28), .A2(n_275), .B1(n_446), .B2(n_531), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_29), .A2(n_102), .B1(n_488), .B2(n_642), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_30), .A2(n_228), .B1(n_441), .B2(n_446), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_31), .A2(n_213), .B1(n_559), .B2(n_561), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_32), .A2(n_118), .B1(n_593), .B2(n_842), .C(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_33), .A2(n_171), .B1(n_676), .B2(n_930), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_34), .A2(n_1166), .B1(n_1190), .B2(n_1191), .Y(n_1165) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_34), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_35), .A2(n_120), .B1(n_526), .B2(n_687), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_36), .Y(n_997) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_37), .A2(n_148), .B1(n_529), .B2(n_1032), .Y(n_1031) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_38), .A2(n_92), .B1(n_543), .B2(n_618), .Y(n_671) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_39), .A2(n_125), .B1(n_422), .B2(n_423), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_40), .A2(n_284), .B1(n_442), .B2(n_589), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_41), .A2(n_265), .B1(n_543), .B2(n_548), .Y(n_1144) );
AOI222xp33_ASAP7_75t_L g832 ( .A1(n_42), .A2(n_211), .B1(n_315), .B2(n_561), .C1(n_618), .C2(n_666), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_43), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_44), .B(n_1028), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_45), .A2(n_329), .B1(n_435), .B2(n_1158), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_46), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_47), .A2(n_84), .B1(n_471), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_48), .A2(n_274), .B1(n_757), .B2(n_930), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_49), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_50), .A2(n_225), .B1(n_616), .B2(n_673), .C(n_872), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_51), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_52), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_53), .A2(n_128), .B1(n_593), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_54), .A2(n_381), .B1(n_676), .B2(n_677), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_55), .A2(n_194), .B1(n_471), .B2(n_1037), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_56), .A2(n_87), .B1(n_967), .B2(n_969), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_57), .B(n_578), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_58), .Y(n_466) );
INVx1_ASAP7_75t_L g793 ( .A(n_60), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_61), .A2(n_155), .B1(n_526), .B2(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g624 ( .A(n_62), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g1188 ( .A1(n_63), .A2(n_176), .B1(n_311), .B2(n_559), .C1(n_560), .C2(n_1189), .Y(n_1188) );
AOI22x1_ASAP7_75t_L g702 ( .A1(n_64), .A2(n_703), .B1(n_730), .B2(n_731), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_64), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_65), .A2(n_95), .B1(n_441), .B2(n_682), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_66), .A2(n_114), .B1(n_435), .B2(n_586), .Y(n_1109) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_67), .A2(n_131), .B1(n_685), .B2(n_686), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_68), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_69), .A2(n_245), .B1(n_589), .B2(n_631), .Y(n_779) );
AO22x1_ASAP7_75t_L g986 ( .A1(n_70), .A2(n_987), .B1(n_1014), .B2(n_1015), .Y(n_986) );
INVx1_ASAP7_75t_L g1014 ( .A(n_70), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_71), .A2(n_104), .B1(n_754), .B2(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_72), .A2(n_328), .B1(n_452), .B2(n_631), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_73), .Y(n_973) );
INVx1_ASAP7_75t_L g869 ( .A(n_74), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_75), .A2(n_204), .B1(n_543), .B2(n_547), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_76), .A2(n_384), .B1(n_941), .B2(n_969), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_77), .B(n_536), .Y(n_944) );
INVx1_ASAP7_75t_L g900 ( .A(n_78), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_79), .A2(n_396), .B1(n_842), .B2(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_80), .A2(n_244), .B1(n_435), .B2(n_899), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g1172 ( .A(n_81), .Y(n_1172) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_82), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_83), .A2(n_347), .B1(n_1086), .B2(n_1111), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_85), .A2(n_390), .B1(n_543), .B2(n_618), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g1052 ( .A(n_86), .Y(n_1052) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_88), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_89), .A2(n_221), .B1(n_782), .B2(n_1086), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_90), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_91), .A2(n_272), .B1(n_593), .B2(n_777), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_93), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_94), .A2(n_220), .B1(n_441), .B2(n_446), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g866 ( .A1(n_96), .A2(n_116), .B1(n_452), .B2(n_471), .C(n_867), .Y(n_866) );
AO22x2_ASAP7_75t_L g426 ( .A1(n_97), .A2(n_273), .B1(n_422), .B2(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g1132 ( .A(n_97), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_98), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_99), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_100), .A2(n_160), .B1(n_848), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_101), .A2(n_250), .B1(n_468), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_103), .A2(n_236), .B1(n_848), .B2(n_849), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_105), .A2(n_295), .B1(n_454), .B2(n_631), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_106), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_107), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_108), .A2(n_287), .B1(n_545), .B2(n_559), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_109), .A2(n_206), .B1(n_535), .B2(n_539), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_111), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_112), .A2(n_387), .B1(n_489), .B2(n_827), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_113), .A2(n_1139), .B1(n_1159), .B2(n_1160), .Y(n_1138) );
CKINVDCx20_ASAP7_75t_R g1159 ( .A(n_113), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_115), .A2(n_277), .B1(n_435), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g873 ( .A(n_117), .Y(n_873) );
XOR2x2_ASAP7_75t_L g911 ( .A(n_119), .B(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g851 ( .A(n_121), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_122), .A2(n_293), .B1(n_651), .B2(n_678), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_123), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_124), .A2(n_281), .B1(n_474), .B2(n_830), .Y(n_837) );
INVx1_ASAP7_75t_L g1136 ( .A(n_125), .Y(n_1136) );
CKINVDCx20_ASAP7_75t_R g1183 ( .A(n_126), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_129), .A2(n_276), .B1(n_710), .B2(n_711), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_130), .A2(n_318), .B1(n_710), .B2(n_842), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_132), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_133), .Y(n_724) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_134), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_135), .B(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_136), .A2(n_291), .B1(n_757), .B2(n_758), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g990 ( .A(n_137), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_139), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_140), .A2(n_162), .B1(n_447), .B2(n_681), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g1170 ( .A(n_141), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_142), .B(n_922), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_143), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_145), .A2(n_364), .B1(n_454), .B2(n_469), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_146), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_147), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_149), .A2(n_154), .B1(n_651), .B2(n_678), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_150), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_151), .A2(n_859), .B1(n_877), .B2(n_878), .Y(n_858) );
INVx1_ASAP7_75t_L g877 ( .A(n_151), .Y(n_877) );
OAI22xp5_ASAP7_75t_SL g1066 ( .A1(n_152), .A2(n_1067), .B1(n_1068), .B2(n_1088), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_152), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_153), .Y(n_1001) );
INVx1_ASAP7_75t_L g868 ( .A(n_156), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_157), .A2(n_362), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_158), .A2(n_243), .B1(n_658), .B2(n_1111), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_159), .A2(n_178), .B1(n_462), .B2(n_1086), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_161), .A2(n_376), .B1(n_689), .B2(n_932), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_163), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_164), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_165), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_166), .A2(n_219), .B1(n_559), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_168), .A2(n_319), .B1(n_553), .B2(n_687), .Y(n_939) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_169), .A2(n_356), .B1(n_689), .B2(n_691), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_170), .A2(n_264), .B1(n_531), .B2(n_754), .Y(n_753) );
AND2x6_ASAP7_75t_L g401 ( .A(n_172), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_172), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_173), .A2(n_298), .B1(n_532), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_174), .A2(n_346), .B1(n_489), .B2(n_561), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_175), .A2(n_278), .B1(n_578), .B2(n_811), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_177), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_180), .A2(n_349), .B1(n_682), .B2(n_796), .Y(n_795) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_181), .A2(n_254), .B1(n_271), .B2(n_489), .C1(n_497), .C2(n_578), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_182), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_184), .A2(n_327), .B1(n_526), .B2(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g633 ( .A(n_185), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_186), .A2(n_353), .B1(n_714), .B2(n_758), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_187), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_188), .A2(n_377), .B1(n_681), .B2(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g1013 ( .A(n_189), .Y(n_1013) );
INVx1_ASAP7_75t_L g814 ( .A(n_190), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g1169 ( .A(n_191), .Y(n_1169) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_192), .A2(n_332), .B1(n_527), .B2(n_758), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_193), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_195), .A2(n_268), .B1(n_441), .B2(n_446), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_196), .Y(n_1179) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_197), .A2(n_260), .B1(n_556), .B2(n_609), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_198), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_199), .A2(n_367), .B1(n_678), .B2(n_775), .Y(n_1060) );
AO22x2_ASAP7_75t_L g421 ( .A1(n_200), .A2(n_261), .B1(n_422), .B2(n_423), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_200), .B(n_1134), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_201), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_202), .A2(n_233), .B1(n_463), .B2(n_532), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_203), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_205), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_207), .A2(n_386), .B1(n_555), .B2(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g1023 ( .A(n_208), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_210), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_214), .B(n_502), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_215), .A2(n_266), .B1(n_551), .B2(n_553), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_216), .Y(n_1072) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_217), .A2(n_359), .B1(n_680), .B2(n_682), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_222), .A2(n_292), .B1(n_616), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_223), .A2(n_323), .B1(n_539), .B2(n_846), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_224), .Y(n_833) );
OA22x2_ASAP7_75t_L g789 ( .A1(n_226), .A2(n_790), .B1(n_791), .B2(n_817), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_226), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_227), .A2(n_313), .B1(n_526), .B2(n_586), .C(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g626 ( .A(n_229), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g1153 ( .A(n_230), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_231), .B(n_846), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_232), .B(n_669), .Y(n_977) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_234), .A2(n_399), .B(n_407), .C(n_1137), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_235), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_237), .B(n_539), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_238), .A2(n_258), .B1(n_502), .B2(n_547), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_240), .A2(n_331), .B1(n_548), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_241), .A2(n_297), .B1(n_529), .B2(n_777), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_242), .A2(n_314), .B1(n_543), .B2(n_648), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_246), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_247), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_248), .Y(n_980) );
INVx1_ASAP7_75t_L g621 ( .A(n_249), .Y(n_621) );
INVx1_ASAP7_75t_L g875 ( .A(n_251), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_252), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g1187 ( .A(n_253), .Y(n_1187) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_255), .A2(n_366), .B1(n_378), .B2(n_497), .C1(n_559), .C2(n_560), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_256), .Y(n_958) );
INVx2_ASAP7_75t_L g406 ( .A(n_257), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_259), .A2(n_294), .B1(n_502), .B2(n_918), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g1147 ( .A(n_262), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_263), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_267), .A2(n_735), .B1(n_736), .B2(n_760), .Y(n_734) );
CKINVDCx14_ASAP7_75t_R g760 ( .A(n_267), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_269), .A2(n_317), .B1(n_561), .B2(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_270), .Y(n_573) );
INVx1_ASAP7_75t_L g1053 ( .A(n_279), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_280), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_282), .A2(n_305), .B1(n_685), .B2(n_758), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_283), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_285), .A2(n_563), .B1(n_596), .B2(n_597), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_285), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_286), .Y(n_741) );
INVx1_ASAP7_75t_L g794 ( .A(n_288), .Y(n_794) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_289), .A2(n_394), .B1(n_473), .B2(n_658), .Y(n_657) );
XOR2x2_ASAP7_75t_L g1018 ( .A(n_290), .B(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g422 ( .A(n_296), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_296), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g1152 ( .A(n_300), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_301), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_302), .A2(n_383), .B1(n_441), .B2(n_446), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_303), .A2(n_354), .B1(n_656), .B2(n_757), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_304), .B(n_536), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_306), .Y(n_1097) );
INVx1_ASAP7_75t_L g865 ( .A(n_307), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g1184 ( .A1(n_308), .A2(n_358), .B1(n_535), .B2(n_673), .C(n_1185), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_309), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g816 ( .A(n_310), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_312), .A2(n_414), .B1(n_519), .B2(n_520), .Y(n_413) );
INVx1_ASAP7_75t_L g519 ( .A(n_312), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_320), .Y(n_477) );
INVx1_ASAP7_75t_L g806 ( .A(n_321), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g1103 ( .A(n_322), .Y(n_1103) );
INVx1_ASAP7_75t_L g1011 ( .A(n_324), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_325), .B(n_616), .Y(n_770) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_326), .A2(n_661), .B1(n_662), .B2(n_693), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_326), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_330), .A2(n_392), .B1(n_536), .B2(n_541), .Y(n_825) );
AND2x2_ASAP7_75t_L g405 ( .A(n_334), .B(n_406), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_335), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_336), .B(n_577), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_337), .Y(n_1099) );
INVx1_ASAP7_75t_L g402 ( .A(n_338), .Y(n_402) );
INVx1_ASAP7_75t_L g854 ( .A(n_339), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_341), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_342), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_343), .A2(n_348), .B1(n_435), .B2(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g1049 ( .A(n_344), .Y(n_1049) );
INVx1_ASAP7_75t_L g629 ( .A(n_345), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_351), .Y(n_1105) );
INVx1_ASAP7_75t_L g862 ( .A(n_352), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_355), .Y(n_992) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_357), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_360), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_361), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_363), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g1181 ( .A(n_368), .Y(n_1181) );
INVx1_ASAP7_75t_L g612 ( .A(n_369), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_370), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_371), .B(n_769), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_372), .B(n_560), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_373), .A2(n_389), .B1(n_551), .B2(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_374), .B(n_539), .Y(n_645) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_375), .B(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_379), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_380), .B(n_615), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_382), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_385), .Y(n_1186) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_388), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_391), .A2(n_1092), .B1(n_1115), .B2(n_1116), .Y(n_1091) );
INVx1_ASAP7_75t_L g1115 ( .A(n_391), .Y(n_1115) );
INVx1_ASAP7_75t_L g801 ( .A(n_393), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_395), .A2(n_955), .B1(n_981), .B2(n_982), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_395), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_397), .Y(n_1047) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_402), .Y(n_1128) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_403), .A2(n_1127), .B(n_1197), .Y(n_1196) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_697), .B1(n_1122), .B2(n_1123), .C(n_1124), .Y(n_407) );
INVx1_ASAP7_75t_L g1123 ( .A(n_408), .Y(n_1123) );
AOI22xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_410), .B1(n_601), .B2(n_696), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_521), .B2(n_600), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g520 ( .A(n_414), .Y(n_520) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_475), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_450), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_433), .B1(n_434), .B2(n_439), .C(n_440), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_417), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_417), .A2(n_1181), .B1(n_1182), .B2(n_1183), .Y(n_1180) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g622 ( .A(n_418), .Y(n_622) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_428), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_420), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g552 ( .A(n_420), .B(n_428), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g864 ( .A(n_420), .B(n_445), .Y(n_864) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_425), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_421), .B(n_426), .Y(n_438) );
INVx2_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
AND2x2_ASAP7_75t_L g493 ( .A(n_421), .B(n_430), .Y(n_493) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_424), .Y(n_427) );
INVx1_ASAP7_75t_L g518 ( .A(n_425), .Y(n_518) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
AND2x2_ASAP7_75t_L g465 ( .A(n_426), .B(n_458), .Y(n_465) );
INVx1_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
AND2x4_ASAP7_75t_L g436 ( .A(n_428), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g464 ( .A(n_428), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g470 ( .A(n_428), .B(n_457), .Y(n_470) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x2_ASAP7_75t_L g445 ( .A(n_429), .B(n_432), .Y(n_445) );
OR2x2_ASAP7_75t_L g456 ( .A(n_429), .B(n_432), .Y(n_456) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g498 ( .A(n_430), .B(n_432), .Y(n_498) );
AND2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g511 ( .A(n_431), .Y(n_511) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_435), .Y(n_711) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g553 ( .A(n_436), .Y(n_553) );
BUFx2_ASAP7_75t_SL g656 ( .A(n_436), .Y(n_656) );
BUFx3_ASAP7_75t_L g692 ( .A(n_436), .Y(n_692) );
BUFx2_ASAP7_75t_SL g758 ( .A(n_436), .Y(n_758) );
BUFx2_ASAP7_75t_L g775 ( .A(n_436), .Y(n_775) );
BUFx3_ASAP7_75t_L g932 ( .A(n_436), .Y(n_932) );
AND2x2_ASAP7_75t_L g777 ( .A(n_437), .B(n_511), .Y(n_777) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x6_ASAP7_75t_L g448 ( .A(n_438), .B(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_442), .Y(n_531) );
INVx5_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g610 ( .A(n_443), .Y(n_610) );
INVx2_ASAP7_75t_L g681 ( .A(n_443), .Y(n_681) );
INVx4_ASAP7_75t_L g798 ( .A(n_443), .Y(n_798) );
INVx3_ASAP7_75t_L g941 ( .A(n_443), .Y(n_941) );
INVx1_ASAP7_75t_L g968 ( .A(n_443), .Y(n_968) );
INVx8_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g474 ( .A(n_445), .B(n_457), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_445), .B(n_465), .Y(n_485) );
AND2x6_ASAP7_75t_L g541 ( .A(n_445), .B(n_465), .Y(n_541) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g532 ( .A(n_447), .Y(n_532) );
BUFx2_ASAP7_75t_L g682 ( .A(n_447), .Y(n_682) );
BUFx2_ASAP7_75t_L g754 ( .A(n_447), .Y(n_754) );
BUFx4f_ASAP7_75t_SL g1008 ( .A(n_447), .Y(n_1008) );
INVx6_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_448), .A2(n_862), .B1(n_863), .B2(n_865), .Y(n_861) );
INVx1_ASAP7_75t_SL g969 ( .A(n_448), .Y(n_969) );
INVx1_ASAP7_75t_L g546 ( .A(n_449), .Y(n_546) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_460), .B1(n_461), .B2(n_466), .C(n_467), .Y(n_450) );
OAI221xp5_ASAP7_75t_SL g1151 ( .A1(n_451), .A2(n_528), .B1(n_1152), .B2(n_1153), .C(n_1154), .Y(n_1151) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g555 ( .A(n_453), .Y(n_555) );
INVx2_ASAP7_75t_L g710 ( .A(n_453), .Y(n_710) );
INVx2_ASAP7_75t_SL g930 ( .A(n_453), .Y(n_930) );
INVx11_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx11_ASAP7_75t_L g590 ( .A(n_454), .Y(n_590) );
AND2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
AND2x4_ASAP7_75t_L g538 ( .A(n_455), .B(n_465), .Y(n_538) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g480 ( .A(n_456), .B(n_481), .Y(n_480) );
AND2x6_ASAP7_75t_L g497 ( .A(n_457), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_461), .A2(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
INVx2_ASAP7_75t_L g594 ( .A(n_464), .Y(n_594) );
BUFx3_ASAP7_75t_L g678 ( .A(n_464), .Y(n_678) );
BUFx3_ASAP7_75t_L g782 ( .A(n_464), .Y(n_782) );
INVx1_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g706 ( .A(n_469), .Y(n_706) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_469), .Y(n_842) );
BUFx3_ASAP7_75t_L g1086 ( .A(n_469), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_SL g526 ( .A(n_470), .Y(n_526) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_470), .Y(n_651) );
INVx2_ASAP7_75t_L g690 ( .A(n_470), .Y(n_690) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx6_ASAP7_75t_L g557 ( .A(n_474), .Y(n_557) );
BUFx3_ASAP7_75t_L g676 ( .A(n_474), .Y(n_676) );
BUFx3_ASAP7_75t_L g899 ( .A(n_474), .Y(n_899) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .C(n_506), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_482), .B2(n_483), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_478), .A2(n_566), .B1(n_567), .B2(n_568), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_478), .A2(n_483), .B1(n_720), .B2(n_721), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_478), .A2(n_804), .B1(n_805), .B2(n_806), .C(n_807), .Y(n_803) );
OAI221xp5_ASAP7_75t_SL g1141 ( .A1(n_478), .A2(n_805), .B1(n_1142), .B2(n_1143), .C(n_1144), .Y(n_1141) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g740 ( .A(n_479), .Y(n_740) );
INVx1_ASAP7_75t_SL g991 ( .A(n_479), .Y(n_991) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_480), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g1096 ( .A(n_480), .Y(n_1096) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g805 ( .A(n_484), .Y(n_805) );
INVx1_ASAP7_75t_SL g993 ( .A(n_484), .Y(n_993) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g570 ( .A(n_485), .Y(n_570) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_494), .B1(n_495), .B2(n_499), .C1(n_500), .C2(n_505), .Y(n_486) );
OAI221xp5_ASAP7_75t_SL g1073 ( .A1(n_487), .A2(n_1022), .B1(n_1074), .B2(n_1075), .C(n_1076), .Y(n_1073) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g996 ( .A(n_488), .Y(n_996) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx4f_ASAP7_75t_SL g559 ( .A(n_490), .Y(n_559) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_490), .Y(n_813) );
BUFx2_ASAP7_75t_L g853 ( .A(n_490), .Y(n_853) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_490), .Y(n_926) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g504 ( .A(n_492), .Y(n_504) );
AND2x4_ASAP7_75t_L g503 ( .A(n_493), .B(n_504), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_493), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g545 ( .A(n_493), .B(n_546), .Y(n_545) );
OAI222xp33_ASAP7_75t_L g722 ( .A1(n_495), .A2(n_574), .B1(n_723), .B2(n_724), .C1(n_725), .C2(n_726), .Y(n_722) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g572 ( .A(n_496), .Y(n_572) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx3_ASAP7_75t_L g666 ( .A(n_497), .Y(n_666) );
INVx4_ASAP7_75t_L g744 ( .A(n_497), .Y(n_744) );
INVx2_ASAP7_75t_L g885 ( .A(n_497), .Y(n_885) );
INVx2_ASAP7_75t_SL g915 ( .A(n_497), .Y(n_915) );
INVx1_ASAP7_75t_L g516 ( .A(n_498), .Y(n_516) );
AND2x4_ASAP7_75t_L g548 ( .A(n_498), .B(n_518), .Y(n_548) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g669 ( .A(n_502), .Y(n_669) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx12f_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_512), .B2(n_513), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_508), .A2(n_513), .B1(n_728), .B2(n_729), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_508), .A2(n_513), .B1(n_979), .B2(n_980), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_508), .A2(n_1000), .B1(n_1001), .B2(n_1002), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_508), .A2(n_1106), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_SL g1104 ( .A(n_509), .Y(n_1104) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_510), .Y(n_581) );
BUFx3_ASAP7_75t_L g874 ( .A(n_510), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_513), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_579) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g1002 ( .A(n_514), .Y(n_1002) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_515), .A2(n_581), .B1(n_748), .B2(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_515), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_515), .A2(n_874), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_515), .Y(n_1106) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
OA22x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_562), .B1(n_598), .B2(n_599), .Y(n_521) );
INVx1_ASAP7_75t_L g599 ( .A(n_522), .Y(n_599) );
NAND4xp75_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .C(n_549), .D(n_558), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
INVx1_ASAP7_75t_L g1182 ( .A(n_526), .Y(n_1182) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g607 ( .A(n_528), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g792 ( .A1(n_528), .A2(n_706), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_792) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_SL g533 ( .A(n_534), .B(n_542), .Y(n_533) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_536), .Y(n_922) );
INVx5_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g616 ( .A(n_537), .Y(n_616) );
INVx2_ASAP7_75t_L g846 ( .A(n_537), .Y(n_846) );
INVx2_ASAP7_75t_L g1028 ( .A(n_537), .Y(n_1028) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_SL g673 ( .A(n_540), .Y(n_673) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
BUFx4f_ASAP7_75t_L g769 ( .A(n_541), .Y(n_769) );
BUFx2_ASAP7_75t_L g924 ( .A(n_541), .Y(n_924) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g808 ( .A(n_544), .Y(n_808) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g827 ( .A(n_545), .Y(n_827) );
BUFx2_ASAP7_75t_L g848 ( .A(n_545), .Y(n_848) );
BUFx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
BUFx2_ASAP7_75t_SL g648 ( .A(n_548), .Y(n_648) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_548), .Y(n_849) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
INVx1_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_551), .Y(n_1158) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
BUFx3_ASAP7_75t_L g687 ( .A(n_552), .Y(n_687) );
BUFx3_ASAP7_75t_L g830 ( .A(n_552), .Y(n_830) );
INVxp67_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g631 ( .A(n_557), .Y(n_631) );
INVx2_ASAP7_75t_L g714 ( .A(n_557), .Y(n_714) );
INVx2_ASAP7_75t_L g1111 ( .A(n_557), .Y(n_1111) );
INVx1_ASAP7_75t_L g574 ( .A(n_559), .Y(n_574) );
INVx1_ASAP7_75t_L g725 ( .A(n_560), .Y(n_725) );
BUFx4f_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
INVx1_ASAP7_75t_L g598 ( .A(n_562), .Y(n_598) );
INVx2_ASAP7_75t_L g597 ( .A(n_563), .Y(n_597) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_583), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_571), .C(n_579), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_568), .A2(n_991), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g613 ( .A(n_570), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_574), .B2(n_575), .C(n_576), .Y(n_571) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_572), .A2(n_640), .B(n_641), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g974 ( .A1(n_574), .A2(n_915), .B1(n_975), .B2(n_976), .C(n_977), .Y(n_974) );
OAI221xp5_ASAP7_75t_SL g1098 ( .A1(n_574), .A2(n_743), .B1(n_1099), .B2(n_1100), .C(n_1101), .Y(n_1098) );
BUFx4f_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_591), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g628 ( .A(n_590), .Y(n_628) );
INVx2_ASAP7_75t_SL g658 ( .A(n_590), .Y(n_658) );
INVx4_ASAP7_75t_L g685 ( .A(n_590), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_590), .A2(n_713), .B1(n_800), .B2(n_801), .C(n_802), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g696 ( .A(n_601), .Y(n_696) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_634), .B1(n_635), .B2(n_695), .Y(n_602) );
INVx2_ASAP7_75t_L g695 ( .A(n_603), .Y(n_695) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_633), .Y(n_603) );
NAND4xp75_ASAP7_75t_L g604 ( .A(n_605), .B(n_611), .C(n_619), .D(n_632), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OA211x2_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_614), .C(n_617), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_613), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_738) );
OA211x2_ASAP7_75t_L g942 ( .A1(n_613), .A2(n_943), .B(n_944), .C(n_945), .Y(n_942) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_625), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g712 ( .A1(n_622), .A2(n_713), .B1(n_715), .B2(n_716), .C(n_717), .Y(n_712) );
OAI221xp5_ASAP7_75t_SL g962 ( .A1(n_622), .A2(n_963), .B1(n_964), .B2(n_965), .C(n_966), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_623), .A2(n_959), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_629), .B2(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_659), .B1(n_660), .B2(n_694), .Y(n_635) );
INVx1_ASAP7_75t_L g694 ( .A(n_636), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_649), .C(n_653), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_644), .Y(n_638) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .C(n_647), .Y(n_644) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
BUFx4f_ASAP7_75t_SL g757 ( .A(n_655), .Y(n_757) );
INVx1_ASAP7_75t_SL g870 ( .A(n_656), .Y(n_870) );
INVx1_ASAP7_75t_L g1178 ( .A(n_658), .Y(n_1178) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g693 ( .A(n_662), .Y(n_693) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_674), .C(n_683), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_670), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_667), .B(n_668), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g764 ( .A1(n_665), .A2(n_765), .B(n_766), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g994 ( .A1(n_665), .A2(n_995), .B1(n_996), .B2(n_997), .C(n_998), .Y(n_994) );
OAI21xp33_ASAP7_75t_L g1048 ( .A1(n_665), .A2(n_1049), .B(n_1050), .Y(n_1048) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g963 ( .A(n_676), .Y(n_963) );
INVx1_ASAP7_75t_L g959 ( .A(n_677), .Y(n_959) );
BUFx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g1174 ( .A(n_682), .Y(n_1174) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g1012 ( .A(n_685), .Y(n_1012) );
BUFx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g781 ( .A(n_690), .Y(n_781) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g1122 ( .A(n_697), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_905), .B2(n_1121), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
XNOR2xp5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_786), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_732), .B2(n_733), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g731 ( .A(n_703), .Y(n_731) );
AND2x2_ASAP7_75t_SL g703 ( .A(n_704), .B(n_718), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_712), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g957 ( .A1(n_706), .A2(n_958), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_713), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_713), .A2(n_1177), .B1(n_1178), .B2(n_1179), .Y(n_1176) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_722), .C(n_727), .Y(n_718) );
OAI222xp33_ASAP7_75t_L g809 ( .A1(n_725), .A2(n_744), .B1(n_810), .B2(n_814), .C1(n_815), .C2(n_816), .Y(n_809) );
OAI222xp33_ASAP7_75t_L g1145 ( .A1(n_725), .A2(n_1022), .B1(n_1146), .B2(n_1147), .C1(n_1148), .C2(n_1149), .Y(n_1145) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
AO22x1_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_761), .B1(n_784), .B2(n_785), .Y(n_733) );
INVx1_ASAP7_75t_L g785 ( .A(n_734), .Y(n_785) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_750), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .C(n_747), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_740), .A2(n_805), .B1(n_972), .B2(n_973), .Y(n_971) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_745), .B(n_746), .Y(n_742) );
OAI21xp5_ASAP7_75t_SL g850 ( .A1(n_743), .A2(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g1189 ( .A(n_743), .Y(n_1189) );
BUFx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx4_ASAP7_75t_L g950 ( .A(n_744), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_755), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
INVx3_ASAP7_75t_SL g784 ( .A(n_761), .Y(n_784) );
AO22x1_ASAP7_75t_L g1118 ( .A1(n_761), .A2(n_784), .B1(n_1040), .B2(n_1041), .Y(n_1118) );
XOR2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_783), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_763), .B(n_772), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_770), .C(n_771), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_778), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_857), .B2(n_904), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_818), .B1(n_855), .B2(n_856), .Y(n_788) );
INVx1_ASAP7_75t_L g855 ( .A(n_789), .Y(n_855) );
INVx1_ASAP7_75t_L g817 ( .A(n_791), .Y(n_817) );
OR4x1_ASAP7_75t_L g791 ( .A(n_792), .B(n_799), .C(n_803), .D(n_809), .Y(n_791) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_798), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_805), .A2(n_1045), .B1(n_1046), .B2(n_1047), .Y(n_1044) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx4_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g856 ( .A(n_818), .Y(n_856) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_834), .Y(n_818) );
XOR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_833), .Y(n_819) );
NAND4xp75_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_828), .D(n_832), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
AND2x2_ASAP7_75t_SL g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g1038 ( .A(n_830), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_834), .A2(n_881), .B1(n_901), .B2(n_902), .Y(n_880) );
INVx2_ASAP7_75t_SL g901 ( .A(n_834), .Y(n_901) );
XOR2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_854), .Y(n_834) );
NOR4xp75_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .C(n_844), .D(n_850), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NAND2x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
NAND2xp5_ASAP7_75t_SL g844 ( .A(n_845), .B(n_847), .Y(n_844) );
INVx1_ASAP7_75t_SL g919 ( .A(n_849), .Y(n_919) );
INVx2_ASAP7_75t_SL g904 ( .A(n_857), .Y(n_904) );
OA22x2_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_879), .B1(n_880), .B2(n_903), .Y(n_857) );
INVx1_ASAP7_75t_L g903 ( .A(n_858), .Y(n_903) );
INVx1_ASAP7_75t_L g878 ( .A(n_859), .Y(n_878) );
AND4x1_ASAP7_75t_L g859 ( .A(n_860), .B(n_866), .C(n_871), .D(n_876), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_863), .A2(n_1005), .B1(n_1006), .B2(n_1007), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_863), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
BUFx2_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_874), .A2(n_1002), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g902 ( .A(n_881), .Y(n_902) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_900), .Y(n_881) );
NAND2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_892), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_888), .Y(n_883) );
OAI21xp5_ASAP7_75t_SL g884 ( .A1(n_885), .A2(n_886), .B(n_887), .Y(n_884) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .C(n_891), .Y(n_888) );
NOR2x1_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g1121 ( .A(n_905), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_907), .B1(n_1063), .B2(n_1120), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .B1(n_983), .B2(n_984), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
XNOR2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_954), .Y(n_909) );
AO22x2_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_936), .B1(n_952), .B2(n_953), .Y(n_910) );
INVx2_ASAP7_75t_L g952 ( .A(n_911), .Y(n_952) );
NAND2xp5_ASAP7_75t_SL g912 ( .A(n_913), .B(n_927), .Y(n_912) );
NOR2xp33_ASAP7_75t_SL g913 ( .A(n_914), .B(n_920), .Y(n_913) );
OAI21xp5_ASAP7_75t_SL g914 ( .A1(n_915), .A2(n_916), .B(n_917), .Y(n_914) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_923), .C(n_925), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g1146 ( .A(n_926), .Y(n_1146) );
NOR2x1_ASAP7_75t_L g927 ( .A(n_928), .B(n_933), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_931), .Y(n_928) );
INVx1_ASAP7_75t_L g1033 ( .A(n_930), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx3_ASAP7_75t_SL g953 ( .A(n_936), .Y(n_953) );
XOR2x2_ASAP7_75t_L g936 ( .A(n_937), .B(n_951), .Y(n_936) );
NAND4xp75_ASAP7_75t_L g937 ( .A(n_938), .B(n_942), .C(n_946), .D(n_949), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
INVx2_ASAP7_75t_L g1022 ( .A(n_950), .Y(n_1022) );
INVx2_ASAP7_75t_L g982 ( .A(n_955), .Y(n_982) );
AND2x2_ASAP7_75t_SL g955 ( .A(n_956), .B(n_970), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_962), .Y(n_956) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
NOR3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_974), .C(n_978), .Y(n_970) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B1(n_1016), .B2(n_1017), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1015 ( .A(n_987), .Y(n_1015) );
AND3x1_ASAP7_75t_L g987 ( .A(n_988), .B(n_1003), .C(n_1009), .Y(n_987) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_994), .C(n_999), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B1(n_992), .B2(n_993), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_993), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_1008), .Y(n_1007) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1040), .B1(n_1041), .B2(n_1062), .Y(n_1017) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1018), .Y(n_1062) );
NAND3x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1030), .C(n_1035), .Y(n_1019) );
NOR2x1_ASAP7_75t_SL g1020 ( .A(n_1021), .B(n_1025), .Y(n_1020) );
OAI21xp5_ASAP7_75t_SL g1021 ( .A1(n_1022), .A2(n_1023), .B(n_1024), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .C(n_1029), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1034), .Y(n_1030) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1039), .Y(n_1035) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_1041), .Y(n_1040) );
XOR2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1061), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1054), .Y(n_1042) );
NOR3xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1048), .C(n_1051), .Y(n_1043) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1058), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1063), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1065), .B1(n_1089), .B2(n_1119), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_SL g1067 ( .A(n_1068), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1080), .Y(n_1068) );
NOR3xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1073), .C(n_1077), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1084), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1087), .Y(n_1084) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1089), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B1(n_1117), .B2(n_1118), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1092), .Y(n_1116) );
AND2x2_ASAP7_75t_SL g1092 ( .A(n_1093), .B(n_1107), .Y(n_1092) );
NOR3xp33_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1098), .C(n_1102), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_1103), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1112), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_SL g1124 ( .A(n_1125), .Y(n_1124) );
NOR2x1_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1130), .Y(n_1125) );
OR2x2_ASAP7_75t_SL g1194 ( .A(n_1126), .B(n_1131), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1129), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1127), .B(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1128), .B(n_1162), .Y(n_1197) );
CKINVDCx16_ASAP7_75t_R g1162 ( .A(n_1129), .Y(n_1162) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
OAI222xp33_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1161), .B1(n_1163), .B2(n_1190), .C1(n_1192), .C2(n_1195), .Y(n_1137) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1139), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1150), .Y(n_1139) );
NOR2xp33_ASAP7_75t_SL g1140 ( .A(n_1141), .B(n_1145), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1155), .Y(n_1150) );
NAND2xp33_ASAP7_75t_SL g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1166), .Y(n_1191) );
AND4x1_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1175), .C(n_1184), .D(n_1188), .Y(n_1166) );
NOR2xp33_ASAP7_75t_SL g1167 ( .A(n_1168), .B(n_1171), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1180), .Y(n_1175) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_1193), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
CKINVDCx20_ASAP7_75t_R g1195 ( .A(n_1196), .Y(n_1195) );
endmodule