module fake_jpeg_15302_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_10),
.C(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_57),
.Y(n_82)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_29),
.B1(n_24),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_38),
.B1(n_49),
.B2(n_40),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_24),
.B1(n_29),
.B2(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_38),
.B1(n_29),
.B2(n_39),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_103),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_53),
.B1(n_28),
.B2(n_54),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_88),
.A3(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_41),
.B1(n_37),
.B2(n_28),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_41),
.B1(n_56),
.B2(n_28),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_97),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_37),
.B1(n_56),
.B2(n_23),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_57),
.B1(n_47),
.B2(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_105),
.Y(n_130)
);

AND2x4_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_48),
.B1(n_25),
.B2(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_108),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_114),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_125),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_45),
.B(n_71),
.C(n_32),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_79),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_151),
.C(n_50),
.Y(n_159)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_143),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_25),
.B(n_31),
.C(n_40),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_146),
.B(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_144),
.Y(n_158)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_63),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_30),
.Y(n_146)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_112),
.B1(n_107),
.B2(n_104),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_86),
.Y(n_151)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_131),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_84),
.B1(n_120),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_138),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_120),
.B1(n_117),
.B2(n_81),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_142),
.B1(n_148),
.B2(n_127),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_50),
.C(n_115),
.Y(n_166)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_132),
.Y(n_193)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_21),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_176),
.C(n_151),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_117),
.B1(n_81),
.B2(n_73),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_73),
.B1(n_109),
.B2(n_115),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_106),
.C(n_97),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_177),
.B(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_162),
.B(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_183),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_146),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_191),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_171),
.B1(n_142),
.B2(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_176),
.B1(n_160),
.B2(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_142),
.B1(n_140),
.B2(n_137),
.Y(n_220)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_150),
.B(n_130),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_141),
.B(n_27),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_161),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_172),
.B(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_145),
.C(n_144),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_199),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_173),
.B(n_170),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_201),
.B(n_217),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_170),
.B(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_164),
.B1(n_150),
.B2(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_216),
.B1(n_225),
.B2(n_23),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_195),
.B1(n_180),
.B2(n_181),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_132),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_221),
.C(n_33),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_223),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_196),
.B1(n_199),
.B2(n_198),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_167),
.B(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

AOI32xp33_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_182),
.A3(n_187),
.B1(n_177),
.B2(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_21),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_106),
.B1(n_42),
.B2(n_27),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_233),
.B1(n_235),
.B2(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_230),
.B(n_214),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_178),
.B1(n_192),
.B2(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_222),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_188),
.B1(n_136),
.B2(n_147),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_245),
.C(n_249),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_200),
.B1(n_203),
.B2(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_42),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_221),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_201),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_147),
.B1(n_124),
.B2(n_0),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_124),
.C(n_21),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_208),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_252),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_263),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_220),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_204),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_266),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_270),
.B(n_202),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_237),
.B(n_228),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_236),
.A2(n_207),
.B(n_203),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_36),
.B(n_35),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_233),
.B1(n_242),
.B2(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_276),
.B(n_265),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_277),
.B(n_258),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_241),
.C(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_280),
.C(n_290),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_249),
.C(n_224),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_225),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_202),
.B1(n_124),
.B2(n_0),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_292),
.B1(n_269),
.B2(n_266),
.Y(n_298)
);

AOI211xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_284),
.B(n_254),
.C(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_256),
.B(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_3),
.B(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_124),
.C(n_36),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_261),
.B(n_264),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_254),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_36),
.C(n_35),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_260),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_257),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_288),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_261),
.B1(n_271),
.B2(n_253),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_272),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_288),
.B(n_281),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_308),
.B1(n_293),
.B2(n_284),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_277),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_262),
.B1(n_272),
.B2(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_302),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_279),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_317),
.C(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_316),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_290),
.C(n_267),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_317),
.B1(n_321),
.B2(n_312),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_255),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_322),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_255),
.B1(n_8),
.B2(n_9),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_33),
.C(n_255),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_255),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_3),
.C(n_8),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_329),
.B(n_16),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_304),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_311),
.A2(n_296),
.B1(n_309),
.B2(n_11),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_333),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_13),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_314),
.B(n_13),
.Y(n_335)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_11),
.B(n_13),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_338),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_334),
.C(n_324),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_343),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_15),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_342),
.Y(n_348)
);

INVx11_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_15),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_344),
.B(n_347),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_336),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_345),
.A2(n_342),
.B1(n_343),
.B2(n_340),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g354 ( 
.A1(n_350),
.A2(n_351),
.B(n_346),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_345),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_348),
.B(n_349),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_354),
.C(n_19),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_355),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_19),
.C(n_17),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_358),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_18),
.C(n_19),
.Y(n_360)
);


endmodule