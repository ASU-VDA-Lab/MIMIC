module real_jpeg_33015_n_2 (n_1, n_0, n_2);

input n_1;
input n_0;

output n_2;

wire n_4;
wire n_3;

AND2x2_ASAP7_75t_L g2 ( 
.A(n_0),
.B(n_3),
.Y(n_2)
);

CKINVDCx5p33_ASAP7_75t_R g4 ( 
.A(n_1),
.Y(n_4)
);

CKINVDCx5p33_ASAP7_75t_R g3 ( 
.A(n_4),
.Y(n_3)
);


endmodule