module fake_jpeg_9151_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_54),
.Y(n_70)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_56),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_34),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_63),
.B1(n_30),
.B2(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_18),
.B1(n_33),
.B2(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_1),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_74),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_73),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_93),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_2),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_2),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_46),
.B1(n_48),
.B2(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_34),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_48),
.B1(n_51),
.B2(n_62),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_115),
.B1(n_122),
.B2(n_90),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_39),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_106),
.C(n_110),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_102),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_58),
.B(n_30),
.C(n_29),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_107),
.B(n_73),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_58),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_38),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_58),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_38),
.C(n_31),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_14),
.B(n_15),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_31),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_93),
.C(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_48),
.B1(n_66),
.B2(n_44),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_73),
.B1(n_88),
.B2(n_53),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_66),
.B1(n_65),
.B2(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_92),
.B1(n_78),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_109),
.B1(n_114),
.B2(n_120),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_116),
.C(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_74),
.B(n_69),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_146),
.B(n_149),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_74),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_142),
.B(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_29),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_76),
.B1(n_37),
.B2(n_65),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_28),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_69),
.B(n_73),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_97),
.B(n_15),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_107),
.B1(n_110),
.B2(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_88),
.B(n_31),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_44),
.B1(n_37),
.B2(n_36),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_119),
.B1(n_112),
.B2(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_158),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_168),
.B1(n_146),
.B2(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_165),
.C(n_124),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_162),
.B1(n_134),
.B2(n_143),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_164),
.B(n_166),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_119),
.B1(n_103),
.B2(n_112),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_103),
.B(n_113),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_19),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_108),
.B(n_27),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_108),
.B(n_27),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_174),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_53),
.C(n_76),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_27),
.C(n_20),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_202),
.Y(n_232)
);

XNOR2x2_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_144),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_194),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_186),
.B(n_188),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_139),
.B1(n_147),
.B2(n_132),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_206),
.B1(n_155),
.B2(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_123),
.B1(n_142),
.B2(n_126),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_193),
.B1(n_176),
.B2(n_179),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_126),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_124),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.C(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_136),
.C(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_127),
.B1(n_140),
.B2(n_137),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_207),
.B1(n_157),
.B2(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_76),
.B1(n_37),
.B2(n_20),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_27),
.B1(n_20),
.B2(n_22),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_212),
.B1(n_206),
.B2(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_155),
.B1(n_154),
.B2(n_181),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_169),
.B(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_215),
.A2(n_217),
.B1(n_219),
.B2(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_226),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_169),
.B(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_196),
.C(n_159),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_170),
.B(n_171),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_178),
.C(n_172),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_176),
.C(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_167),
.B1(n_174),
.B2(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_175),
.B1(n_168),
.B2(n_22),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_234),
.C(n_193),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_191),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_233),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_246),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_232),
.Y(n_237)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_204),
.B1(n_200),
.B2(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_250),
.B1(n_213),
.B2(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_19),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_26),
.Y(n_271)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_185),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_211),
.A2(n_167),
.B1(n_207),
.B2(n_209),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_2),
.B(n_3),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_255),
.B(n_217),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_253),
.B1(n_31),
.B2(n_26),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_175),
.B1(n_22),
.B2(n_5),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_214),
.C(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_264),
.C(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_271),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_214),
.C(n_224),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_213),
.B1(n_227),
.B2(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_239),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_229),
.C(n_234),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_211),
.C(n_11),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_11),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_245),
.C(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_261),
.B1(n_269),
.B2(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_256),
.B1(n_263),
.B2(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_245),
.C(n_247),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_251),
.C(n_26),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_253),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_244),
.C(n_240),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_8),
.B1(n_13),
.B2(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_252),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_284),
.B(n_9),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_250),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_266),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_275),
.C(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_26),
.C(n_4),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_9),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_9),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_6),
.C(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_303),
.B(n_10),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_8),
.B(n_12),
.Y(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_304),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_290),
.C(n_3),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_7),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_10),
.B(n_14),
.C(n_3),
.D(n_4),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_285),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_310),
.B1(n_302),
.B2(n_297),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_309),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.C(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_311),
.B1(n_300),
.B2(n_4),
.Y(n_318)
);


endmodule