module real_jpeg_1022_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_249;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_185;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_98),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_47),
.B1(n_51),
.B2(n_98),
.Y(n_210)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_37),
.B1(n_39),
.B2(n_135),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_135),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_47),
.B1(n_51),
.B2(n_135),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_37),
.B1(n_39),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_4),
.A2(n_47),
.B1(n_51),
.B2(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_161),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_5),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_5),
.A2(n_26),
.B(n_170),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_65),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_39),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_47),
.C(n_50),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_206),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_5),
.B(n_88),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_45),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_58),
.Y(n_107)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_10),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_10),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_10),
.A2(n_29),
.B1(n_47),
.B2(n_51),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_37),
.B1(n_39),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_47),
.B1(n_51),
.B2(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_180),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_13),
.A2(n_47),
.B1(n_51),
.B2(n_180),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_14),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_14),
.A2(n_37),
.B1(n_39),
.B2(n_160),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_160),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_14),
.A2(n_47),
.B1(n_51),
.B2(n_160),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_16),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_16),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_16),
.A2(n_41),
.B1(n_47),
.B2(n_51),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_21),
.B(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_81),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_22),
.A2(n_74),
.B1(n_75),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_23),
.A2(n_24),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_44),
.C(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_34),
.A3(n_39),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_30),
.A2(n_36),
.B1(n_40),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_30),
.A2(n_36),
.B1(n_97),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_30),
.A2(n_36),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_30),
.A2(n_36),
.B1(n_179),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_31),
.A2(n_134),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_33),
.B(n_37),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_36),
.Y(n_161)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_39),
.B1(n_66),
.B2(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_37),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_39),
.A2(n_55),
.A3(n_66),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_59),
.B1(n_60),
.B2(n_73),
.Y(n_43)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_44),
.A2(n_73),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_52),
.B(n_57),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_52),
.B1(n_57),
.B2(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_52),
.B1(n_80),
.B2(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_45),
.A2(n_52),
.B1(n_94),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_45),
.A2(n_52),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_45),
.A2(n_52),
.B1(n_202),
.B2(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_45),
.A2(n_52),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_45),
.A2(n_52),
.B1(n_230),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_46),
.A2(n_128),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_46),
.A2(n_153),
.B1(n_201),
.B2(n_242),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_47),
.B(n_258),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_52),
.Y(n_153)
);

AO22x2_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_54),
.B(n_68),
.Y(n_207)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_55),
.B(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_65),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_71),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_78),
.B1(n_106),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_64),
.A2(n_106),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_64),
.A2(n_106),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_64),
.A2(n_106),
.B1(n_176),
.B2(n_192),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_64),
.A2(n_106),
.B1(n_191),
.B2(n_239),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_81),
.B(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_95),
.B(n_96),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_82),
.A2(n_83),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_95),
.B1(n_96),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_87),
.B1(n_124),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_85),
.A2(n_87),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_85),
.A2(n_87),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_86),
.A2(n_88),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_86),
.A2(n_88),
.B1(n_173),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_86),
.A2(n_88),
.B1(n_210),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_86),
.A2(n_88),
.B1(n_206),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_86),
.A2(n_88),
.B1(n_260),
.B2(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_298),
.B(n_303),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_162),
.B(n_297),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_144),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_117),
.B(n_144),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_136),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_118),
.B(n_138),
.C(n_143),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_132),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_120),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_132),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_149),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.C(n_158),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_151),
.B(n_154),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_158),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_185),
.B(n_296),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_183),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_164),
.B(n_183),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_182),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_165),
.B(n_182),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_167),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.C(n_178),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_168),
.B(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_172),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_175),
.B(n_178),
.Y(n_286)
);

AOI31xp33_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_280),
.A3(n_289),
.B(n_293),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_225),
.B(n_279),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_212),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_212),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_199),
.C(n_203),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_194),
.C(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_203),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_217),
.B(n_220),
.C(n_224),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_274),
.B(n_278),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_243),
.B(n_273),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_232),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_238),
.C(n_241),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_254),
.B(n_272),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_266),
.B(n_271),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_261),
.B(n_265),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_302),
.Y(n_303)
);


endmodule