module fake_netlist_6_4437_n_359 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_359);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;

output n_359;

wire n_52;
wire n_91;
wire n_326;
wire n_256;
wire n_209;
wire n_63;
wire n_223;
wire n_278;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_22;
wire n_208;
wire n_68;
wire n_316;
wire n_28;
wire n_304;
wire n_212;
wire n_50;
wire n_144;
wire n_125;
wire n_168;
wire n_297;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_350;
wire n_78;
wire n_84;
wire n_142;
wire n_143;
wire n_180;
wire n_62;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_67;
wire n_246;
wire n_38;
wire n_289;
wire n_59;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_353;
wire n_65;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_71;
wire n_74;
wire n_229;
wire n_305;
wire n_72;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_35;
wire n_183;
wire n_79;
wire n_338;
wire n_56;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_39;
wire n_344;
wire n_73;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_20;
wire n_155;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_218;
wire n_70;
wire n_234;
wire n_37;
wire n_82;
wire n_27;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_58;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_48;
wire n_25;
wire n_93;
wire n_80;
wire n_196;
wire n_352;
wire n_107;
wire n_89;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_69;
wire n_293;
wire n_31;
wire n_334;
wire n_53;
wire n_44;
wire n_232;
wire n_163;
wire n_46;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_83;
wire n_323;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_32;
wire n_66;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_23;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_33;
wire n_61;
wire n_237;
wire n_244;
wire n_76;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_40;
wire n_240;
wire n_139;
wire n_319;
wire n_41;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_30;
wire n_275;
wire n_43;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_21;
wire n_193;
wire n_269;
wire n_346;
wire n_88;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_49;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_90;
wire n_347;
wire n_24;
wire n_54;
wire n_328;
wire n_87;
wire n_195;
wire n_285;
wire n_85;
wire n_99;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_19;
wire n_47;
wire n_29;
wire n_75;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_81;
wire n_36;
wire n_26;
wire n_55;
wire n_267;
wire n_339;
wire n_315;
wire n_64;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_60;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_51;
wire n_283;

INVx1_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_19),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_6),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_36),
.Y(n_51)
);

AO21x2_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_41),
.B(n_32),
.Y(n_52)
);

BUFx8_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_22),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_26),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_33),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_38),
.B1(n_47),
.B2(n_28),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_37),
.B1(n_23),
.B2(n_30),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_21),
.B1(n_23),
.B2(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_10),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_12),
.B(n_63),
.C(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_51),
.B(n_59),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_54),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_60),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_54),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_R g92 ( 
.A(n_54),
.B(n_55),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx8_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_52),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_55),
.B(n_54),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_55),
.B1(n_65),
.B2(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_65),
.B(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_65),
.B(n_87),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_72),
.B(n_82),
.C(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_87),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_90),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_70),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_90),
.B(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_87),
.B(n_80),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_90),
.B1(n_86),
.B2(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_68),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_88),
.B(n_92),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI211xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_86),
.B(n_94),
.C(n_68),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_R g142 ( 
.A(n_97),
.B(n_94),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI21x1_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_108),
.B(n_127),
.Y(n_144)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_68),
.B(n_94),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_68),
.B1(n_85),
.B2(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_85),
.B1(n_105),
.B2(n_104),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

AO32x2_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_116),
.A3(n_126),
.B1(n_101),
.B2(n_124),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_104),
.B(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_85),
.B(n_114),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_100),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_122),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_112),
.B(n_103),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_109),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_126),
.B1(n_116),
.B2(n_122),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_116),
.B1(n_124),
.B2(n_101),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_150),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_124),
.B(n_116),
.C(n_109),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_114),
.B(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

AND2x6_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_96),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_99),
.B1(n_120),
.B2(n_114),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_120),
.B(n_85),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_120),
.B1(n_99),
.B2(n_85),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_85),
.B1(n_99),
.B2(n_136),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_85),
.B(n_157),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_137),
.B1(n_152),
.B2(n_155),
.C(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_155),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_147),
.B(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_143),
.B1(n_149),
.B2(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_143),
.B1(n_149),
.B2(n_140),
.C(n_128),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_149),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_140),
.B(n_134),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_151),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_140),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_130),
.B1(n_140),
.B2(n_134),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_151),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_164),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_151),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_164),
.Y(n_217)
);

OAI33xp33_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_172),
.A3(n_177),
.B1(n_169),
.B2(n_135),
.B3(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

AO31x2_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_205),
.A3(n_171),
.B(n_193),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_151),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_201),
.Y(n_224)
);

OAI321xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_173),
.A3(n_175),
.B1(n_184),
.B2(n_179),
.C(n_170),
.Y(n_225)
);

AOI211xp5_ASAP7_75t_SL g226 ( 
.A1(n_211),
.A2(n_174),
.B(n_186),
.C(n_187),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_187),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_187),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_182),
.B1(n_132),
.B2(n_135),
.C(n_154),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_210),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_210),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_192),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_192),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_200),
.B(n_194),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_209),
.C(n_207),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_200),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_202),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_229),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_202),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_198),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_229),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_198),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_209),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_217),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_247),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_227),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_221),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_221),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_213),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_219),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_221),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_219),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_231),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_236),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_225),
.B(n_237),
.C(n_226),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_237),
.A3(n_239),
.B1(n_242),
.B2(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_236),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_256),
.Y(n_286)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_239),
.A3(n_252),
.B1(n_248),
.B2(n_246),
.C1(n_251),
.C2(n_249),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_242),
.B1(n_209),
.B2(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_248),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_252),
.Y(n_290)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_252),
.A3(n_212),
.B1(n_251),
.B2(n_208),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_253),
.B(n_224),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_271),
.Y(n_298)
);

AOI221xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_263),
.B1(n_218),
.B2(n_256),
.C(n_268),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_260),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_268),
.Y(n_302)
);

OAI222xp33_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_260),
.B1(n_270),
.B2(n_273),
.C1(n_253),
.C2(n_264),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_253),
.B1(n_198),
.B2(n_252),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_278),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_R g312 ( 
.A(n_302),
.B(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_286),
.Y(n_313)
);

AOI221xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_281),
.B1(n_288),
.B2(n_291),
.C(n_290),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_253),
.B1(n_270),
.B2(n_198),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_287),
.B1(n_277),
.B2(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_285),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_291),
.B(n_142),
.Y(n_323)
);

NOR4xp25_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_309),
.C(n_310),
.D(n_301),
.Y(n_324)
);

AOI221xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_310),
.B1(n_300),
.B2(n_273),
.C(n_274),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_300),
.B(n_275),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

AOI211xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_274),
.B(n_264),
.C(n_251),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_203),
.C(n_208),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_198),
.B1(n_203),
.B2(n_193),
.Y(n_330)
);

NAND5xp2_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_232),
.C(n_145),
.D(n_142),
.E(n_198),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_319),
.A2(n_201),
.B(n_190),
.Y(n_332)
);

OAI211xp5_ASAP7_75t_SL g333 ( 
.A1(n_317),
.A2(n_134),
.B(n_132),
.C(n_153),
.Y(n_333)
);

OAI311xp33_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_221),
.A3(n_198),
.B1(n_134),
.C1(n_130),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_138),
.B(n_144),
.C(n_156),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_322),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_315),
.C(n_145),
.Y(n_339)
);

AND2x4_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_198),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_198),
.B1(n_130),
.B2(n_167),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_337),
.A2(n_324),
.B1(n_326),
.B2(n_328),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

NAND4xp25_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_331),
.C(n_330),
.D(n_333),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_334),
.Y(n_345)
);

NAND4xp25_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_132),
.C(n_154),
.D(n_135),
.Y(n_346)
);

OR3x1_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_340),
.C(n_341),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_167),
.B1(n_160),
.B2(n_153),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_221),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_167),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_350),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_349),
.B1(n_153),
.B2(n_134),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_356),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

AOI222xp33_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.C1(n_144),
.C2(n_138),
.Y(n_359)
);


endmodule