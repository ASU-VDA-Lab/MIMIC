module fake_jpeg_12934_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_67),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_25),
.B1(n_35),
.B2(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_52),
.B(n_65),
.Y(n_98)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_31),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_73),
.B1(n_25),
.B2(n_35),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_6),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_6),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_28),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_76),
.B(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_84),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_89),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_108),
.B1(n_64),
.B2(n_32),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_21),
.B(n_34),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_104),
.B(n_79),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_20),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_32),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_126),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_40),
.B1(n_70),
.B2(n_42),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_58),
.B1(n_68),
.B2(n_55),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_69),
.B1(n_28),
.B2(n_33),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_139),
.B(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_81),
.B(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_33),
.B1(n_36),
.B2(n_12),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_75),
.B(n_10),
.C(n_11),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_133),
.C(n_151),
.Y(n_157)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_10),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_127),
.Y(n_159)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_12),
.B(n_13),
.C(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_36),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_137),
.Y(n_163)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_82),
.A2(n_95),
.B(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_36),
.B1(n_99),
.B2(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_143),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_114),
.B1(n_80),
.B2(n_96),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_148),
.B1(n_104),
.B2(n_77),
.Y(n_153)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_85),
.A2(n_90),
.B1(n_102),
.B2(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_102),
.B1(n_100),
.B2(n_86),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_116),
.Y(n_169)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_74),
.B(n_79),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_132),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_117),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_151),
.C(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_119),
.B(n_130),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_148),
.B(n_139),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_189),
.B(n_179),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_120),
.B1(n_140),
.B2(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_196),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_177),
.B(n_154),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_192),
.C(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_149),
.C(n_135),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_191),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_131),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_146),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_145),
.Y(n_192)
);

NOR4xp25_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_158),
.C(n_161),
.D(n_153),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_128),
.B1(n_129),
.B2(n_169),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_156),
.B1(n_171),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_179),
.B1(n_172),
.B2(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_186),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_185),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_171),
.B1(n_176),
.B2(n_152),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_199),
.B(n_168),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_214),
.Y(n_224)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_164),
.B1(n_176),
.B2(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_206),
.C(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_215),
.C(n_206),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_222),
.C(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_227),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_187),
.C(n_190),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_203),
.A3(n_205),
.B1(n_202),
.B2(n_210),
.C1(n_194),
.C2(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_184),
.C(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_236),
.C(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_189),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_240),
.Y(n_247)
);

AOI21x1_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_225),
.B(n_217),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_225),
.B(n_183),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_224),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_208),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_248),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_240),
.B(n_207),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_216),
.B1(n_188),
.B2(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_239),
.A3(n_212),
.B1(n_191),
.B2(n_182),
.C1(n_180),
.C2(n_160),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_244),
.Y(n_252)
);

OAI31xp33_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_245),
.A3(n_212),
.B(n_168),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_212),
.Y(n_255)
);


endmodule