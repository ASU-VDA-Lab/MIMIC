module fake_jpeg_23344_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_31),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_50),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_23),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_36),
.B1(n_22),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_66),
.B1(n_71),
.B2(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_22),
.B1(n_35),
.B2(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_28),
.B1(n_37),
.B2(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_28),
.B1(n_37),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_27),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_37),
.B1(n_33),
.B2(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_85),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_25),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_34),
.B1(n_28),
.B2(n_31),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_32),
.B1(n_19),
.B2(n_3),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_32),
.B(n_19),
.C(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_101),
.Y(n_123)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_96),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_23),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_2),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_107),
.Y(n_134)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_53),
.B(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_53),
.B(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_32),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_50),
.B(n_20),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_18),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_57),
.B1(n_66),
.B2(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_1),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_61),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_82),
.Y(n_144)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_126),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_114),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_77),
.C(n_66),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_138),
.C(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_128),
.Y(n_166)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_70),
.B1(n_52),
.B2(n_58),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_91),
.B1(n_104),
.B2(n_94),
.Y(n_182)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_136),
.Y(n_171)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_145),
.B1(n_154),
.B2(n_117),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_66),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_99),
.Y(n_159)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_56),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_99),
.Y(n_156)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_103),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_54),
.B(n_52),
.C(n_73),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_153),
.B(n_104),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_100),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_78),
.B1(n_56),
.B2(n_6),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_113),
.B(n_88),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_175),
.B(n_123),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_164),
.B(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_113),
.B1(n_96),
.B2(n_99),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_177),
.B1(n_179),
.B2(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_162),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_184),
.B1(n_140),
.B2(n_143),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_4),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_5),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_168),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_121),
.B(n_89),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_128),
.B(n_131),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_180),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_107),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_111),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_109),
.B1(n_92),
.B2(n_93),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_106),
.B1(n_100),
.B2(n_97),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_185),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_206),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_151),
.B(n_145),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_145),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_156),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_140),
.B1(n_136),
.B2(n_131),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_139),
.B1(n_126),
.B2(n_122),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_169),
.A2(n_112),
.B1(n_148),
.B2(n_133),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_112),
.B1(n_6),
.B2(n_8),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_179),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_184),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_219),
.B(n_235),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_238),
.Y(n_243)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_241),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_215),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_231),
.B(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_158),
.Y(n_235)
);

XOR2x2_ASAP7_75t_SL g236 ( 
.A(n_190),
.B(n_169),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_239),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_159),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_190),
.C(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_174),
.B(n_155),
.C(n_164),
.D(n_167),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

NAND5xp2_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_164),
.C(n_167),
.D(n_175),
.E(n_172),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_246),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_193),
.B1(n_207),
.B2(n_194),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_251),
.B1(n_253),
.B2(n_258),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_194),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_214),
.B1(n_205),
.B2(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_193),
.B1(n_197),
.B2(n_204),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_182),
.B1(n_199),
.B2(n_208),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.C(n_256),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_213),
.C(n_209),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_225),
.A2(n_229),
.B1(n_232),
.B2(n_163),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_212),
.B(n_170),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_259),
.A2(n_230),
.B(n_223),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_216),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_228),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_262),
.A2(n_274),
.B1(n_278),
.B2(n_253),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_234),
.C(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_267),
.C(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_229),
.C(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_272),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_240),
.C(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_241),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_227),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_228),
.C(n_160),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_173),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_160),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_245),
.B1(n_250),
.B2(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

AO22x1_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_264),
.B1(n_268),
.B2(n_12),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_248),
.B(n_251),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_265),
.B(n_264),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_248),
.B1(n_187),
.B2(n_183),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_5),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_290),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_8),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_276),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_285),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.C(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_10),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_287),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_286),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_305),
.C(n_307),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_308),
.C(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_290),
.C(n_281),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_293),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_301),
.B1(n_300),
.B2(n_293),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_316),
.A3(n_11),
.B1(n_13),
.B2(n_16),
.C1(n_17),
.C2(n_301),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_312),
.B(n_311),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_317),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);


endmodule