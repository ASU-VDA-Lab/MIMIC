module fake_jpeg_2250_n_142 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_34),
.Y(n_51)
);

BUFx2_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_3),
.B1(n_6),
.B2(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_27),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_19),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_56),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_57),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_21),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_24),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_71),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_19),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_64),
.B1(n_74),
.B2(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_81),
.B1(n_67),
.B2(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_45),
.B1(n_33),
.B2(n_41),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_30),
.B(n_51),
.C(n_62),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_104),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_107),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_82),
.C(n_79),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_116),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_82),
.B(n_81),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_82),
.B1(n_84),
.B2(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_91),
.C(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_124),
.B(n_112),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_115),
.C(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_124),
.C(n_114),
.Y(n_133)
);

BUFx12f_ASAP7_75t_SL g127 ( 
.A(n_121),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_133),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_97),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_108),
.B(n_97),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_104),
.B(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_108),
.B1(n_97),
.B2(n_95),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.C(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_87),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_87),
.Y(n_142)
);


endmodule