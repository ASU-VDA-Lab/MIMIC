module fake_aes_5341_n_28 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
BUFx6f_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
NAND2xp33_ASAP7_75t_SL g11 ( .A(n_6), .B(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_15) );
OR2x6_ASAP7_75t_L g16 ( .A(n_12), .B(n_0), .Y(n_16) );
AOI22xp33_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_11), .B1(n_10), .B2(n_2), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AOI31xp33_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_15), .A3(n_16), .B(n_1), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_10), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_23), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI222xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_7), .B1(n_10), .B2(n_25), .C1(n_11), .C2(n_24), .Y(n_28) );
endmodule