module fake_jpeg_29752_n_49 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_49);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_17),
.B2(n_22),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_32),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_9),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_40),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_12),
.Y(n_43)
);

OA21x2_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_45),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_44),
.C(n_45),
.Y(n_49)
);


endmodule