module fake_netlist_1_10412_n_666 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_666);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_82), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_73), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_69), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_43), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_12), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_47), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_14), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_35), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_22), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_25), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_27), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_54), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_20), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_11), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_5), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_87), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_80), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_63), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_2), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_55), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_64), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_37), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_34), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_41), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_88), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_124), .B(n_0), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_124), .B(n_1), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_110), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_109), .A2(n_39), .B(n_85), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_94), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_93), .B(n_1), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_105), .B(n_2), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_110), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_102), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_105), .B(n_3), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_94), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_102), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_108), .B(n_3), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_100), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_108), .B(n_4), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_99), .B(n_6), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_137), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_150), .B(n_112), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_141), .B(n_109), .Y(n_161) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_130), .B(n_121), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_141), .A2(n_106), .B1(n_98), .B2(n_126), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
AND2x4_ASAP7_75t_SL g165 ( .A(n_146), .B(n_101), .Y(n_165) );
BUFx10_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_144), .B(n_122), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_129), .B(n_112), .Y(n_168) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_153), .A2(n_138), .B(n_117), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_144), .B(n_95), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_145), .B(n_122), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_143), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_145), .B(n_90), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_129), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_146), .B(n_93), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_146), .B(n_96), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_151), .B(n_114), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_170), .B(n_149), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
NOR3xp33_ASAP7_75t_SL g194 ( .A(n_158), .B(n_113), .C(n_138), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_182), .A2(n_139), .B1(n_142), .B2(n_149), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
AND3x1_ASAP7_75t_L g198 ( .A(n_160), .B(n_147), .C(n_139), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_182), .B(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_170), .B(n_142), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_157), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_168), .B(n_165), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_166), .B(n_89), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_170), .A2(n_126), .B1(n_96), .B2(n_98), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_168), .B(n_183), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_170), .A2(n_147), .B1(n_116), .B2(n_106), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g209 ( .A(n_170), .B(n_136), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_162), .A2(n_136), .B(n_117), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_166), .B(n_91), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_178), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_165), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_166), .B(n_92), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_183), .A2(n_116), .B1(n_104), .B2(n_114), .Y(n_215) );
BUFx12f_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_183), .A2(n_118), .B1(n_115), .B2(n_119), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_168), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_178), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_166), .B(n_97), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_187), .B(n_136), .Y(n_223) );
BUFx6f_ASAP7_75t_SL g224 ( .A(n_188), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_187), .B(n_119), .Y(n_225) );
BUFx12f_ASAP7_75t_L g226 ( .A(n_158), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_178), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_175), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_186), .B(n_107), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_175), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_187), .A2(n_118), .B1(n_128), .B2(n_123), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_118), .B1(n_127), .B2(n_123), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_165), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_230), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_191), .B(n_165), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_220), .A2(n_188), .B1(n_175), .B2(n_180), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_191), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_199), .B(n_175), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_195), .A2(n_190), .B1(n_189), .B2(n_163), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_230), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_179), .B1(n_162), .B2(n_169), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_230), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_191), .B(n_175), .Y(n_245) );
AOI21xp33_ASAP7_75t_L g246 ( .A1(n_203), .A2(n_179), .B(n_169), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_207), .B(n_175), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_223), .A2(n_176), .B(n_189), .C(n_190), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_203), .B(n_169), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_216), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_230), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_223), .A2(n_174), .B(n_159), .C(n_171), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_232), .A2(n_164), .B(n_171), .C(n_174), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_191), .B(n_111), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_195), .A2(n_163), .B1(n_176), .B2(n_164), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_200), .B(n_188), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_193), .B(n_169), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_228), .B(n_125), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_232), .A2(n_188), .B(n_161), .C(n_167), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_213), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_197), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_196), .B(n_188), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_224), .Y(n_266) );
CKINVDCx11_ASAP7_75t_R g267 ( .A(n_226), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_225), .B(n_188), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_233), .A2(n_161), .B(n_167), .C(n_127), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_208), .A2(n_118), .B1(n_128), .B2(n_120), .C(n_152), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_225), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_198), .A2(n_169), .B1(n_118), .B2(n_128), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_226), .B(n_118), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_184), .B(n_177), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_208), .A2(n_120), .B1(n_121), .B2(n_184), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_197), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_233), .A2(n_173), .B(n_184), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_225), .A2(n_154), .B(n_152), .C(n_135), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
OAI222xp33_ASAP7_75t_L g281 ( .A1(n_273), .A2(n_235), .B1(n_217), .B2(n_234), .C1(n_209), .C2(n_215), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_239), .B(n_225), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_275), .A2(n_209), .B(n_234), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_275), .A2(n_209), .B(n_231), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_280), .B(n_197), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_250), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_237), .B(n_235), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_266), .B(n_205), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_249), .A2(n_192), .B(n_202), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_277), .Y(n_291) );
OR2x6_ASAP7_75t_L g292 ( .A(n_266), .B(n_211), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_248), .A2(n_206), .B(n_194), .C(n_222), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_244), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_237), .B(n_214), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_248), .A2(n_217), .B(n_192), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_280), .B(n_202), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
AOI21x1_ASAP7_75t_L g299 ( .A1(n_278), .A2(n_135), .B(n_152), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_262), .B(n_215), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_239), .B(n_229), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_249), .A2(n_259), .B(n_279), .C(n_246), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_242), .Y(n_304) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_252), .A2(n_154), .B(n_135), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_253), .B(n_212), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_279), .A2(n_212), .B(n_219), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_259), .B(n_219), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_201), .Y(n_309) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_261), .A2(n_154), .B(n_132), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_268), .B(n_201), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_278), .A2(n_227), .B(n_221), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_276), .A2(n_227), .B(n_221), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_241), .A2(n_218), .B(n_204), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g315 ( .A(n_280), .B(n_204), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_251), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_303), .A2(n_254), .B(n_247), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_308), .A2(n_269), .B(n_257), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_301), .A2(n_238), .B1(n_243), .B2(n_245), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_281), .A2(n_264), .B1(n_272), .B2(n_238), .C(n_271), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g322 ( .A1(n_293), .A2(n_267), .B(n_255), .C(n_265), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_282), .A2(n_240), .B1(n_258), .B2(n_274), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_282), .B(n_245), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_281), .A2(n_253), .B1(n_270), .B2(n_260), .C(n_256), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_308), .A2(n_274), .B1(n_218), .B2(n_121), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_295), .A2(n_274), .B1(n_121), .B2(n_9), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_7), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_290), .A2(n_131), .B1(n_132), .B2(n_156), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_295), .A2(n_173), .B1(n_184), .B2(n_177), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_295), .A2(n_173), .B1(n_184), .B2(n_177), .Y(n_333) );
BUFx12f_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_314), .A2(n_132), .B(n_131), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_290), .A2(n_172), .B(n_185), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_316), .Y(n_337) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_288), .B(n_287), .C(n_302), .Y(n_338) );
NOR2x1p5_ASAP7_75t_L g339 ( .A(n_300), .B(n_8), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_309), .B(n_10), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_299), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_300), .B(n_177), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_302), .A2(n_295), .B1(n_292), .B2(n_289), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_295), .A2(n_131), .B(n_11), .Y(n_344) );
OAI222xp33_ASAP7_75t_L g345 ( .A1(n_289), .A2(n_10), .B1(n_13), .B2(n_15), .C1(n_16), .C2(n_17), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_322), .B(n_306), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_329), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_334), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_319), .B(n_300), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_332), .B(n_310), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_332), .B(n_316), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_337), .B(n_310), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_337), .B(n_310), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_310), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_317), .B(n_314), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_335), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_342), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_328), .B(n_310), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_330), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_305), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_340), .B(n_305), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_305), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_345), .A2(n_311), .B1(n_306), .B2(n_298), .C(n_304), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_318), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_330), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_331), .B(n_300), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_347), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_371), .A2(n_323), .B1(n_321), .B2(n_325), .C(n_338), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_349), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_371), .A2(n_327), .B1(n_324), .B2(n_344), .C(n_323), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_352), .B(n_305), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_357), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_352), .B(n_305), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_352), .B(n_296), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
NOR2x1p5_ASAP7_75t_L g388 ( .A(n_368), .B(n_334), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_368), .A2(n_326), .B1(n_333), .B2(n_289), .C(n_292), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_357), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_354), .B(n_314), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_362), .B(n_289), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_355), .B(n_283), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_359), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_363), .B(n_283), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_363), .B(n_283), .Y(n_401) );
INVx5_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_363), .B(n_284), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_370), .B(n_296), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_369), .B(n_326), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_370), .B(n_296), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_372), .A2(n_284), .B(n_336), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_401), .B(n_365), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_401), .B(n_365), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_401), .B(n_365), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_400), .B(n_366), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_400), .B(n_366), .Y(n_416) );
NAND2x1_ASAP7_75t_L g417 ( .A(n_399), .B(n_369), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_398), .B(n_366), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_398), .B(n_367), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_387), .B(n_372), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_387), .B(n_351), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_392), .B(n_356), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_398), .B(n_367), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_367), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_393), .B(n_351), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_393), .B(n_351), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_402), .B(n_362), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_394), .B(n_351), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_394), .B(n_356), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_403), .B(n_385), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_399), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_403), .B(n_358), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_376), .A2(n_346), .B(n_353), .C(n_358), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_404), .B(n_353), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_403), .B(n_360), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_385), .B(n_364), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_389), .A2(n_348), .B(n_374), .C(n_297), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_385), .B(n_374), .Y(n_446) );
OAI21x1_ASAP7_75t_L g447 ( .A1(n_407), .A2(n_361), .B(n_373), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_380), .B(n_364), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_380), .B(n_364), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
AOI211x1_ASAP7_75t_SL g452 ( .A1(n_386), .A2(n_373), .B(n_297), .C(n_156), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_373), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_378), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_405), .B(n_361), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_378), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_378), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_381), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_388), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_432), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_446), .A2(n_407), .B(n_376), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_439), .A2(n_389), .B1(n_374), .B2(n_379), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_429), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_437), .Y(n_469) );
NOR2x1p5_ASAP7_75t_L g470 ( .A(n_461), .B(n_395), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_436), .B(n_408), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_436), .B(n_408), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_423), .B(n_386), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_432), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
NAND2xp33_ASAP7_75t_L g478 ( .A(n_461), .B(n_388), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_425), .B(n_391), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_411), .B(n_391), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_458), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_411), .B(n_381), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
NOR2xp33_ASAP7_75t_SL g486 ( .A(n_445), .B(n_402), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_432), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_425), .B(n_379), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_415), .B(n_381), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_417), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_430), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_433), .B(n_395), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_412), .B(n_382), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_412), .B(n_382), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_420), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_414), .B(n_382), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_414), .B(n_384), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_423), .B(n_384), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_435), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_434), .B(n_384), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_447), .A2(n_396), .B(n_402), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_431), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_418), .B(n_390), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_434), .B(n_390), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
NAND2x1_ASAP7_75t_L g506 ( .A(n_453), .B(n_390), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_418), .B(n_397), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_419), .B(n_397), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_419), .B(n_397), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_424), .B(n_402), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_433), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_454), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_422), .B(n_396), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_424), .B(n_402), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_427), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_433), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_415), .B(n_410), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_428), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_416), .B(n_438), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_514), .Y(n_523) );
AOI211x1_ASAP7_75t_L g524 ( .A1(n_465), .A2(n_441), .B(n_416), .C(n_438), .Y(n_524) );
INVxp33_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_522), .B(n_441), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_522), .B(n_516), .Y(n_527) );
OAI322xp33_ASAP7_75t_L g528 ( .A1(n_488), .A2(n_455), .A3(n_457), .B1(n_449), .B2(n_443), .C1(n_451), .C2(n_460), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_489), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_482), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_506), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_466), .A2(n_374), .B1(n_444), .B2(n_450), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_479), .A2(n_457), .B(n_455), .C(n_456), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_467), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g535 ( .A1(n_463), .A2(n_452), .A3(n_444), .B1(n_448), .B2(n_450), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_491), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_502), .Y(n_537) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_467), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_487), .A2(n_402), .B1(n_396), .B2(n_448), .Y(n_540) );
NAND2x1_ASAP7_75t_L g541 ( .A(n_490), .B(n_361), .Y(n_541) );
OA21x2_ASAP7_75t_SL g542 ( .A1(n_475), .A2(n_402), .B(n_15), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_478), .A2(n_292), .B1(n_410), .B2(n_447), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
AOI21xp33_ASAP7_75t_SL g546 ( .A1(n_490), .A2(n_13), .B(n_16), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_477), .B(n_18), .Y(n_547) );
NAND2xp33_ASAP7_75t_SL g548 ( .A(n_487), .B(n_410), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_518), .A2(n_156), .B1(n_306), .B2(n_311), .C(n_410), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_521), .B(n_18), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_462), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_499), .B(n_19), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_464), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_478), .A2(n_292), .B1(n_306), .B2(n_315), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_481), .B(n_156), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_486), .A2(n_292), .B(n_312), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_484), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_520), .A2(n_156), .B1(n_284), .B2(n_21), .C1(n_22), .C2(n_20), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_481), .B(n_156), .Y(n_559) );
OAI322xp33_ASAP7_75t_L g560 ( .A1(n_471), .A2(n_19), .A3(n_21), .B1(n_342), .B2(n_291), .C1(n_285), .C2(n_304), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_468), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_469), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_520), .B(n_312), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_513), .B(n_312), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_512), .A2(n_342), .B1(n_286), .B2(n_315), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_513), .A2(n_291), .B(n_285), .C(n_304), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_493), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_494), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_483), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_494), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_519), .B(n_313), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g575 ( .A1(n_519), .A2(n_291), .B1(n_285), .B2(n_298), .C1(n_185), .C2(n_172), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_524), .B(n_480), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_557), .Y(n_577) );
OAI321xp33_ASAP7_75t_L g578 ( .A1(n_542), .A2(n_517), .A3(n_515), .B1(n_472), .B2(n_476), .C(n_473), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_526), .B(n_496), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_555), .B(n_509), .Y(n_580) );
XNOR2xp5_ASAP7_75t_L g581 ( .A(n_525), .B(n_509), .Y(n_581) );
O2A1O1Ixp5_ASAP7_75t_SL g582 ( .A1(n_545), .A2(n_497), .B(n_503), .C(n_507), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_523), .B(n_510), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_534), .A2(n_472), .B(n_476), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g585 ( .A1(n_534), .A2(n_474), .B1(n_501), .B2(n_500), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_530), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_536), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_537), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_559), .B(n_510), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_539), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_527), .B(n_474), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_532), .B(n_498), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_551), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_553), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_528), .A2(n_515), .B1(n_511), .B2(n_508), .C(n_485), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_532), .B(n_504), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_529), .Y(n_598) );
OA22x2_ASAP7_75t_L g599 ( .A1(n_538), .A2(n_492), .B1(n_508), .B2(n_485), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_538), .A2(n_504), .B1(n_500), .B2(n_498), .Y(n_600) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_571), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_561), .Y(n_602) );
AOI32xp33_ASAP7_75t_L g603 ( .A1(n_552), .A2(n_492), .A3(n_511), .B1(n_313), .B2(n_298), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_566), .B(n_492), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_567), .B(n_313), .Y(n_606) );
OA22x2_ASAP7_75t_L g607 ( .A1(n_540), .A2(n_307), .B1(n_24), .B2(n_26), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_552), .A2(n_286), .B1(n_185), .B2(n_172), .C(n_177), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_569), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_548), .B(n_185), .C(n_172), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_543), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_583), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_578), .A2(n_547), .B1(n_550), .B2(n_535), .C1(n_563), .C2(n_571), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_576), .A2(n_547), .B(n_531), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g615 ( .A1(n_603), .A2(n_546), .B(n_558), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_599), .B(n_574), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_599), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_582), .B(n_549), .C(n_533), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_576), .A2(n_570), .B1(n_572), .B2(n_565), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_578), .A2(n_560), .B(n_565), .C(n_568), .Y(n_620) );
XOR2x2_ASAP7_75t_L g621 ( .A(n_581), .B(n_554), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_611), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_598), .B(n_564), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_607), .A2(n_556), .B(n_568), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_585), .A2(n_573), .B1(n_544), .B2(n_575), .C(n_541), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_607), .A2(n_307), .B(n_173), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_580), .B(n_23), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_593), .A2(n_307), .B1(n_173), .B2(n_181), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_597), .A2(n_181), .B1(n_29), .B2(n_30), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_596), .A2(n_181), .B1(n_31), .B2(n_32), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_608), .A2(n_181), .B1(n_33), .B2(n_38), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_610), .A2(n_28), .B(n_42), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_584), .B1(n_601), .B2(n_586), .C(n_591), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g635 ( .A1(n_614), .A2(n_592), .A3(n_600), .B1(n_579), .B2(n_583), .C1(n_605), .C2(n_590), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_615), .A2(n_587), .B1(n_588), .B2(n_589), .C(n_609), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_612), .B(n_604), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_625), .A2(n_602), .B1(n_595), .B2(n_594), .Y(n_638) );
NAND4xp75_ASAP7_75t_L g639 ( .A(n_630), .B(n_606), .C(n_45), .D(n_46), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_613), .B(n_44), .C(n_48), .D(n_49), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_623), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_619), .A2(n_50), .B(n_51), .C(n_52), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_617), .A2(n_181), .B1(n_56), .B2(n_57), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_613), .B(n_181), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_632), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_620), .A2(n_181), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_638), .A2(n_624), .B1(n_621), .B2(n_618), .C(n_616), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_644), .B(n_618), .C(n_633), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_646), .B(n_629), .C(n_631), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_640), .A2(n_627), .B1(n_622), .B2(n_628), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_634), .B(n_626), .C(n_65), .Y(n_651) );
AND3x4_ASAP7_75t_L g652 ( .A(n_635), .B(n_53), .C(n_67), .Y(n_652) );
CKINVDCx16_ASAP7_75t_R g653 ( .A(n_641), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_652), .B(n_639), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_648), .B(n_636), .C(n_642), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_647), .B(n_637), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_655), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_657), .B(n_651), .C(n_649), .D(n_650), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_656), .A2(n_645), .B(n_643), .Y(n_660) );
OAI22x1_ASAP7_75t_L g661 ( .A1(n_658), .A2(n_654), .B1(n_71), .B2(n_72), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_659), .A2(n_181), .B1(n_75), .B2(n_76), .C(n_77), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g663 ( .A(n_661), .B(n_660), .Y(n_663) );
OA22x2_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_662), .B1(n_78), .B2(n_79), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_181), .B1(n_81), .B2(n_83), .Y(n_665) );
AO21x2_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_68), .B(n_86), .Y(n_666) );
endmodule