module fake_jpeg_31652_n_109 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_53),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_45),
.B1(n_36),
.B2(n_43),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_57),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_41),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_44),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_72),
.C(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_74),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_37),
.B(n_31),
.C(n_13),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_1),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_2),
.B(n_3),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_10),
.B1(n_17),
.B2(n_21),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_5),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_30),
.B1(n_11),
.B2(n_16),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_6),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_93),
.B(n_77),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_94),
.B1(n_79),
.B2(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_100),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_87),
.C(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_96),
.B(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_96),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_79),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_94),
.C(n_25),
.Y(n_109)
);


endmodule