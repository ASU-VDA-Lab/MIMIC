module real_aes_9139_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g190 ( .A1(n_0), .A2(n_191), .B(n_192), .C(n_196), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_1), .B(n_186), .Y(n_197) );
INVx1_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_3), .B(n_151), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_4), .A2(n_132), .B(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_5), .A2(n_137), .B(n_142), .C(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_6), .A2(n_132), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_7), .B(n_186), .Y(n_471) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_165), .B(n_215), .Y(n_214) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_10), .A2(n_137), .B(n_142), .C(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g526 ( .A(n_11), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_12), .B(n_41), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_13), .B(n_195), .Y(n_503) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_15), .B(n_151), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_16), .A2(n_152), .B(n_511), .C(n_513), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_17), .B(n_186), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_18), .B(n_179), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_19), .A2(n_142), .B(n_173), .C(n_178), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_20), .A2(n_194), .B(n_209), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_21), .B(n_195), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_22), .A2(n_78), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_22), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_23), .B(n_195), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_24), .Y(n_452) );
INVx1_ASAP7_75t_L g477 ( .A(n_25), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_26), .A2(n_142), .B(n_178), .C(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_27), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_28), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_29), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_29), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_30), .Y(n_732) );
INVx1_ASAP7_75t_L g553 ( .A(n_31), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_32), .A2(n_132), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_34), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_35), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_36), .A2(n_194), .B(n_468), .C(n_470), .Y(n_467) );
INVxp67_ASAP7_75t_L g554 ( .A(n_37), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_38), .B(n_220), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_39), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_40), .A2(n_142), .B(n_178), .C(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_42), .A2(n_196), .B(n_524), .C(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_43), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_44), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_45), .B(n_151), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_46), .B(n_132), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_47), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_48), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_48), .A2(n_97), .B1(n_480), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_49), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_50), .A2(n_140), .B(n_155), .C(n_229), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_51), .A2(n_89), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_51), .Y(n_741) );
INVx1_ASAP7_75t_L g193 ( .A(n_52), .Y(n_193) );
INVx1_ASAP7_75t_L g230 ( .A(n_53), .Y(n_230) );
INVx1_ASAP7_75t_L g489 ( .A(n_54), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_55), .B(n_132), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_56), .A2(n_105), .B1(n_117), .B2(n_754), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_57), .Y(n_182) );
CKINVDCx14_ASAP7_75t_R g522 ( .A(n_58), .Y(n_522) );
INVx1_ASAP7_75t_L g138 ( .A(n_59), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_60), .B(n_132), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_61), .B(n_186), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_62), .A2(n_177), .B(n_240), .C(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g160 ( .A(n_63), .Y(n_160) );
INVx1_ASAP7_75t_SL g469 ( .A(n_64), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_65), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_66), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_67), .B(n_186), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_68), .B(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g455 ( .A(n_69), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_70), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_71), .B(n_148), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_72), .A2(n_142), .B(n_155), .C(n_266), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_73), .Y(n_238) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_75), .A2(n_132), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_76), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_77), .A2(n_132), .B(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_78), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_79), .A2(n_171), .B(n_549), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_80), .Y(n_474) );
INVx1_ASAP7_75t_L g509 ( .A(n_81), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_82), .B(n_147), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_83), .A2(n_720), .B1(n_726), .B2(n_727), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_83), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_84), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_85), .A2(n_132), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g512 ( .A(n_86), .Y(n_512) );
INVx2_ASAP7_75t_L g158 ( .A(n_87), .Y(n_158) );
INVx1_ASAP7_75t_L g502 ( .A(n_88), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_89), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_90), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_91), .B(n_195), .Y(n_207) );
OR2x2_ASAP7_75t_L g112 ( .A(n_92), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g122 ( .A(n_92), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_93), .A2(n_142), .B(n_155), .C(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_94), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
INVxp67_ASAP7_75t_L g243 ( .A(n_96), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_97), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_98), .B(n_165), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_99), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g202 ( .A(n_100), .Y(n_202) );
INVx1_ASAP7_75t_L g267 ( .A(n_101), .Y(n_267) );
INVx2_ASAP7_75t_L g492 ( .A(n_102), .Y(n_492) );
AND2x2_ASAP7_75t_L g232 ( .A(n_103), .B(n_157), .Y(n_232) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g754 ( .A(n_107), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_112), .Y(n_749) );
INVx2_ASAP7_75t_L g753 ( .A(n_112), .Y(n_753) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_113), .B(n_122), .Y(n_731) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_114), .A2(n_119), .B1(n_728), .B2(n_732), .Y(n_118) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AO221x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_733), .B1(n_737), .B2(n_746), .C(n_750), .Y(n_117) );
XOR2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_719), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_123), .B1(n_442), .B2(n_443), .Y(n_120) );
INVx1_ASAP7_75t_L g442 ( .A(n_121), .Y(n_442) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XOR2xp5_ASAP7_75t_L g738 ( .A(n_124), .B(n_739), .Y(n_738) );
OR3x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_356), .C(n_399), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_283), .C(n_313), .D(n_330), .E(n_345), .Y(n_125) );
AOI221xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_198), .B1(n_245), .B2(n_251), .C(n_255), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_167), .Y(n_127) );
OR2x2_ASAP7_75t_L g260 ( .A(n_128), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_128), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_128), .B(n_253), .Y(n_335) );
OR2x2_ASAP7_75t_L g347 ( .A(n_128), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_128), .B(n_306), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_128), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_128), .B(n_284), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_128), .B(n_292), .Y(n_398) );
AND2x2_ASAP7_75t_L g430 ( .A(n_128), .B(n_184), .Y(n_430) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_128), .Y(n_438) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_129), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g257 ( .A(n_129), .B(n_233), .Y(n_257) );
BUFx2_ASAP7_75t_L g280 ( .A(n_129), .Y(n_280) );
AND2x2_ASAP7_75t_L g309 ( .A(n_129), .B(n_168), .Y(n_309) );
AND2x2_ASAP7_75t_L g364 ( .A(n_129), .B(n_261), .Y(n_364) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_139), .B(n_157), .Y(n_130) );
BUFx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_133), .B(n_137), .Y(n_203) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g210 ( .A(n_135), .Y(n_210) );
INVx1_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g220 ( .A(n_136), .Y(n_220) );
INVx4_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
BUFx3_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_141), .A2(n_156), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_141), .A2(n_156), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_141), .A2(n_156), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_141), .A2(n_156), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_141), .A2(n_156), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_141), .A2(n_156), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_141), .A2(n_156), .B(n_550), .C(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_143), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_147), .A2(n_153), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_147), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g501 ( .A1(n_147), .A2(n_457), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g241 ( .A(n_149), .Y(n_241) );
INVx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_151), .B(n_243), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_151), .A2(n_176), .B(n_477), .C(n_478), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_151), .A2(n_241), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_152), .B(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx1_ASAP7_75t_L g513 ( .A(n_154), .Y(n_513) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_157), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_157), .A2(n_203), .B(n_474), .C(n_475), .Y(n_473) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_157), .A2(n_520), .B(n_527), .Y(n_519) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g166 ( .A(n_158), .B(n_159), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx3_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_211), .Y(n_200) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_164), .A2(n_264), .B(n_272), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_164), .B(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_164), .A2(n_451), .B(n_458), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_164), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_164), .B(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_165), .A2(n_216), .B(n_217), .Y(n_215) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_167), .B(n_318), .Y(n_327) );
OAI32xp33_ASAP7_75t_L g341 ( .A1(n_167), .A2(n_277), .A3(n_342), .B1(n_343), .B2(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_167), .B(n_343), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_167), .B(n_260), .Y(n_384) );
INVx1_ASAP7_75t_SL g413 ( .A(n_167), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_167), .B(n_200), .C(n_364), .D(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
INVx5_ASAP7_75t_L g254 ( .A(n_168), .Y(n_254) );
AND2x2_ASAP7_75t_L g284 ( .A(n_168), .B(n_185), .Y(n_284) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_168), .Y(n_363) );
AND2x2_ASAP7_75t_L g433 ( .A(n_168), .B(n_380), .Y(n_433) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_181), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_172), .B(n_179), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_177), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_180), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_183), .A2(n_498), .B(n_504), .Y(n_497) );
AND2x4_ASAP7_75t_L g306 ( .A(n_184), .B(n_254), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_184), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g340 ( .A(n_184), .B(n_261), .Y(n_340) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g253 ( .A(n_185), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g292 ( .A(n_185), .B(n_263), .Y(n_292) );
AND2x2_ASAP7_75t_L g301 ( .A(n_185), .B(n_262), .Y(n_301) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_194), .B(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g524 ( .A(n_195), .Y(n_524) );
INVx2_ASAP7_75t_L g457 ( .A(n_196), .Y(n_457) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_198), .A2(n_370), .B1(n_372), .B2(n_374), .C1(n_377), .C2(n_378), .Y(n_369) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_222), .Y(n_198) );
AND2x2_ASAP7_75t_L g302 ( .A(n_199), .B(n_303), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_199), .B(n_280), .C(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
INVx5_ASAP7_75t_SL g250 ( .A(n_200), .Y(n_250) );
OAI322xp33_ASAP7_75t_L g255 ( .A1(n_200), .A2(n_256), .A3(n_258), .B1(n_259), .B2(n_274), .C1(n_277), .C2(n_279), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_200), .B(n_248), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_200), .B(n_234), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_203), .A2(n_452), .B(n_453), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_203), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_221), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g547 ( .A(n_213), .Y(n_547) );
INVx2_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_214), .B(n_224), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_222), .B(n_287), .Y(n_342) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g321 ( .A(n_223), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
OR2x2_ASAP7_75t_L g249 ( .A(n_224), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_224), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g289 ( .A(n_224), .B(n_234), .Y(n_289) );
AND2x2_ASAP7_75t_L g312 ( .A(n_224), .B(n_248), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_224), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g328 ( .A(n_224), .B(n_287), .Y(n_328) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_224), .B(n_296), .Y(n_386) );
INVx5_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g276 ( .A(n_225), .B(n_250), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_225), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g303 ( .A(n_225), .B(n_234), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_225), .B(n_350), .Y(n_391) );
OR2x2_ASAP7_75t_L g407 ( .A(n_225), .B(n_351), .Y(n_407) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_225), .B(n_368), .Y(n_414) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_225), .Y(n_421) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
AND2x2_ASAP7_75t_L g275 ( .A(n_233), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g325 ( .A(n_233), .B(n_248), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_233), .B(n_250), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_233), .B(n_287), .Y(n_409) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_234), .B(n_250), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_234), .B(n_248), .Y(n_297) );
OR2x2_ASAP7_75t_L g351 ( .A(n_234), .B(n_248), .Y(n_351) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_247), .Y(n_368) );
INVxp67_ASAP7_75t_L g390 ( .A(n_234), .Y(n_390) );
AND2x2_ASAP7_75t_L g417 ( .A(n_234), .B(n_287), .Y(n_417) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_234), .Y(n_424) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_235), .A2(n_464), .B(n_471), .Y(n_463) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_235), .A2(n_487), .B(n_493), .Y(n_486) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_235), .A2(n_507), .B(n_514), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_240), .A2(n_267), .B(n_268), .C(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_241), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_241), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_247), .B(n_298), .Y(n_371) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g287 ( .A(n_248), .B(n_250), .Y(n_287) );
OR2x2_ASAP7_75t_L g354 ( .A(n_248), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g298 ( .A(n_249), .Y(n_298) );
OR2x2_ASAP7_75t_L g359 ( .A(n_249), .B(n_351), .Y(n_359) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g258 ( .A(n_253), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_253), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g259 ( .A(n_254), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_254), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_254), .B(n_261), .Y(n_294) );
INVx2_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
AND2x2_ASAP7_75t_L g352 ( .A(n_254), .B(n_292), .Y(n_352) );
AND2x2_ASAP7_75t_L g377 ( .A(n_254), .B(n_301), .Y(n_377) );
INVx1_ASAP7_75t_L g329 ( .A(n_259), .Y(n_329) );
INVx2_ASAP7_75t_SL g316 ( .A(n_260), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g380 ( .A(n_263), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_271), .Y(n_264) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g470 ( .A(n_270), .Y(n_470) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g349 ( .A(n_276), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_276), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_276), .A2(n_358), .B1(n_360), .B2(n_365), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_276), .B(n_368), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_277), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g311 ( .A(n_278), .Y(n_311) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g293 ( .A(n_280), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_280), .B(n_284), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_280), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g343 ( .A(n_282), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_290), .C(n_304), .Y(n_283) );
INVx1_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_284), .A2(n_416), .B1(n_418), .B2(n_419), .C(n_422), .Y(n_415) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g434 ( .A(n_287), .Y(n_434) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_322), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .B(n_295), .C(n_299), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_297), .A2(n_298), .A3(n_361), .B1(n_398), .B2(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AND2x2_ASAP7_75t_L g440 ( .A(n_300), .B(n_339), .Y(n_440) );
AND2x2_ASAP7_75t_L g387 ( .A(n_301), .B(n_339), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_301), .B(n_309), .Y(n_405) );
AOI31xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_307), .A3(n_308), .B(n_310), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_306), .B(n_318), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_306), .B(n_316), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_306), .A2(n_336), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_332), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B1(n_323), .B2(n_326), .C1(n_328), .C2(n_329), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g396 ( .A(n_315), .Y(n_396) );
INVx1_ASAP7_75t_L g418 ( .A(n_318), .Y(n_418) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_321), .A2(n_432), .B1(n_434), .B2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g337 ( .A(n_322), .Y(n_337) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_336), .B2(n_338), .C(n_341), .Y(n_330) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g375 ( .A(n_333), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g427 ( .A(n_333), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g402 ( .A(n_338), .Y(n_402) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
INVx1_ASAP7_75t_L g348 ( .A(n_340), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_343), .B(n_430), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_352), .B2(n_353), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g439 ( .A(n_352), .Y(n_439) );
INVxp33_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_354), .B(n_398), .Y(n_397) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_389), .A3(n_390), .B1(n_391), .B2(n_392), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_369), .C(n_381), .D(n_393), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
NAND2xp33_ASAP7_75t_SL g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_364), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_394), .B1(n_411), .B2(n_414), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g429 ( .A(n_380), .B(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_385), .B2(n_387), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_390), .B(n_421), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_410), .C(n_425), .D(n_436), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B(n_406), .C(n_408), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g441 ( .A(n_428), .Y(n_441) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B(n_441), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_674), .Y(n_443) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_611), .C(n_645), .D(n_661), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_446), .B(n_540), .C(n_575), .D(n_591), .Y(n_445) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_481), .B1(n_515), .B2(n_528), .C1(n_533), .C2(n_539), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g707 ( .A1(n_448), .A2(n_708), .A3(n_709), .B(n_711), .Y(n_707) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_460), .Y(n_448) );
AND2x2_ASAP7_75t_L g682 ( .A(n_449), .B(n_462), .Y(n_682) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g532 ( .A(n_450), .Y(n_532) );
AND2x2_ASAP7_75t_L g539 ( .A(n_450), .B(n_472), .Y(n_539) );
AND2x2_ASAP7_75t_L g596 ( .A(n_450), .B(n_463), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_460), .B(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_461), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_461), .B(n_543), .Y(n_586) );
AND2x2_ASAP7_75t_L g679 ( .A(n_461), .B(n_619), .Y(n_679) );
OAI321xp33_ASAP7_75t_L g713 ( .A1(n_461), .A2(n_532), .A3(n_686), .B1(n_714), .B2(n_716), .C(n_717), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_461), .B(n_518), .C(n_626), .D(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
AND2x2_ASAP7_75t_L g581 ( .A(n_462), .B(n_530), .Y(n_581) );
AND2x2_ASAP7_75t_L g600 ( .A(n_462), .B(n_532), .Y(n_600) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g556 ( .A(n_463), .B(n_472), .Y(n_556) );
AND2x2_ASAP7_75t_L g642 ( .A(n_463), .B(n_530), .Y(n_642) );
INVx3_ASAP7_75t_SL g530 ( .A(n_472), .Y(n_530) );
AND2x2_ASAP7_75t_L g574 ( .A(n_472), .B(n_561), .Y(n_574) );
OR2x2_ASAP7_75t_L g607 ( .A(n_472), .B(n_532), .Y(n_607) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_472), .Y(n_614) );
AND2x2_ASAP7_75t_L g643 ( .A(n_472), .B(n_531), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_472), .B(n_616), .Y(n_658) );
AND2x2_ASAP7_75t_L g690 ( .A(n_472), .B(n_682), .Y(n_690) );
AND2x2_ASAP7_75t_L g699 ( .A(n_472), .B(n_544), .Y(n_699) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_479), .Y(n_472) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
INVx1_ASAP7_75t_SL g667 ( .A(n_483), .Y(n_667) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g535 ( .A(n_484), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g517 ( .A(n_485), .B(n_496), .Y(n_517) );
AND2x2_ASAP7_75t_L g603 ( .A(n_485), .B(n_519), .Y(n_603) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g573 ( .A(n_486), .B(n_506), .Y(n_573) );
OR2x2_ASAP7_75t_L g584 ( .A(n_486), .B(n_519), .Y(n_584) );
AND2x2_ASAP7_75t_L g610 ( .A(n_486), .B(n_519), .Y(n_610) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_486), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_494), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_494), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g583 ( .A(n_495), .B(n_584), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g669 ( .A1(n_495), .A2(n_573), .A3(n_579), .B1(n_610), .B2(n_660), .C1(n_670), .C2(n_672), .Y(n_669) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_496), .B(n_518), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_496), .B(n_519), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_496), .B(n_536), .Y(n_590) );
AND2x2_ASAP7_75t_L g644 ( .A(n_496), .B(n_610), .Y(n_644) );
INVx1_ASAP7_75t_L g648 ( .A(n_496), .Y(n_648) );
AND2x2_ASAP7_75t_L g660 ( .A(n_496), .B(n_506), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_496), .B(n_535), .Y(n_692) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_506), .Y(n_557) );
BUFx3_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
AND3x2_ASAP7_75t_L g653 ( .A(n_497), .B(n_633), .C(n_654), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_506), .B(n_517), .C(n_518), .Y(n_516) );
INVx1_ASAP7_75t_SL g536 ( .A(n_506), .Y(n_536) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_506), .Y(n_638) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g632 ( .A(n_517), .B(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g639 ( .A(n_517), .Y(n_639) );
AND2x2_ASAP7_75t_L g677 ( .A(n_518), .B(n_655), .Y(n_677) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g558 ( .A(n_519), .Y(n_558) );
AND2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_536), .Y(n_633) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OR2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g696 ( .A(n_530), .B(n_596), .Y(n_696) );
AND2x2_ASAP7_75t_L g710 ( .A(n_530), .B(n_532), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_531), .B(n_544), .Y(n_651) );
AND2x2_ASAP7_75t_L g698 ( .A(n_531), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g578 ( .A(n_532), .B(n_544), .Y(n_578) );
INVx1_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
AND2x2_ASAP7_75t_L g619 ( .A(n_532), .B(n_544), .Y(n_619) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_534), .A2(n_662), .B1(n_666), .B2(n_668), .C(n_669), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_537), .Y(n_534) );
AND2x2_ASAP7_75t_L g565 ( .A(n_535), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_538), .B(n_572), .Y(n_715) );
AOI322xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_557), .A3(n_558), .B1(n_559), .B2(n_565), .C1(n_567), .C2(n_574), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_556), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_543), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_543), .B(n_606), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_543), .A2(n_556), .B(n_630), .C(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_543), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_543), .B(n_600), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_543), .B(n_682), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_543), .B(n_710), .Y(n_709) );
BUFx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_544), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_544), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g671 ( .A(n_544), .B(n_558), .Y(n_671) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B(n_555), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_546), .A2(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g563 ( .A(n_548), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_555), .Y(n_564) );
INVx1_ASAP7_75t_L g646 ( .A(n_556), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_556), .A2(n_581), .A3(n_657), .B(n_659), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_556), .B(n_562), .Y(n_708) );
INVx1_ASAP7_75t_SL g569 ( .A(n_557), .Y(n_569) );
AND2x2_ASAP7_75t_L g602 ( .A(n_557), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g683 ( .A(n_557), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g568 ( .A(n_558), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
AND2x2_ASAP7_75t_L g620 ( .A(n_558), .B(n_573), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_558), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g712 ( .A(n_558), .B(n_660), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_560), .B(n_630), .Y(n_703) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g599 ( .A(n_562), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g617 ( .A(n_562), .Y(n_617) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_568), .B(n_570), .Y(n_567) );
OAI211xp5_ASAP7_75t_SL g611 ( .A1(n_569), .A2(n_612), .B(n_618), .C(n_634), .Y(n_611) );
OR2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_667), .Y(n_686) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g623 ( .A(n_571), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_571), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g592 ( .A(n_573), .B(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_582), .C(n_585), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g626 ( .A(n_578), .Y(n_626) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_581), .B(n_619), .Y(n_624) );
INVx1_ASAP7_75t_L g630 ( .A(n_581), .Y(n_630) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g589 ( .A(n_584), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g622 ( .A(n_584), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g684 ( .A(n_584), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_587), .B(n_589), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_587), .A2(n_598), .B(n_601), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B(n_597), .C(n_604), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_592), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_595), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g608 ( .A(n_596), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_598), .A2(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_603), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g628 ( .A(n_603), .Y(n_628) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_608), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g659 ( .A(n_610), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_616), .B(n_642), .Y(n_668) );
AND2x2_ASAP7_75t_L g681 ( .A(n_616), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g695 ( .A(n_616), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g705 ( .A(n_616), .B(n_643), .Y(n_705) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_621), .C(n_629), .Y(n_618) );
INVx1_ASAP7_75t_L g665 ( .A(n_619), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_627), .Y(n_621) );
OR2x2_ASAP7_75t_L g627 ( .A(n_623), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_623), .B(n_684), .Y(n_706) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g700 ( .A(n_633), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_640), .B1(n_643), .B2(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g718 ( .A(n_638), .Y(n_718) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g664 ( .A(n_642), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B(n_649), .C(n_656), .Y(n_645) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_664), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR5xp2_ASAP7_75t_L g674 ( .A(n_675), .B(n_693), .C(n_701), .D(n_707), .E(n_713), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_678), .B(n_680), .C(n_687), .Y(n_675) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B(n_685), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_690), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .B(n_700), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g716 ( .A(n_696), .Y(n_716) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g727 ( .A(n_720), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g747 ( .A(n_736), .Y(n_747) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_742), .B1(n_743), .B2(n_745), .Y(n_737) );
INVx1_ASAP7_75t_L g745 ( .A(n_738), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule