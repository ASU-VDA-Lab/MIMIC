module fake_jpeg_17431_n_125 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_13),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_11),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_22),
.B1(n_18),
.B2(n_23),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_53),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_16),
.B1(n_22),
.B2(n_1),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_16),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_44),
.C(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_26),
.C(n_17),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_54),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_23),
.CI(n_26),
.CON(n_49),
.SN(n_49)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_52),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_3),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_63),
.B(n_59),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_38),
.B1(n_36),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_78),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_50),
.B1(n_67),
.B2(n_80),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_64),
.C(n_55),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_42),
.C(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.C(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_94),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_57),
.C(n_51),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_51),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_50),
.C(n_81),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_66),
.C(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_68),
.B1(n_70),
.B2(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_71),
.B(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_93),
.C(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_117),
.B(n_95),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_102),
.C(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_111),
.B1(n_104),
.B2(n_112),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_113),
.B(n_108),
.C(n_109),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_121),
.B(n_119),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_114),
.C(n_87),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_124),
.C(n_106),
.Y(n_125)
);


endmodule