module fake_jpeg_11489_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_50),
.B1(n_66),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_52),
.B1(n_53),
.B2(n_64),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_53),
.Y(n_89)
);

NAND2x1p5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_49),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_50),
.B1(n_66),
.B2(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_79),
.B(n_86),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_63),
.B(n_57),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_63),
.B1(n_57),
.B2(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_107),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_53),
.B1(n_64),
.B2(n_52),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_60),
.B(n_1),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_0),
.B(n_2),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_91),
.B1(n_77),
.B2(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_3),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_122),
.B(n_125),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_6),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_127),
.B1(n_131),
.B2(n_14),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_8),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_11),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_30),
.A3(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_23),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_136),
.C(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_106),
.B1(n_12),
.B2(n_13),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_143),
.B1(n_145),
.B2(n_131),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_22),
.B(n_40),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_45),
.C(n_38),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_27),
.C(n_35),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_119),
.B1(n_113),
.B2(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.C(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_137),
.B(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.C(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_148),
.B1(n_140),
.B2(n_135),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_157),
.B(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_136),
.B1(n_133),
.B2(n_149),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_36),
.A3(n_31),
.B1(n_32),
.B2(n_148),
.C1(n_117),
.C2(n_119),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_117),
.Y(n_161)
);


endmodule