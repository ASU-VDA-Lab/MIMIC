module fake_jpeg_23967_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_27),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_64),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_12),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_14),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_40),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_24),
.B1(n_18),
.B2(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_19),
.B1(n_29),
.B2(n_6),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_12),
.B1(n_38),
.B2(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_81),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_84),
.B(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_47),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_61),
.B1(n_58),
.B2(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_107),
.B(n_71),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_106),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_46),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_90),
.B(n_74),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_73),
.C(n_70),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_126),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_112),
.B(n_117),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_106),
.B(n_104),
.C(n_107),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_95),
.B1(n_109),
.B2(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_103),
.B1(n_106),
.B2(n_118),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_115),
.B1(n_102),
.B2(n_101),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_105),
.B(n_97),
.C(n_110),
.D(n_79),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_101),
.C(n_70),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_76),
.B(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

OAI21x1_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_128),
.B(n_125),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_128),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_146),
.B(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_125),
.B1(n_78),
.B2(n_95),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_149),
.B(n_151),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_144),
.C(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_145),
.B(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_140),
.C(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_128),
.B1(n_143),
.B2(n_138),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_160),
.B(n_154),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_143),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_126),
.B1(n_155),
.B2(n_143),
.C(n_134),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_158),
.Y(n_164)
);


endmodule