module fake_jpeg_20610_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_41),
.Y(n_74)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_58),
.B1(n_77),
.B2(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_83),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_23),
.B1(n_19),
.B2(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_68),
.B1(n_76),
.B2(n_79),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_23),
.B1(n_19),
.B2(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_28),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_34),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_36),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_20),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_20),
.B1(n_29),
.B2(n_2),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_88),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_0),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_36),
.A2(n_0),
.B(n_1),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_4),
.C(n_5),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_108),
.B1(n_96),
.B2(n_100),
.Y(n_142)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_83),
.C(n_73),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_62),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_7),
.B(n_8),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_7),
.Y(n_111)
);

AO22x2_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_9),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_107),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_125),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_64),
.B(n_48),
.C(n_58),
.D(n_77),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_112),
.B(n_103),
.C(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_116),
.C(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_57),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_54),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_147),
.B(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_144),
.Y(n_153)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_145),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_52),
.B1(n_86),
.B2(n_78),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_142),
.B1(n_51),
.B2(n_78),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_96),
.A2(n_86),
.B1(n_52),
.B2(n_49),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_148),
.B1(n_93),
.B2(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_49),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_111),
.Y(n_145)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_67),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_60),
.B1(n_56),
.B2(n_51),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_154),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_112),
.B1(n_113),
.B2(n_117),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_130),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_97),
.B(n_90),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_158),
.B(n_167),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_97),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_146),
.C(n_134),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_110),
.B(n_57),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_116),
.B1(n_110),
.B2(n_12),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_166),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_144),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.C(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_9),
.C(n_11),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_183),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_193),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_137),
.A3(n_134),
.B1(n_130),
.B2(n_122),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_136),
.B1(n_122),
.B2(n_119),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_195),
.B(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_11),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_211),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_192),
.B1(n_194),
.B2(n_171),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_170),
.C(n_155),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_180),
.C(n_192),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_163),
.B1(n_153),
.B2(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_179),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_180),
.B(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_187),
.C(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_205),
.C(n_162),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_203),
.B1(n_178),
.B2(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_211),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_223),
.Y(n_239)
);

AOI321xp33_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_208),
.A3(n_204),
.B1(n_202),
.B2(n_209),
.C(n_201),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_233),
.C(n_225),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_196),
.C(n_157),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_220),
.C(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_239),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_217),
.Y(n_238)
);

OAI221xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_151),
.B1(n_164),
.B2(n_198),
.C(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_221),
.C(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_228),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_234),
.B(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.C(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_190),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_241),
.C(n_237),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_238),
.B(n_210),
.C(n_198),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_253),
.A2(n_254),
.B(n_182),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_228),
.B(n_189),
.Y(n_254)
);

AOI321xp33_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_250),
.A3(n_191),
.B1(n_182),
.B2(n_176),
.C(n_151),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);


endmodule