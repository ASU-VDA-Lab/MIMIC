module real_aes_2181_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g270 ( .A(n_0), .B(n_219), .Y(n_270) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_1), .A2(n_53), .B1(n_90), .B2(n_101), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_2), .A2(n_7), .B1(n_135), .B2(n_140), .Y(n_134) );
INVx1_ASAP7_75t_L g188 ( .A(n_3), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_4), .B(n_204), .Y(n_203) );
NAND2xp33_ASAP7_75t_SL g314 ( .A(n_5), .B(n_210), .Y(n_314) );
INVx1_ASAP7_75t_L g306 ( .A(n_6), .Y(n_306) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_8), .A2(n_18), .B1(n_90), .B2(n_98), .Y(n_97) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_9), .A2(n_11), .B1(n_171), .B2(n_172), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_9), .Y(n_171) );
AND2x2_ASAP7_75t_L g198 ( .A(n_10), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g172 ( .A(n_11), .Y(n_172) );
INVx2_ASAP7_75t_L g200 ( .A(n_12), .Y(n_200) );
AOI221x1_ASAP7_75t_L g309 ( .A1(n_13), .A2(n_212), .B1(n_310), .B2(n_312), .C(n_313), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_14), .B(n_204), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_15), .A2(n_212), .B(n_217), .Y(n_211) );
AOI221xp5_ASAP7_75t_SL g280 ( .A1(n_16), .A2(n_32), .B1(n_204), .B2(n_212), .C(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_17), .B(n_219), .Y(n_218) );
OAI221xp5_ASAP7_75t_L g180 ( .A1(n_18), .A2(n_53), .B1(n_56), .B2(n_181), .C(n_183), .Y(n_180) );
OR2x2_ASAP7_75t_L g201 ( .A(n_19), .B(n_68), .Y(n_201) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_19), .A2(n_68), .B(n_200), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_20), .B(n_221), .Y(n_297) );
INVxp67_ASAP7_75t_L g308 ( .A(n_21), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_22), .Y(n_102) );
AND2x2_ASAP7_75t_L g243 ( .A(n_23), .B(n_233), .Y(n_243) );
INVx3_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_25), .A2(n_44), .B1(n_124), .B2(n_128), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_26), .A2(n_54), .B1(n_160), .B2(n_164), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_27), .A2(n_63), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_27), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_27), .A2(n_212), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_28), .B(n_221), .Y(n_282) );
INVx1_ASAP7_75t_SL g91 ( .A(n_29), .Y(n_91) );
INVx1_ASAP7_75t_L g190 ( .A(n_30), .Y(n_190) );
AND2x2_ASAP7_75t_L g210 ( .A(n_30), .B(n_188), .Y(n_210) );
AND2x2_ASAP7_75t_L g213 ( .A(n_30), .B(n_214), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_31), .A2(n_61), .B1(n_145), .B2(n_148), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_33), .A2(n_60), .B1(n_212), .B2(n_257), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_34), .A2(n_71), .B1(n_154), .B2(n_157), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_35), .B(n_219), .Y(n_241) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_36), .A2(n_56), .B1(n_90), .B2(n_94), .Y(n_93) );
AND2x2_ASAP7_75t_L g273 ( .A(n_37), .B(n_233), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_38), .A2(n_42), .B1(n_115), .B2(n_119), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_39), .B(n_233), .Y(n_284) );
INVx1_ASAP7_75t_L g207 ( .A(n_40), .Y(n_207) );
INVx1_ASAP7_75t_L g216 ( .A(n_40), .Y(n_216) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_43), .B(n_204), .Y(n_242) );
AND2x2_ASAP7_75t_L g234 ( .A(n_45), .B(n_233), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_46), .B(n_221), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_47), .A2(n_80), .B1(n_166), .B2(n_167), .Y(n_79) );
INVx1_ASAP7_75t_L g166 ( .A(n_47), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_48), .B(n_219), .Y(n_230) );
AND2x2_ASAP7_75t_SL g298 ( .A(n_49), .B(n_199), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_50), .A2(n_212), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_51), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_52), .B(n_248), .Y(n_261) );
INVxp33_ASAP7_75t_L g185 ( .A(n_53), .Y(n_185) );
INVx1_ASAP7_75t_L g209 ( .A(n_55), .Y(n_209) );
INVx1_ASAP7_75t_L g214 ( .A(n_55), .Y(n_214) );
INVxp67_ASAP7_75t_L g184 ( .A(n_56), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_57), .A2(n_80), .B1(n_167), .B2(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_57), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_58), .B(n_204), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_59), .A2(n_62), .B1(n_204), .B2(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g175 ( .A(n_63), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_64), .B(n_219), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_65), .B(n_219), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_66), .A2(n_69), .B1(n_104), .B2(n_109), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_67), .A2(n_212), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_70), .B(n_221), .Y(n_229) );
INVxp67_ASAP7_75t_L g311 ( .A(n_72), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_73), .B(n_204), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_74), .B(n_221), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_75), .A2(n_212), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g509 ( .A(n_75), .Y(n_509) );
BUFx2_ASAP7_75t_SL g182 ( .A(n_76), .Y(n_182) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_177), .B1(n_191), .B2(n_505), .C(n_506), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_168), .Y(n_78) );
INVxp67_ASAP7_75t_SL g167 ( .A(n_80), .Y(n_167) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_80), .Y(n_510) );
AND2x4_ASAP7_75t_L g80 ( .A(n_81), .B(n_132), .Y(n_80) );
NOR2xp67_ASAP7_75t_L g81 ( .A(n_82), .B(n_113), .Y(n_81) );
OAI21xp5_ASAP7_75t_SL g82 ( .A1(n_83), .A2(n_102), .B(n_103), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx4_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
INVx6_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x4_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g130 ( .A(n_87), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_88), .Y(n_112) );
INVx2_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
OAI22x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_90), .Y(n_101) );
INVx2_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
AND2x2_ASAP7_75t_L g126 ( .A(n_93), .B(n_127), .Y(n_126) );
BUFx2_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
AND2x2_ASAP7_75t_L g147 ( .A(n_95), .B(n_126), .Y(n_147) );
AND2x4_ASAP7_75t_L g156 ( .A(n_95), .B(n_107), .Y(n_156) );
AND2x4_ASAP7_75t_L g163 ( .A(n_95), .B(n_151), .Y(n_163) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x4_ASAP7_75t_L g106 ( .A(n_97), .B(n_99), .Y(n_106) );
AND2x2_ASAP7_75t_L g111 ( .A(n_97), .B(n_100), .Y(n_111) );
INVx1_ASAP7_75t_L g118 ( .A(n_97), .Y(n_118) );
INVxp67_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g117 ( .A(n_100), .B(n_118), .Y(n_117) );
BUFx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x4_ASAP7_75t_L g125 ( .A(n_106), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g165 ( .A(n_106), .B(n_151), .Y(n_165) );
AND2x2_ASAP7_75t_L g116 ( .A(n_107), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g151 ( .A(n_108), .B(n_127), .Y(n_151) );
BUFx12f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x4_ASAP7_75t_L g142 ( .A(n_111), .B(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g158 ( .A(n_111), .B(n_151), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_123), .Y(n_113) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g139 ( .A(n_117), .B(n_126), .Y(n_139) );
AND2x4_ASAP7_75t_L g150 ( .A(n_117), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_118), .Y(n_122) );
BUFx4f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx6_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_152), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_144), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_159), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx8_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_167), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B1(n_173), .B2(n_176), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_173), .Y(n_176) );
CKINVDCx14_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
AND3x1_ASAP7_75t_SL g179 ( .A(n_180), .B(n_186), .C(n_189), .Y(n_179) );
INVxp67_ASAP7_75t_L g514 ( .A(n_180), .Y(n_514) );
CKINVDCx8_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_186), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_186), .A2(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g253 ( .A(n_187), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_SL g520 ( .A(n_187), .B(n_189), .Y(n_520) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g215 ( .A(n_188), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_189), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g258 ( .A(n_190), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_435), .Y(n_192) );
NOR4xp25_ASAP7_75t_SL g193 ( .A(n_194), .B(n_328), .C(n_372), .D(n_399), .Y(n_193) );
OAI221xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_289), .B1(n_299), .B2(n_316), .C(n_318), .Y(n_194) );
AOI32xp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_244), .A3(n_262), .B1(n_274), .B2(n_285), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_196), .B(n_471), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_196), .A2(n_441), .B1(n_499), .B2(n_502), .Y(n_498) );
AND2x4_ASAP7_75t_SL g196 ( .A(n_197), .B(n_224), .Y(n_196) );
INVx5_ASAP7_75t_L g288 ( .A(n_197), .Y(n_288) );
OR2x2_ASAP7_75t_L g317 ( .A(n_197), .B(n_287), .Y(n_317) );
AND2x4_ASAP7_75t_L g319 ( .A(n_197), .B(n_236), .Y(n_319) );
INVx2_ASAP7_75t_L g334 ( .A(n_197), .Y(n_334) );
OR2x2_ASAP7_75t_L g346 ( .A(n_197), .B(n_245), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_197), .B(n_235), .Y(n_353) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_197), .B(n_276), .Y(n_395) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_197), .Y(n_452) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AND2x4_ASAP7_75t_L g223 ( .A(n_200), .B(n_201), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_211), .B(n_223), .Y(n_202) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_210), .Y(n_204) );
INVx1_ASAP7_75t_L g315 ( .A(n_205), .Y(n_315) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
AND2x6_ASAP7_75t_L g219 ( .A(n_206), .B(n_214), .Y(n_219) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g221 ( .A(n_208), .B(n_216), .Y(n_221) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx5_ASAP7_75t_L g222 ( .A(n_210), .Y(n_222) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_212), .Y(n_505) );
AND2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
BUFx3_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
INVx2_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
AND2x4_ASAP7_75t_L g257 ( .A(n_215), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_222), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_222), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_222), .A2(n_270), .B(n_271), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_222), .A2(n_282), .B(n_283), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_222), .A2(n_296), .B(n_297), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_223), .B(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_223), .B(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_223), .B(n_311), .Y(n_310) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_223), .B(n_314), .C(n_315), .Y(n_313) );
INVx3_ASAP7_75t_SL g347 ( .A(n_224), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_224), .B(n_288), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g481 ( .A1(n_224), .A2(n_352), .A3(n_382), .B1(n_412), .B2(n_447), .Y(n_481) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
AND2x2_ASAP7_75t_L g321 ( .A(n_225), .B(n_245), .Y(n_321) );
OR2x2_ASAP7_75t_L g337 ( .A(n_225), .B(n_236), .Y(n_337) );
INVx1_ASAP7_75t_L g360 ( .A(n_225), .Y(n_360) );
INVx2_ASAP7_75t_L g376 ( .A(n_225), .Y(n_376) );
AND2x2_ASAP7_75t_L g413 ( .A(n_225), .B(n_276), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_225), .B(n_236), .Y(n_432) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_225), .Y(n_501) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_234), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_232), .A2(n_237), .B(n_243), .Y(n_236) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_232), .A2(n_237), .B(n_243), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_233), .Y(n_232) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_233), .A2(n_280), .B(n_284), .Y(n_279) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g468 ( .A(n_236), .B(n_245), .Y(n_468) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_236), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
OR2x2_ASAP7_75t_L g316 ( .A(n_244), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g322 ( .A(n_244), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_244), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g497 ( .A(n_244), .B(n_366), .Y(n_497) );
BUFx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g426 ( .A(n_245), .B(n_376), .Y(n_426) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B(n_261), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_248), .A2(n_293), .B(n_294), .Y(n_292) );
BUFx4f_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g266 ( .A(n_249), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_252), .A2(n_257), .B1(n_305), .B2(n_307), .Y(n_304) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g525 ( .A(n_253), .Y(n_525) );
INVx1_ASAP7_75t_L g524 ( .A(n_255), .Y(n_524) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_262), .B(n_393), .Y(n_495) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_263), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_264), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
AND2x2_ASAP7_75t_L g326 ( .A(n_264), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_264), .B(n_302), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_264), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g384 ( .A(n_264), .Y(n_384) );
OR2x2_ASAP7_75t_L g403 ( .A(n_264), .B(n_330), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_264), .Y(n_410) );
NOR2xp33_ASAP7_75t_R g462 ( .A(n_264), .B(n_291), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_264), .B(n_303), .Y(n_466) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_273), .Y(n_265) );
INVx4_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_272), .Y(n_267) );
AOI32xp33_ASAP7_75t_L g489 ( .A1(n_274), .A2(n_325), .A3(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g356 ( .A(n_276), .Y(n_356) );
AND2x4_ASAP7_75t_L g375 ( .A(n_276), .B(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_276), .B(n_347), .Y(n_404) );
OR2x2_ASAP7_75t_L g458 ( .A(n_276), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g416 ( .A(n_277), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g474 ( .A(n_277), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_278), .B(n_291), .Y(n_440) );
AND2x2_ASAP7_75t_L g477 ( .A(n_278), .B(n_443), .Y(n_477) );
INVx2_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
INVx2_ASAP7_75t_L g330 ( .A(n_279), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_279), .B(n_291), .Y(n_350) );
INVx1_ASAP7_75t_L g381 ( .A(n_279), .Y(n_381) );
OR2x2_ASAP7_75t_L g407 ( .A(n_279), .B(n_291), .Y(n_407) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_279), .Y(n_459) );
BUFx3_ASAP7_75t_L g488 ( .A(n_279), .Y(n_488) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g357 ( .A(n_286), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_286), .B(n_375), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_286), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_287), .B(n_360), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_287), .A2(n_356), .B(n_374), .Y(n_389) );
OAI32xp33_ASAP7_75t_L g411 ( .A1(n_288), .A2(n_412), .A3(n_414), .B1(n_416), .B2(n_418), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_288), .B(n_375), .Y(n_484) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g417 ( .A(n_290), .Y(n_417) );
NOR2x1p5_ASAP7_75t_L g487 ( .A(n_290), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g301 ( .A(n_291), .B(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_SL g325 ( .A(n_291), .B(n_303), .Y(n_325) );
OR2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
AND2x2_ASAP7_75t_L g382 ( .A(n_291), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g393 ( .A(n_291), .B(n_303), .Y(n_393) );
OR2x2_ASAP7_75t_L g455 ( .A(n_291), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g472 ( .A(n_291), .B(n_403), .Y(n_472) );
INVx1_ASAP7_75t_L g504 ( .A(n_291), .Y(n_504) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_298), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_300), .B(n_381), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_301), .B(n_415), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g419 ( .A1(n_301), .A2(n_420), .B1(n_425), .B2(n_427), .C1(n_430), .C2(n_433), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_301), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g447 ( .A(n_301), .B(n_326), .Y(n_447) );
AND2x2_ASAP7_75t_L g409 ( .A(n_302), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g424 ( .A(n_302), .B(n_329), .Y(n_424) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_303), .B(n_330), .Y(n_362) );
AND2x4_ASAP7_75t_L g383 ( .A(n_303), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g443 ( .A(n_303), .B(n_364), .Y(n_443) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_309), .Y(n_303) );
INVx1_ASAP7_75t_SL g323 ( .A(n_317), .Y(n_323) );
NAND2xp33_ASAP7_75t_SL g492 ( .A(n_317), .B(n_347), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_322), .C(n_324), .Y(n_318) );
INVx2_ASAP7_75t_SL g369 ( .A(n_319), .Y(n_369) );
AND2x2_ASAP7_75t_L g373 ( .A(n_320), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_321), .B(n_369), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_321), .A2(n_359), .B(n_395), .C(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g471 ( .A(n_321), .B(n_452), .Y(n_471) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x4_ASAP7_75t_L g370 ( .A(n_325), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g475 ( .A(n_325), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B(n_338), .C(n_365), .Y(n_328) );
INVx2_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
OR2x2_ASAP7_75t_L g387 ( .A(n_329), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_333), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g425 ( .A(n_333), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_333), .B(n_413), .Y(n_479) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_335), .A2(n_438), .B1(n_439), .B2(n_441), .C1(n_444), .C2(n_447), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_336), .A2(n_401), .B1(n_404), .B2(n_405), .C(n_411), .Y(n_400) );
AND2x2_ASAP7_75t_L g438 ( .A(n_336), .B(n_395), .Y(n_438) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp33_ASAP7_75t_SL g351 ( .A(n_337), .B(n_352), .Y(n_351) );
AOI221x1_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_348), .B2(n_351), .C(n_354), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g491 ( .A(n_341), .B(n_429), .Y(n_491) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g349 ( .A(n_342), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
OAI32xp33_ASAP7_75t_L g457 ( .A1(n_347), .A2(n_388), .A3(n_458), .B1(n_460), .B2(n_464), .Y(n_457) );
OAI21xp33_ASAP7_75t_SL g476 ( .A1(n_348), .A2(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_361), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
OR2x2_ASAP7_75t_L g358 ( .A(n_356), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g431 ( .A(n_356), .B(n_432), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_360), .A2(n_386), .B1(n_389), .B2(n_390), .C(n_394), .Y(n_385) );
INVx1_ASAP7_75t_L g461 ( .A(n_360), .Y(n_461) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_360), .Y(n_467) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_369), .B(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_377), .B(n_385), .Y(n_372) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_376), .Y(n_446) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_379), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g398 ( .A(n_381), .Y(n_398) );
INVx1_ASAP7_75t_L g388 ( .A(n_383), .Y(n_388) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_383), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_383), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_383), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g402 ( .A(n_393), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_398), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_400), .B(n_419), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g415 ( .A(n_403), .Y(n_415) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_SL g429 ( .A(n_407), .Y(n_429) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_409), .B(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_410), .Y(n_423) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g434 ( .A(n_426), .Y(n_434) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
NOR4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_469), .C(n_480), .D(n_493), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_448), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_438), .A2(n_449), .B(n_454), .C(n_457), .Y(n_448) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_453), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g460 ( .A1(n_451), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_468), .B(n_500), .Y(n_499) );
OAI221xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_472), .B1(n_473), .B2(n_474), .C(n_476), .Y(n_469) );
INVx1_ASAP7_75t_SL g473 ( .A(n_471), .Y(n_473) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_482), .C(n_489), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp33_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OAI222xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_509), .B1(n_511), .B2(n_515), .C1(n_518), .C2(n_521), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
endmodule