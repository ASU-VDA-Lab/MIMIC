module real_jpeg_21194_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_2),
.B1(n_38),
.B2(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_38),
.B1(n_60),
.B2(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_7),
.B1(n_40),
.B2(n_57),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_40),
.B(n_63),
.C(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_46),
.B(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_3),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_61),
.B(n_62),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_34),
.B(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_58),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_57),
.B(n_59),
.C(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_57),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_36)
);

BUFx3_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_107),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_106),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_93),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_42),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_21),
.A2(n_22),
.B1(n_47),
.B2(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_21),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_22),
.A2(n_25),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_22),
.B(n_40),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_29),
.A2(n_30),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_29),
.A2(n_30),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_30),
.B(n_87),
.C(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_30),
.B(n_158),
.C(n_165),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_31),
.B(n_36),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_33),
.A2(n_34),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_34),
.A2(n_35),
.B(n_40),
.C(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_36),
.B(n_40),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_40),
.B(n_73),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_40),
.A2(n_61),
.B(n_75),
.C(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_44),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_48),
.A2(n_49),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_48),
.A2(n_49),
.B1(n_101),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_49),
.B(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_49),
.B(n_101),
.C(n_143),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B(n_52),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_68),
.B2(n_69),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_54),
.A2(n_55),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_101),
.C(n_103),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B(n_64),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_58),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_73),
.B(n_74),
.C(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_74),
.Y(n_78)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_92),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_89),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_137),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2x1_ASAP7_75t_R g127 ( 
.A(n_87),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_128),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_87),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_89),
.A2(n_90),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_126),
.C(n_161),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.C(n_100),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_95),
.B(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_100),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_101),
.A2(n_103),
.B1(n_153),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_103),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_182),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_178),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_167),
.B(n_177),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_155),
.B(n_166),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_140),
.B(n_154),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_131),
.B(n_139),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_122),
.B(n_130),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B(n_129),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_151),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_151),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);


endmodule