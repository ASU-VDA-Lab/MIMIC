module fake_aes_10314_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx4_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
BUFx2_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_14), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AOI22xp5_ASAP7_75t_SL g23 ( .A1(n_18), .A2(n_13), .B1(n_12), .B2(n_16), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_21), .B(n_13), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_18), .B1(n_21), .B2(n_19), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_23), .B(n_18), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_18), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B1(n_18), .B2(n_21), .Y(n_29) );
OAI21xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_19), .B(n_20), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_20), .B1(n_19), .B2(n_21), .C(n_12), .Y(n_31) );
OAI221xp5_ASAP7_75t_SL g32 ( .A1(n_29), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_3), .Y(n_32) );
AOI221xp5_ASAP7_75t_SL g33 ( .A1(n_30), .A2(n_1), .B1(n_2), .B2(n_4), .C(n_16), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
INVxp33_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g38 ( .A(n_35), .Y(n_38) );
AOI222xp33_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_8), .B1(n_9), .B2(n_11), .C1(n_34), .C2(n_38), .Y(n_39) );
endmodule