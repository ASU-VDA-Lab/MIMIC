module fake_jpeg_31380_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_11),
.B(n_14),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_79),
.B(n_81),
.Y(n_83)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_20),
.B1(n_45),
.B2(n_44),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_57),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_72),
.B(n_4),
.C(n_5),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_96),
.Y(n_108)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_74),
.B1(n_51),
.B2(n_65),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_114),
.B1(n_113),
.B2(n_109),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_65),
.B1(n_64),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_28),
.B1(n_43),
.B2(n_41),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_54),
.B(n_56),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_105),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_58),
.B(n_53),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_6),
.B(n_7),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_63),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_3),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_113),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_67),
.B(n_71),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_117),
.B(n_9),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_55),
.B1(n_59),
.B2(n_69),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_97),
.B1(n_78),
.B2(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_110),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_78),
.B(n_5),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_19),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_12),
.C(n_15),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_125),
.B1(n_16),
.B2(n_17),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_7),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_8),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_131),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_9),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_134),
.B(n_12),
.C(n_14),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

OAI322xp33_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_124),
.A3(n_129),
.B1(n_135),
.B2(n_134),
.C1(n_120),
.C2(n_37),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_27),
.C(n_29),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_133),
.C(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_150),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_133),
.C(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_145),
.C(n_143),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_137),
.B1(n_138),
.B2(n_146),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_153),
.B(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_151),
.Y(n_157)
);

OAI331xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_138),
.A3(n_147),
.B1(n_137),
.B2(n_34),
.B3(n_36),
.C1(n_47),
.Y(n_158)
);

AOI221xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_136),
.B1(n_32),
.B2(n_33),
.C(n_31),
.Y(n_159)
);


endmodule