module fake_netlist_6_1585_n_13275 (n_992, n_2542, n_1671, n_1, n_2817, n_801, n_1613, n_1234, n_1458, n_2576, n_1199, n_1674, n_741, n_1027, n_1351, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_2157, n_2332, n_212, n_700, n_50, n_1307, n_2003, n_1038, n_578, n_1581, n_1003, n_365, n_168, n_1237, n_1061, n_2353, n_2534, n_1357, n_1853, n_77, n_783, n_2451, n_1738, n_2243, n_798, n_188, n_1575, n_1854, n_2324, n_1923, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_2260, n_677, n_1708, n_805, n_1151, n_396, n_1739, n_350, n_78, n_2051, n_2317, n_1380, n_2359, n_442, n_480, n_142, n_2847, n_1402, n_2557, n_1688, n_1691, n_1975, n_1009, n_1743, n_62, n_1930, n_2405, n_1160, n_883, n_2647, n_1238, n_1991, n_2570, n_2179, n_2386, n_1724, n_1032, n_2336, n_1247, n_1547, n_2521, n_1553, n_893, n_1099, n_2491, n_1264, n_1192, n_471, n_1844, n_424, n_1700, n_1555, n_1415, n_2211, n_1370, n_1786, n_369, n_287, n_2382, n_2672, n_2291, n_415, n_830, n_2299, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_1371, n_2886, n_200, n_1985, n_447, n_2838, n_2184, n_1803, n_1172, n_852, n_2509, n_71, n_229, n_2513, n_1590, n_2645, n_1532, n_2313, n_2628, n_1393, n_1517, n_1867, n_1704, n_1078, n_250, n_544, n_1711, n_2247, n_1140, n_2630, n_1444, n_1670, n_1603, n_2344, n_1579, n_35, n_2365, n_2470, n_2321, n_1263, n_2019, n_836, n_375, n_2074, n_2447, n_522, n_2919, n_2129, n_2340, n_1261, n_945, n_2286, n_1649, n_2018, n_2094, n_1903, n_1511, n_1143, n_2356, n_2399, n_1422, n_1232, n_1772, n_1572, n_616, n_658, n_1874, n_1119, n_2865, n_2825, n_2013, n_428, n_1433, n_1902, n_1842, n_1620, n_2044, n_1954, n_1735, n_2510, n_1541, n_1300, n_641, n_2480, n_2739, n_822, n_693, n_1313, n_2791, n_1056, n_2212, n_758, n_516, n_1455, n_2418, n_2864, n_1163, n_2729, n_1180, n_2256, n_2582, n_943, n_1798, n_1550, n_2703, n_491, n_2786, n_1591, n_42, n_772, n_2806, n_1344, n_2730, n_2495, n_666, n_371, n_940, n_770, n_567, n_1781, n_1971, n_2058, n_2090, n_2603, n_405, n_213, n_2660, n_538, n_2173, n_2004, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_1345, n_1820, n_2873, n_494, n_539, n_493, n_155, n_2880, n_2394, n_2108, n_45, n_454, n_1421, n_2836, n_1936, n_638, n_1404, n_1211, n_2124, n_381, n_2378, n_887, n_1660, n_1961, n_112, n_1280, n_713, n_2655, n_1400, n_2625, n_2843, n_126, n_1467, n_58, n_976, n_2155, n_224, n_2686, n_48, n_1445, n_2364, n_2551, n_1526, n_1560, n_734, n_1088, n_1894, n_196, n_1231, n_2599, n_1978, n_2085, n_917, n_574, n_9, n_2370, n_2612, n_907, n_6, n_1446, n_14, n_2591, n_659, n_1815, n_2214, n_407, n_913, n_1658, n_2593, n_808, n_867, n_1230, n_473, n_1193, n_1967, n_1054, n_559, n_2613, n_1333, n_2496, n_44, n_2708, n_1648, n_1911, n_1956, n_163, n_1644, n_2011, n_2725, n_2277, n_1558, n_1732, n_281, n_551, n_699, n_1986, n_2300, n_564, n_2397, n_451, n_824, n_279, n_686, n_757, n_594, n_1641, n_2113, n_1918, n_2190, n_2907, n_577, n_166, n_2735, n_1843, n_619, n_2268, n_1367, n_1336, n_521, n_2778, n_2850, n_572, n_395, n_813, n_1909, n_2080, n_1481, n_323, n_606, n_1441, n_818, n_1123, n_1309, n_92, n_2104, n_513, n_645, n_1381, n_331, n_1699, n_916, n_2093, n_2633, n_483, n_102, n_2207, n_1970, n_2770, n_608, n_261, n_2101, n_2696, n_630, n_2059, n_32, n_2198, n_541, n_512, n_2669, n_2073, n_2273, n_121, n_433, n_2546, n_792, n_2522, n_476, n_2792, n_2, n_1328, n_1957, n_2917, n_219, n_2616, n_1907, n_2529, n_264, n_263, n_1162, n_860, n_1530, n_788, n_939, n_1543, n_821, n_2811, n_938, n_1302, n_1068, n_1599, n_329, n_982, n_2674, n_2832, n_549, n_1762, n_1910, n_1075, n_408, n_932, n_2831, n_61, n_237, n_1876, n_1895, n_2123, n_1697, n_2143, n_243, n_979, n_1873, n_905, n_1866, n_1680, n_117, n_175, n_322, n_993, n_2692, n_689, n_2031, n_354, n_2130, n_1330, n_1413, n_1605, n_2228, n_134, n_1988, n_1278, n_547, n_2455, n_2876, n_558, n_2654, n_2469, n_1064, n_1396, n_634, n_2355, n_136, n_966, n_2908, n_764, n_2751, n_2764, n_1663, n_2895, n_2009, n_692, n_733, n_1793, n_1233, n_1289, n_2714, n_2245, n_487, n_241, n_30, n_2068, n_1107, n_2866, n_2457, n_1014, n_1290, n_1703, n_2580, n_882, n_2176, n_2072, n_1354, n_2821, n_586, n_423, n_1865, n_1875, n_1701, n_2459, n_318, n_1111, n_1713, n_715, n_2678, n_1251, n_1265, n_2711, n_88, n_1726, n_1950, n_530, n_1563, n_1912, n_277, n_2434, n_1982, n_2878, n_618, n_1297, n_1662, n_1312, n_199, n_1167, n_1359, n_2818, n_2428, n_674, n_871, n_922, n_268, n_1335, n_1760, n_1927, n_210, n_2028, n_1069, n_2664, n_5, n_1664, n_1722, n_612, n_2641, n_178, n_247, n_1165, n_355, n_702, n_347, n_2008, n_2749, n_2192, n_2254, n_2345, n_1926, n_1175, n_328, n_1386, n_2311, n_1896, n_429, n_1747, n_1012, n_195, n_780, n_675, n_2624, n_903, n_1540, n_1977, n_1802, n_1504, n_2350, n_2804, n_2453, n_286, n_254, n_2193, n_2676, n_1655, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_1801, n_1886, n_2092, n_2347, n_1654, n_816, n_1157, n_1750, n_1462, n_1188, n_1752, n_877, n_1813, n_2514, n_2206, n_604, n_2810, n_2319, n_2519, n_825, n_728, n_2916, n_1063, n_1588, n_2467, n_26, n_2602, n_2468, n_55, n_267, n_1124, n_1624, n_515, n_2096, n_1965, n_2476, n_598, n_696, n_1515, n_961, n_437, n_1082, n_1317, n_2733, n_2824, n_593, n_514, n_687, n_697, n_890, n_637, n_2377, n_295, n_701, n_2178, n_950, n_388, n_190, n_2812, n_484, n_2644, n_2036, n_2152, n_1709, n_2652, n_2411, n_2525, n_1825, n_2393, n_1757, n_1796, n_170, n_2657, n_1792, n_891, n_2067, n_2136, n_2409, n_2082, n_2252, n_1412, n_2497, n_2687, n_949, n_1630, n_678, n_2887, n_283, n_2075, n_2194, n_2619, n_91, n_2763, n_2762, n_1987, n_507, n_968, n_909, n_1369, n_881, n_2271, n_1008, n_760, n_1546, n_2583, n_590, n_63, n_2606, n_362, n_148, n_2279, n_161, n_22, n_462, n_1033, n_1052, n_2794, n_1296, n_2663, n_1990, n_2391, n_304, n_2431, n_694, n_2150, n_1294, n_1420, n_125, n_1634, n_2078, n_297, n_595, n_627, n_1767, n_1779, n_524, n_1465, n_342, n_2622, n_1858, n_1044, n_2658, n_2665, n_2165, n_2133, n_1712, n_1391, n_449, n_131, n_1523, n_2558, n_2750, n_2775, n_1208, n_2893, n_1164, n_1295, n_1627, n_2728, n_2349, n_2684, n_2712, n_1072, n_1527, n_1495, n_1438, n_495, n_815, n_1100, n_585, n_1487, n_2691, n_840, n_2913, n_874, n_1756, n_1128, n_2493, n_382, n_673, n_2230, n_2705, n_1969, n_2690, n_1071, n_1067, n_1565, n_1493, n_2145, n_1968, n_898, n_255, n_284, n_1952, n_865, n_2573, n_2646, n_925, n_1932, n_1101, n_15, n_1026, n_1880, n_2535, n_2631, n_38, n_289, n_1364, n_2436, n_615, n_2870, n_1249, n_2706, n_59, n_1293, n_2693, n_1127, n_1512, n_2151, n_1451, n_320, n_108, n_639, n_963, n_794, n_2767, n_727, n_894, n_1839, n_2341, n_685, n_1765, n_353, n_2707, n_605, n_1514, n_1863, n_826, n_1646, n_872, n_1139, n_1714, n_86, n_104, n_718, n_1018, n_1521, n_1366, n_542, n_847, n_644, n_682, n_851, n_2537, n_2897, n_305, n_72, n_2554, n_996, n_532, n_173, n_1308, n_2089, n_1376, n_1513, n_2747, n_413, n_791, n_1913, n_510, n_837, n_2097, n_79, n_2170, n_1488, n_2853, n_1808, n_948, n_2517, n_2713, n_704, n_2148, n_977, n_2339, n_1005, n_1947, n_2765, n_2861, n_536, n_1788, n_1999, n_2731, n_622, n_147, n_2590, n_2643, n_1469, n_2060, n_2608, n_1838, n_2638, n_1835, n_1766, n_1776, n_1959, n_2002, n_581, n_2650, n_2138, n_765, n_432, n_987, n_1492, n_2414, n_1340, n_1771, n_2316, n_631, n_720, n_153, n_842, n_2262, n_1707, n_2239, n_1432, n_156, n_145, n_2208, n_843, n_656, n_989, n_2604, n_2407, n_1277, n_2816, n_797, n_2689, n_1473, n_2191, n_1723, n_2717, n_1246, n_1878, n_2574, n_899, n_189, n_738, n_2012, n_1304, n_1035, n_294, n_2842, n_499, n_2675, n_1426, n_705, n_11, n_1004, n_1176, n_2134, n_1529, n_2335, n_2473, n_1022, n_614, n_529, n_2069, n_2307, n_2362, n_425, n_684, n_2539, n_2667, n_2698, n_1431, n_1615, n_1474, n_1571, n_1809, n_1577, n_2297, n_1181, n_2119, n_1822, n_37, n_486, n_947, n_1117, n_2489, n_1087, n_1448, n_1992, n_648, n_657, n_1049, n_2771, n_2445, n_2057, n_2103, n_2605, n_1666, n_2772, n_1505, n_803, n_290, n_118, n_1717, n_926, n_1817, n_2449, n_927, n_2610, n_1849, n_2848, n_919, n_2868, n_1698, n_478, n_2231, n_929, n_107, n_2520, n_1228, n_417, n_2857, n_446, n_89, n_1568, n_1490, n_2372, n_777, n_1299, n_272, n_2896, n_526, n_2718, n_2639, n_1183, n_1436, n_2898, n_2251, n_1384, n_69, n_2494, n_2501, n_2238, n_293, n_2368, n_53, n_458, n_1070, n_2403, n_2837, n_998, n_16, n_717, n_1665, n_18, n_2524, n_154, n_1383, n_2460, n_1178, n_98, n_2127, n_1424, n_2338, n_1073, n_1000, n_796, n_252, n_1195, n_2137, n_1626, n_1507, n_2482, n_184, n_552, n_2532, n_1358, n_1811, n_1388, n_216, n_2481, n_912, n_1857, n_1519, n_2144, n_745, n_1284, n_1604, n_2296, n_2424, n_1142, n_2849, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1774, n_2354, n_2682, n_2589, n_1395, n_2110, n_2199, n_2661, n_731, n_2877, n_1502, n_1659, n_1955, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_2442, n_312, n_1791, n_1368, n_66, n_1418, n_958, n_292, n_1250, n_100, n_1137, n_1897, n_2064, n_880, n_2053, n_2259, n_2121, n_2773, n_2545, n_889, n_2432, n_2710, n_150, n_1478, n_589, n_1310, n_819, n_2294, n_1363, n_2581, n_1334, n_1942, n_1966, n_767, n_1314, n_600, n_964, n_831, n_1837, n_2218, n_2788, n_477, n_2435, n_954, n_864, n_2504, n_2797, n_2623, n_1110, n_2213, n_1410, n_399, n_2389, n_1440, n_124, n_2132, n_2892, n_2063, n_1382, n_1534, n_1564, n_1736, n_211, n_2748, n_1483, n_1834, n_2331, n_1372, n_231, n_2292, n_2860, n_2330, n_40, n_1457, n_505, n_1719, n_319, n_1339, n_1787, n_2701, n_2475, n_537, n_2511, n_1993, n_2281, n_1427, n_311, n_2416, n_2745, n_2617, n_2776, n_1466, n_10, n_403, n_1919, n_1080, n_723, n_1877, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1939, n_2030, n_1769, n_1220, n_2323, n_1893, n_556, n_2784, n_2209, n_2301, n_162, n_2387, n_1755, n_1602, n_2421, n_1136, n_2618, n_2025, n_2357, n_2846, n_2464, n_128, n_1125, n_970, n_2488, n_2224, n_1980, n_642, n_995, n_276, n_1159, n_2329, n_1092, n_2237, n_441, n_221, n_1060, n_1951, n_2250, n_444, n_146, n_1252, n_1784, n_1223, n_303, n_511, n_193, n_1286, n_1773, n_1775, n_2115, n_2410, n_2552, n_1053, n_2374, n_416, n_1681, n_520, n_418, n_1093, n_113, n_1783, n_1533, n_1597, n_2780, n_4, n_266, n_296, n_2596, n_2274, n_775, n_651, n_1153, n_439, n_1618, n_217, n_518, n_1531, n_2828, n_1185, n_453, n_215, n_2384, n_1745, n_914, n_759, n_2724, n_1831, n_426, n_317, n_2585, n_2621, n_1653, n_2352, n_1679, n_1625, n_90, n_2601, n_2160, n_54, n_1453, n_2146, n_2226, n_2131, n_488, n_2502, n_2801, n_497, n_2920, n_773, n_1901, n_920, n_99, n_1374, n_2556, n_2648, n_1315, n_1647, n_13, n_2575, n_2754, n_1224, n_2783, n_2306, n_1614, n_1459, n_1892, n_1933, n_2462, n_1135, n_1169, n_1179, n_2889, n_401, n_324, n_1617, n_335, n_1470, n_2550, n_463, n_1243, n_848, n_120, n_2732, n_301, n_274, n_1096, n_2249, n_1091, n_1917, n_2000, n_1580, n_2227, n_2270, n_2822, n_1425, n_36, n_1881, n_1267, n_1281, n_1806, n_983, n_2023, n_427, n_2572, n_2204, n_1520, n_496, n_2720, n_2159, n_906, n_1390, n_688, n_2289, n_1077, n_1733, n_2315, n_1419, n_2863, n_351, n_259, n_1731, n_177, n_2158, n_2087, n_1855, n_1636, n_1437, n_2135, n_1645, n_1832, n_385, n_1687, n_1439, n_2328, n_1323, n_2859, n_2202, n_858, n_2049, n_1331, n_613, n_736, n_2627, n_501, n_956, n_960, n_2276, n_663, n_856, n_2803, n_2100, n_379, n_778, n_1668, n_2777, n_1134, n_2830, n_2781, n_410, n_1129, n_554, n_602, n_1696, n_2829, n_1995, n_1594, n_2181, n_664, n_1869, n_171, n_2911, n_1764, n_169, n_1429, n_2826, n_1610, n_1889, n_2379, n_435, n_1905, n_2016, n_2343, n_793, n_326, n_587, n_1593, n_580, n_762, n_1030, n_1202, n_1937, n_465, n_1790, n_1778, n_1635, n_1079, n_341, n_2515, n_1744, n_828, n_2139, n_2142, n_607, n_316, n_419, n_28, n_1551, n_2448, n_1103, n_2875, n_2555, n_144, n_2219, n_1203, n_2851, n_820, n_2327, n_951, n_106, n_2201, n_725, n_952, n_999, n_358, n_1254, n_160, n_2841, n_2420, n_186, n_0, n_368, n_575, n_994, n_2263, n_2304, n_1508, n_2487, n_732, n_974, n_2240, n_392, n_2278, n_2656, n_2538, n_724, n_2597, n_2375, n_1934, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_1728, n_557, n_2756, n_1871, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1661, n_1275, n_2884, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_421, n_1468, n_2855, n_1859, n_2102, n_2563, n_238, n_1095, n_2024, n_1595, n_202, n_2156, n_1718, n_1749, n_1683, n_1916, n_2598, n_597, n_280, n_1270, n_2549, n_1187, n_610, n_1403, n_1669, n_1852, n_1024, n_1768, n_2153, n_2544, n_2381, n_198, n_1847, n_2052, n_179, n_248, n_2302, n_517, n_1667, n_667, n_1206, n_621, n_1037, n_1397, n_1279, n_1115, n_750, n_901, n_1499, n_468, n_2755, n_923, n_504, n_1409, n_1841, n_2637, n_2823, n_1639, n_1623, n_183, n_1015, n_1503, n_2819, n_466, n_2526, n_2423, n_1057, n_2548, n_603, n_991, n_2785, n_1657, n_235, n_1126, n_2412, n_1997, n_2636, n_340, n_710, n_1108, n_1818, n_2439, n_2404, n_1182, n_1298, n_2559, n_2177, n_39, n_2595, n_2088, n_73, n_1611, n_785, n_2740, n_746, n_609, n_1601, n_1960, n_2694, n_2061, n_1686, n_2757, n_2337, n_2401, n_101, n_167, n_1356, n_1589, n_127, n_2309, n_2900, n_2607, n_1740, n_2737, n_1497, n_2890, n_1168, n_1216, n_1943, n_133, n_1320, n_2716, n_96, n_2452, n_1430, n_1316, n_1287, n_2722, n_1452, n_2854, n_2499, n_1622, n_1586, n_2543, n_2264, n_302, n_1694, n_380, n_1535, n_2486, n_137, n_2571, n_1596, n_20, n_1190, n_1734, n_397, n_2902, n_1983, n_1938, n_2498, n_122, n_2220, n_2577, n_34, n_1262, n_2472, n_218, n_1891, n_2171, n_1213, n_70, n_2235, n_1350, n_1673, n_2232, n_1715, n_172, n_1443, n_1272, n_2392, n_2894, n_2790, n_239, n_2037, n_97, n_2808, n_2298, n_782, n_2326, n_1539, n_490, n_220, n_809, n_1043, n_1797, n_1608, n_986, n_2305, n_2120, n_80, n_1472, n_2050, n_2373, n_2164, n_2402, n_2225, n_1081, n_402, n_1870, n_352, n_1692, n_800, n_1084, n_1171, n_460, n_2169, n_2371, n_1827, n_1361, n_1864, n_2006, n_1491, n_2187, n_662, n_374, n_1152, n_1840, n_1705, n_450, n_2904, n_2244, n_2586, n_1684, n_921, n_2446, n_1346, n_711, n_1642, n_579, n_1352, n_2789, n_2872, n_937, n_2257, n_1682, n_2017, n_370, n_1695, n_1828, n_2046, n_2272, n_2699, n_2200, n_650, n_1046, n_2560, n_1940, n_1979, n_2760, n_2704, n_1145, n_330, n_1121, n_1102, n_1963, n_2738, n_972, n_1405, n_2376, n_258, n_1406, n_456, n_2766, n_1332, n_260, n_2670, n_313, n_2700, n_624, n_962, n_1041, n_2346, n_565, n_356, n_1569, n_936, n_1883, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_2342, n_2167, n_2084, n_2882, n_2541, n_654, n_411, n_2518, n_2458, n_152, n_1222, n_599, n_776, n_321, n_1823, n_2479, n_105, n_2782, n_227, n_1974, n_2673, n_2456, n_1720, n_2527, n_204, n_482, n_934, n_1637, n_2635, n_1407, n_1795, n_2768, n_2871, n_420, n_2688, n_1341, n_394, n_1456, n_1845, n_1489, n_164, n_2314, n_23, n_942, n_2798, n_2852, n_1524, n_543, n_2229, n_1964, n_2288, n_1920, n_2753, n_2099, n_1496, n_1271, n_1545, n_2007, n_2039, n_1946, n_1355, n_1225, n_1544, n_1485, n_2258, n_325, n_1640, n_804, n_464, n_1846, n_2406, n_533, n_2390, n_806, n_879, n_959, n_2310, n_2506, n_584, n_2141, n_2562, n_244, n_2642, n_1343, n_1522, n_76, n_2734, n_548, n_1782, n_94, n_282, n_2383, n_2626, n_1676, n_833, n_1830, n_2351, n_1567, n_523, n_1319, n_707, n_345, n_1900, n_799, n_1548, n_1155, n_2536, n_139, n_2196, n_41, n_2629, n_273, n_1633, n_2195, n_2809, n_787, n_2172, n_2835, n_1416, n_1528, n_2820, n_2293, n_1146, n_2021, n_2454, n_2114, n_159, n_1086, n_1066, n_1948, n_157, n_2125, n_2026, n_1282, n_2561, n_550, n_2567, n_2322, n_275, n_652, n_2154, n_2727, n_560, n_1906, n_1484, n_1241, n_1321, n_1672, n_569, n_2533, n_1758, n_2283, n_2869, n_2422, n_1925, n_737, n_1318, n_1914, n_1235, n_1229, n_2759, n_2361, n_306, n_1292, n_1373, n_21, n_2266, n_346, n_3, n_2427, n_1029, n_1447, n_2388, n_2056, n_790, n_2611, n_2901, n_138, n_1706, n_1498, n_2653, n_2417, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_2189, n_2680, n_2246, n_1047, n_1984, n_2236, n_1385, n_431, n_24, n_459, n_1269, n_1931, n_2083, n_2834, n_502, n_2668, n_672, n_2441, n_1257, n_1751, n_2840, n_285, n_1375, n_1941, n_85, n_2128, n_655, n_706, n_1045, n_1650, n_786, n_1794, n_1236, n_1962, n_1559, n_1725, n_1928, n_2398, n_1872, n_834, n_19, n_29, n_2695, n_75, n_743, n_766, n_430, n_1741, n_1325, n_1002, n_1746, n_1949, n_545, n_2671, n_489, n_2761, n_2885, n_2793, n_2715, n_2888, n_1804, n_1727, n_251, n_2508, n_1019, n_636, n_2054, n_729, n_110, n_151, n_876, n_774, n_2845, n_1337, n_660, n_2062, n_2041, n_438, n_1477, n_1360, n_2839, n_1860, n_2856, n_1904, n_2874, n_1200, n_2070, n_2588, n_479, n_1607, n_1353, n_1777, n_1908, n_1454, n_2484, n_2348, n_2614, n_2126, n_869, n_1154, n_1113, n_1600, n_2833, n_2253, n_2758, n_2366, n_646, n_528, n_391, n_1098, n_1329, n_2045, n_817, n_2261, n_2216, n_2210, n_262, n_187, n_897, n_846, n_2066, n_841, n_1476, n_2516, n_1001, n_508, n_1800, n_2241, n_1050, n_1411, n_1463, n_2903, n_2827, n_1177, n_332, n_1150, n_1742, n_1562, n_1690, n_398, n_1191, n_1826, n_566, n_1023, n_1882, n_1076, n_1118, n_194, n_57, n_1007, n_1807, n_1929, n_1378, n_2369, n_855, n_1592, n_1759, n_2719, n_1814, n_1631, n_52, n_591, n_1377, n_1879, n_256, n_853, n_440, n_695, n_1542, n_2587, n_875, n_209, n_367, n_680, n_1678, n_2569, n_661, n_2400, n_1716, n_278, n_1256, n_671, n_1953, n_7, n_933, n_740, n_703, n_978, n_2752, n_384, n_1976, n_2905, n_1291, n_1217, n_751, n_749, n_1824, n_310, n_1628, n_1324, n_1399, n_2122, n_2109, n_1435, n_969, n_988, n_2140, n_1065, n_2796, n_2507, n_84, n_1401, n_2358, n_1255, n_568, n_1516, n_143, n_1536, n_180, n_2163, n_2186, n_2029, n_2815, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_2528, n_2814, n_214, n_246, n_2787, n_1338, n_1097, n_2395, n_935, n_781, n_789, n_1554, n_1130, n_181, n_1810, n_182, n_573, n_769, n_2380, n_676, n_327, n_1120, n_832, n_1583, n_1730, n_2295, n_555, n_389, n_814, n_2746, n_1643, n_2020, n_2500, n_2269, n_1729, n_669, n_2290, n_2048, n_176, n_114, n_300, n_222, n_2005, n_747, n_74, n_2565, n_1389, n_1105, n_721, n_1461, n_742, n_535, n_691, n_372, n_2076, n_2736, n_111, n_2883, n_314, n_1408, n_378, n_1196, n_377, n_1598, n_863, n_2175, n_601, n_2182, n_338, n_2910, n_1283, n_2385, n_918, n_748, n_506, n_1114, n_1785, n_56, n_763, n_1147, n_1848, n_360, n_1754, n_2149, n_2396, n_1506, n_119, n_2584, n_1652, n_1812, n_957, n_1994, n_895, n_866, n_1227, n_2450, n_2485, n_2284, n_191, n_2566, n_387, n_2287, n_452, n_744, n_971, n_2702, n_946, n_344, n_2906, n_761, n_1303, n_2769, n_1205, n_2492, n_1258, n_2438, n_2914, n_1392, n_174, n_1173, n_1924, n_525, n_2463, n_2881, n_1677, n_1116, n_611, n_1570, n_1702, n_1219, n_1780, n_1689, n_8, n_2180, n_2858, n_2679, n_1174, n_1944, n_1016, n_1347, n_795, n_1501, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_2117, n_2234, n_2779, n_2685, n_1083, n_109, n_445, n_1561, n_2741, n_930, n_888, n_2275, n_1112, n_2465, n_2620, n_2081, n_2168, n_2568, n_234, n_2022, n_1945, n_2203, n_910, n_1656, n_1721, n_1460, n_911, n_2112, n_2255, n_82, n_1464, n_27, n_236, n_653, n_1737, n_2430, n_1414, n_752, n_908, n_2649, n_2721, n_944, n_2034, n_576, n_1028, n_2106, n_472, n_2862, n_270, n_2265, n_2615, n_414, n_2683, n_1922, n_563, n_2032, n_2744, n_1011, n_2474, n_1566, n_1215, n_2437, n_25, n_93, n_839, n_2444, n_2743, n_708, n_1973, n_2267, n_668, n_626, n_990, n_1500, n_779, n_1537, n_1821, n_2205, n_1104, n_854, n_1058, n_2312, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_2242, n_1509, n_103, n_1693, n_1109, n_185, n_2222, n_712, n_348, n_1276, n_376, n_2015, n_2118, n_2111, n_2466, n_390, n_2915, n_2530, n_1148, n_31, n_2188, n_2505, n_334, n_1989, n_1161, n_2609, n_1085, n_232, n_2802, n_2014, n_2042, n_46, n_1239, n_771, n_1584, n_2425, n_470, n_475, n_924, n_298, n_1582, n_492, n_2318, n_2408, n_1149, n_265, n_1184, n_2483, n_228, n_719, n_1972, n_2592, n_1525, n_2594, n_455, n_2666, n_1585, n_1851, n_363, n_1799, n_1090, n_2147, n_2564, n_592, n_1816, n_2503, n_2433, n_1518, n_829, n_1156, n_1362, n_393, n_984, n_2600, n_1829, n_503, n_2035, n_1450, n_1638, n_132, n_868, n_570, n_859, n_2033, n_406, n_735, n_1789, n_2531, n_1770, n_878, n_620, n_130, n_519, n_2523, n_307, n_469, n_1218, n_2413, n_500, n_1482, n_981, n_714, n_1349, n_291, n_1144, n_2071, n_357, n_2429, n_985, n_2233, n_2440, n_2723, n_481, n_997, n_1710, n_2800, n_2161, n_1301, n_2805, n_802, n_561, n_33, n_980, n_2681, n_1306, n_2010, n_2282, n_1651, n_1198, n_2360, n_2047, n_2651, n_2095, n_1609, n_2174, n_2799, n_436, n_116, n_2334, n_409, n_1244, n_1685, n_1763, n_1998, n_1574, n_2426, n_2490, n_2844, n_240, n_756, n_2303, n_1619, n_2478, n_1981, n_2285, n_1606, n_810, n_1133, n_635, n_95, n_1194, n_2742, n_2640, n_1051, n_253, n_1552, n_2918, n_583, n_1996, n_2367, n_249, n_201, n_2867, n_1039, n_1442, n_2726, n_1034, n_2043, n_1480, n_1158, n_2909, n_2248, n_754, n_941, n_975, n_1031, n_115, n_1305, n_2363, n_2578, n_553, n_43, n_849, n_2662, n_753, n_1753, n_2795, n_2471, n_467, n_2540, n_269, n_359, n_973, n_2807, n_1921, n_1479, n_1055, n_1675, n_2197, n_2217, n_582, n_2065, n_2879, n_861, n_857, n_967, n_571, n_2215, n_2461, n_271, n_404, n_2001, n_158, n_2107, n_1884, n_206, n_2040, n_679, n_633, n_1170, n_665, n_1629, n_2221, n_588, n_225, n_1260, n_308, n_309, n_1819, n_2055, n_1010, n_2553, n_149, n_1040, n_915, n_632, n_1166, n_2038, n_812, n_2891, n_1131, n_2634, n_1761, n_2709, n_534, n_1578, n_1006, n_1861, n_373, n_87, n_1632, n_1890, n_1805, n_2477, n_257, n_1557, n_1888, n_2280, n_1833, n_730, n_1311, n_1494, n_2325, n_670, n_203, n_1850, n_1898, n_2443, n_2697, n_2308, n_2162, n_1868, n_207, n_2333, n_2079, n_1089, n_1887, n_1587, n_2512, n_1365, n_1417, n_205, n_1242, n_2086, n_2185, n_1836, n_2774, n_681, n_1226, n_1274, n_1486, n_2166, n_412, n_2899, n_640, n_1322, n_81, n_965, n_1899, n_1428, n_1616, n_1576, n_1856, n_1862, n_1958, n_2077, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_2632, n_422, n_2579, n_722, n_862, n_2105, n_135, n_165, n_2098, n_540, n_1423, n_2813, n_1935, n_2027, n_457, n_2223, n_2091, n_364, n_1915, n_629, n_1621, n_1748, n_2547, n_2415, n_900, n_1449, n_531, n_827, n_2912, n_60, n_361, n_2659, n_1025, n_2419, n_2116, n_336, n_2320, n_12, n_1885, n_2677, n_1013, n_1259, n_192, n_2183, n_1538, n_51, n_649, n_1612, n_1240, n_13275);

input n_992;
input n_2542;
input n_1671;
input n_1;
input n_2817;
input n_801;
input n_1613;
input n_1234;
input n_1458;
input n_2576;
input n_1199;
input n_1674;
input n_741;
input n_1027;
input n_1351;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_2157;
input n_2332;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_2003;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_2353;
input n_2534;
input n_1357;
input n_1853;
input n_77;
input n_783;
input n_2451;
input n_1738;
input n_2243;
input n_798;
input n_188;
input n_1575;
input n_1854;
input n_2324;
input n_1923;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_2260;
input n_677;
input n_1708;
input n_805;
input n_1151;
input n_396;
input n_1739;
input n_350;
input n_78;
input n_2051;
input n_2317;
input n_1380;
input n_2359;
input n_442;
input n_480;
input n_142;
input n_2847;
input n_1402;
input n_2557;
input n_1688;
input n_1691;
input n_1975;
input n_1009;
input n_1743;
input n_62;
input n_1930;
input n_2405;
input n_1160;
input n_883;
input n_2647;
input n_1238;
input n_1991;
input n_2570;
input n_2179;
input n_2386;
input n_1724;
input n_1032;
input n_2336;
input n_1247;
input n_1547;
input n_2521;
input n_1553;
input n_893;
input n_1099;
input n_2491;
input n_1264;
input n_1192;
input n_471;
input n_1844;
input n_424;
input n_1700;
input n_1555;
input n_1415;
input n_2211;
input n_1370;
input n_1786;
input n_369;
input n_287;
input n_2382;
input n_2672;
input n_2291;
input n_415;
input n_830;
input n_2299;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_2886;
input n_200;
input n_1985;
input n_447;
input n_2838;
input n_2184;
input n_1803;
input n_1172;
input n_852;
input n_2509;
input n_71;
input n_229;
input n_2513;
input n_1590;
input n_2645;
input n_1532;
input n_2313;
input n_2628;
input n_1393;
input n_1517;
input n_1867;
input n_1704;
input n_1078;
input n_250;
input n_544;
input n_1711;
input n_2247;
input n_1140;
input n_2630;
input n_1444;
input n_1670;
input n_1603;
input n_2344;
input n_1579;
input n_35;
input n_2365;
input n_2470;
input n_2321;
input n_1263;
input n_2019;
input n_836;
input n_375;
input n_2074;
input n_2447;
input n_522;
input n_2919;
input n_2129;
input n_2340;
input n_1261;
input n_945;
input n_2286;
input n_1649;
input n_2018;
input n_2094;
input n_1903;
input n_1511;
input n_1143;
input n_2356;
input n_2399;
input n_1422;
input n_1232;
input n_1772;
input n_1572;
input n_616;
input n_658;
input n_1874;
input n_1119;
input n_2865;
input n_2825;
input n_2013;
input n_428;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2044;
input n_1954;
input n_1735;
input n_2510;
input n_1541;
input n_1300;
input n_641;
input n_2480;
input n_2739;
input n_822;
input n_693;
input n_1313;
input n_2791;
input n_1056;
input n_2212;
input n_758;
input n_516;
input n_1455;
input n_2418;
input n_2864;
input n_1163;
input n_2729;
input n_1180;
input n_2256;
input n_2582;
input n_943;
input n_1798;
input n_1550;
input n_2703;
input n_491;
input n_2786;
input n_1591;
input n_42;
input n_772;
input n_2806;
input n_1344;
input n_2730;
input n_2495;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_1781;
input n_1971;
input n_2058;
input n_2090;
input n_2603;
input n_405;
input n_213;
input n_2660;
input n_538;
input n_2173;
input n_2004;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_1345;
input n_1820;
input n_2873;
input n_494;
input n_539;
input n_493;
input n_155;
input n_2880;
input n_2394;
input n_2108;
input n_45;
input n_454;
input n_1421;
input n_2836;
input n_1936;
input n_638;
input n_1404;
input n_1211;
input n_2124;
input n_381;
input n_2378;
input n_887;
input n_1660;
input n_1961;
input n_112;
input n_1280;
input n_713;
input n_2655;
input n_1400;
input n_2625;
input n_2843;
input n_126;
input n_1467;
input n_58;
input n_976;
input n_2155;
input n_224;
input n_2686;
input n_48;
input n_1445;
input n_2364;
input n_2551;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_1894;
input n_196;
input n_1231;
input n_2599;
input n_1978;
input n_2085;
input n_917;
input n_574;
input n_9;
input n_2370;
input n_2612;
input n_907;
input n_6;
input n_1446;
input n_14;
input n_2591;
input n_659;
input n_1815;
input n_2214;
input n_407;
input n_913;
input n_1658;
input n_2593;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1967;
input n_1054;
input n_559;
input n_2613;
input n_1333;
input n_2496;
input n_44;
input n_2708;
input n_1648;
input n_1911;
input n_1956;
input n_163;
input n_1644;
input n_2011;
input n_2725;
input n_2277;
input n_1558;
input n_1732;
input n_281;
input n_551;
input n_699;
input n_1986;
input n_2300;
input n_564;
input n_2397;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_1641;
input n_2113;
input n_1918;
input n_2190;
input n_2907;
input n_577;
input n_166;
input n_2735;
input n_1843;
input n_619;
input n_2268;
input n_1367;
input n_1336;
input n_521;
input n_2778;
input n_2850;
input n_572;
input n_395;
input n_813;
input n_1909;
input n_2080;
input n_1481;
input n_323;
input n_606;
input n_1441;
input n_818;
input n_1123;
input n_1309;
input n_92;
input n_2104;
input n_513;
input n_645;
input n_1381;
input n_331;
input n_1699;
input n_916;
input n_2093;
input n_2633;
input n_483;
input n_102;
input n_2207;
input n_1970;
input n_2770;
input n_608;
input n_261;
input n_2101;
input n_2696;
input n_630;
input n_2059;
input n_32;
input n_2198;
input n_541;
input n_512;
input n_2669;
input n_2073;
input n_2273;
input n_121;
input n_433;
input n_2546;
input n_792;
input n_2522;
input n_476;
input n_2792;
input n_2;
input n_1328;
input n_1957;
input n_2917;
input n_219;
input n_2616;
input n_1907;
input n_2529;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_1530;
input n_788;
input n_939;
input n_1543;
input n_821;
input n_2811;
input n_938;
input n_1302;
input n_1068;
input n_1599;
input n_329;
input n_982;
input n_2674;
input n_2832;
input n_549;
input n_1762;
input n_1910;
input n_1075;
input n_408;
input n_932;
input n_2831;
input n_61;
input n_237;
input n_1876;
input n_1895;
input n_2123;
input n_1697;
input n_2143;
input n_243;
input n_979;
input n_1873;
input n_905;
input n_1866;
input n_1680;
input n_117;
input n_175;
input n_322;
input n_993;
input n_2692;
input n_689;
input n_2031;
input n_354;
input n_2130;
input n_1330;
input n_1413;
input n_1605;
input n_2228;
input n_134;
input n_1988;
input n_1278;
input n_547;
input n_2455;
input n_2876;
input n_558;
input n_2654;
input n_2469;
input n_1064;
input n_1396;
input n_634;
input n_2355;
input n_136;
input n_966;
input n_2908;
input n_764;
input n_2751;
input n_2764;
input n_1663;
input n_2895;
input n_2009;
input n_692;
input n_733;
input n_1793;
input n_1233;
input n_1289;
input n_2714;
input n_2245;
input n_487;
input n_241;
input n_30;
input n_2068;
input n_1107;
input n_2866;
input n_2457;
input n_1014;
input n_1290;
input n_1703;
input n_2580;
input n_882;
input n_2176;
input n_2072;
input n_1354;
input n_2821;
input n_586;
input n_423;
input n_1865;
input n_1875;
input n_1701;
input n_2459;
input n_318;
input n_1111;
input n_1713;
input n_715;
input n_2678;
input n_1251;
input n_1265;
input n_2711;
input n_88;
input n_1726;
input n_1950;
input n_530;
input n_1563;
input n_1912;
input n_277;
input n_2434;
input n_1982;
input n_2878;
input n_618;
input n_1297;
input n_1662;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_2818;
input n_2428;
input n_674;
input n_871;
input n_922;
input n_268;
input n_1335;
input n_1760;
input n_1927;
input n_210;
input n_2028;
input n_1069;
input n_2664;
input n_5;
input n_1664;
input n_1722;
input n_612;
input n_2641;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_2008;
input n_2749;
input n_2192;
input n_2254;
input n_2345;
input n_1926;
input n_1175;
input n_328;
input n_1386;
input n_2311;
input n_1896;
input n_429;
input n_1747;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_2624;
input n_903;
input n_1540;
input n_1977;
input n_1802;
input n_1504;
input n_2350;
input n_2804;
input n_2453;
input n_286;
input n_254;
input n_2193;
input n_2676;
input n_1655;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_1801;
input n_1886;
input n_2092;
input n_2347;
input n_1654;
input n_816;
input n_1157;
input n_1750;
input n_1462;
input n_1188;
input n_1752;
input n_877;
input n_1813;
input n_2514;
input n_2206;
input n_604;
input n_2810;
input n_2319;
input n_2519;
input n_825;
input n_728;
input n_2916;
input n_1063;
input n_1588;
input n_2467;
input n_26;
input n_2602;
input n_2468;
input n_55;
input n_267;
input n_1124;
input n_1624;
input n_515;
input n_2096;
input n_1965;
input n_2476;
input n_598;
input n_696;
input n_1515;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_2733;
input n_2824;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_2377;
input n_295;
input n_701;
input n_2178;
input n_950;
input n_388;
input n_190;
input n_2812;
input n_484;
input n_2644;
input n_2036;
input n_2152;
input n_1709;
input n_2652;
input n_2411;
input n_2525;
input n_1825;
input n_2393;
input n_1757;
input n_1796;
input n_170;
input n_2657;
input n_1792;
input n_891;
input n_2067;
input n_2136;
input n_2409;
input n_2082;
input n_2252;
input n_1412;
input n_2497;
input n_2687;
input n_949;
input n_1630;
input n_678;
input n_2887;
input n_283;
input n_2075;
input n_2194;
input n_2619;
input n_91;
input n_2763;
input n_2762;
input n_1987;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_2271;
input n_1008;
input n_760;
input n_1546;
input n_2583;
input n_590;
input n_63;
input n_2606;
input n_362;
input n_148;
input n_2279;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_2794;
input n_1296;
input n_2663;
input n_1990;
input n_2391;
input n_304;
input n_2431;
input n_694;
input n_2150;
input n_1294;
input n_1420;
input n_125;
input n_1634;
input n_2078;
input n_297;
input n_595;
input n_627;
input n_1767;
input n_1779;
input n_524;
input n_1465;
input n_342;
input n_2622;
input n_1858;
input n_1044;
input n_2658;
input n_2665;
input n_2165;
input n_2133;
input n_1712;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_2558;
input n_2750;
input n_2775;
input n_1208;
input n_2893;
input n_1164;
input n_1295;
input n_1627;
input n_2728;
input n_2349;
input n_2684;
input n_2712;
input n_1072;
input n_1527;
input n_1495;
input n_1438;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_1487;
input n_2691;
input n_840;
input n_2913;
input n_874;
input n_1756;
input n_1128;
input n_2493;
input n_382;
input n_673;
input n_2230;
input n_2705;
input n_1969;
input n_2690;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_2145;
input n_1968;
input n_898;
input n_255;
input n_284;
input n_1952;
input n_865;
input n_2573;
input n_2646;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_1026;
input n_1880;
input n_2535;
input n_2631;
input n_38;
input n_289;
input n_1364;
input n_2436;
input n_615;
input n_2870;
input n_1249;
input n_2706;
input n_59;
input n_1293;
input n_2693;
input n_1127;
input n_1512;
input n_2151;
input n_1451;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_2767;
input n_727;
input n_894;
input n_1839;
input n_2341;
input n_685;
input n_1765;
input n_353;
input n_2707;
input n_605;
input n_1514;
input n_1863;
input n_826;
input n_1646;
input n_872;
input n_1139;
input n_1714;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_1521;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_2537;
input n_2897;
input n_305;
input n_72;
input n_2554;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_2089;
input n_1376;
input n_1513;
input n_2747;
input n_413;
input n_791;
input n_1913;
input n_510;
input n_837;
input n_2097;
input n_79;
input n_2170;
input n_1488;
input n_2853;
input n_1808;
input n_948;
input n_2517;
input n_2713;
input n_704;
input n_2148;
input n_977;
input n_2339;
input n_1005;
input n_1947;
input n_2765;
input n_2861;
input n_536;
input n_1788;
input n_1999;
input n_2731;
input n_622;
input n_147;
input n_2590;
input n_2643;
input n_1469;
input n_2060;
input n_2608;
input n_1838;
input n_2638;
input n_1835;
input n_1766;
input n_1776;
input n_1959;
input n_2002;
input n_581;
input n_2650;
input n_2138;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_2414;
input n_1340;
input n_1771;
input n_2316;
input n_631;
input n_720;
input n_153;
input n_842;
input n_2262;
input n_1707;
input n_2239;
input n_1432;
input n_156;
input n_145;
input n_2208;
input n_843;
input n_656;
input n_989;
input n_2604;
input n_2407;
input n_1277;
input n_2816;
input n_797;
input n_2689;
input n_1473;
input n_2191;
input n_1723;
input n_2717;
input n_1246;
input n_1878;
input n_2574;
input n_899;
input n_189;
input n_738;
input n_2012;
input n_1304;
input n_1035;
input n_294;
input n_2842;
input n_499;
input n_2675;
input n_1426;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_2134;
input n_1529;
input n_2335;
input n_2473;
input n_1022;
input n_614;
input n_529;
input n_2069;
input n_2307;
input n_2362;
input n_425;
input n_684;
input n_2539;
input n_2667;
input n_2698;
input n_1431;
input n_1615;
input n_1474;
input n_1571;
input n_1809;
input n_1577;
input n_2297;
input n_1181;
input n_2119;
input n_1822;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_2489;
input n_1087;
input n_1448;
input n_1992;
input n_648;
input n_657;
input n_1049;
input n_2771;
input n_2445;
input n_2057;
input n_2103;
input n_2605;
input n_1666;
input n_2772;
input n_1505;
input n_803;
input n_290;
input n_118;
input n_1717;
input n_926;
input n_1817;
input n_2449;
input n_927;
input n_2610;
input n_1849;
input n_2848;
input n_919;
input n_2868;
input n_1698;
input n_478;
input n_2231;
input n_929;
input n_107;
input n_2520;
input n_1228;
input n_417;
input n_2857;
input n_446;
input n_89;
input n_1568;
input n_1490;
input n_2372;
input n_777;
input n_1299;
input n_272;
input n_2896;
input n_526;
input n_2718;
input n_2639;
input n_1183;
input n_1436;
input n_2898;
input n_2251;
input n_1384;
input n_69;
input n_2494;
input n_2501;
input n_2238;
input n_293;
input n_2368;
input n_53;
input n_458;
input n_1070;
input n_2403;
input n_2837;
input n_998;
input n_16;
input n_717;
input n_1665;
input n_18;
input n_2524;
input n_154;
input n_1383;
input n_2460;
input n_1178;
input n_98;
input n_2127;
input n_1424;
input n_2338;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_2137;
input n_1626;
input n_1507;
input n_2482;
input n_184;
input n_552;
input n_2532;
input n_1358;
input n_1811;
input n_1388;
input n_216;
input n_2481;
input n_912;
input n_1857;
input n_1519;
input n_2144;
input n_745;
input n_1284;
input n_1604;
input n_2296;
input n_2424;
input n_1142;
input n_2849;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1774;
input n_2354;
input n_2682;
input n_2589;
input n_1395;
input n_2110;
input n_2199;
input n_2661;
input n_731;
input n_2877;
input n_1502;
input n_1659;
input n_1955;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_2442;
input n_312;
input n_1791;
input n_1368;
input n_66;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_1897;
input n_2064;
input n_880;
input n_2053;
input n_2259;
input n_2121;
input n_2773;
input n_2545;
input n_889;
input n_2432;
input n_2710;
input n_150;
input n_1478;
input n_589;
input n_1310;
input n_819;
input n_2294;
input n_1363;
input n_2581;
input n_1334;
input n_1942;
input n_1966;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_1837;
input n_2218;
input n_2788;
input n_477;
input n_2435;
input n_954;
input n_864;
input n_2504;
input n_2797;
input n_2623;
input n_1110;
input n_2213;
input n_1410;
input n_399;
input n_2389;
input n_1440;
input n_124;
input n_2132;
input n_2892;
input n_2063;
input n_1382;
input n_1534;
input n_1564;
input n_1736;
input n_211;
input n_2748;
input n_1483;
input n_1834;
input n_2331;
input n_1372;
input n_231;
input n_2292;
input n_2860;
input n_2330;
input n_40;
input n_1457;
input n_505;
input n_1719;
input n_319;
input n_1339;
input n_1787;
input n_2701;
input n_2475;
input n_537;
input n_2511;
input n_1993;
input n_2281;
input n_1427;
input n_311;
input n_2416;
input n_2745;
input n_2617;
input n_2776;
input n_1466;
input n_10;
input n_403;
input n_1919;
input n_1080;
input n_723;
input n_1877;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1939;
input n_2030;
input n_1769;
input n_1220;
input n_2323;
input n_1893;
input n_556;
input n_2784;
input n_2209;
input n_2301;
input n_162;
input n_2387;
input n_1755;
input n_1602;
input n_2421;
input n_1136;
input n_2618;
input n_2025;
input n_2357;
input n_2846;
input n_2464;
input n_128;
input n_1125;
input n_970;
input n_2488;
input n_2224;
input n_1980;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_2329;
input n_1092;
input n_2237;
input n_441;
input n_221;
input n_1060;
input n_1951;
input n_2250;
input n_444;
input n_146;
input n_1252;
input n_1784;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1773;
input n_1775;
input n_2115;
input n_2410;
input n_2552;
input n_1053;
input n_2374;
input n_416;
input n_1681;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1783;
input n_1533;
input n_1597;
input n_2780;
input n_4;
input n_266;
input n_296;
input n_2596;
input n_2274;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_1618;
input n_217;
input n_518;
input n_1531;
input n_2828;
input n_1185;
input n_453;
input n_215;
input n_2384;
input n_1745;
input n_914;
input n_759;
input n_2724;
input n_1831;
input n_426;
input n_317;
input n_2585;
input n_2621;
input n_1653;
input n_2352;
input n_1679;
input n_1625;
input n_90;
input n_2601;
input n_2160;
input n_54;
input n_1453;
input n_2146;
input n_2226;
input n_2131;
input n_488;
input n_2502;
input n_2801;
input n_497;
input n_2920;
input n_773;
input n_1901;
input n_920;
input n_99;
input n_1374;
input n_2556;
input n_2648;
input n_1315;
input n_1647;
input n_13;
input n_2575;
input n_2754;
input n_1224;
input n_2783;
input n_2306;
input n_1614;
input n_1459;
input n_1892;
input n_1933;
input n_2462;
input n_1135;
input n_1169;
input n_1179;
input n_2889;
input n_401;
input n_324;
input n_1617;
input n_335;
input n_1470;
input n_2550;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_2732;
input n_301;
input n_274;
input n_1096;
input n_2249;
input n_1091;
input n_1917;
input n_2000;
input n_1580;
input n_2227;
input n_2270;
input n_2822;
input n_1425;
input n_36;
input n_1881;
input n_1267;
input n_1281;
input n_1806;
input n_983;
input n_2023;
input n_427;
input n_2572;
input n_2204;
input n_1520;
input n_496;
input n_2720;
input n_2159;
input n_906;
input n_1390;
input n_688;
input n_2289;
input n_1077;
input n_1733;
input n_2315;
input n_1419;
input n_2863;
input n_351;
input n_259;
input n_1731;
input n_177;
input n_2158;
input n_2087;
input n_1855;
input n_1636;
input n_1437;
input n_2135;
input n_1645;
input n_1832;
input n_385;
input n_1687;
input n_1439;
input n_2328;
input n_1323;
input n_2859;
input n_2202;
input n_858;
input n_2049;
input n_1331;
input n_613;
input n_736;
input n_2627;
input n_501;
input n_956;
input n_960;
input n_2276;
input n_663;
input n_856;
input n_2803;
input n_2100;
input n_379;
input n_778;
input n_1668;
input n_2777;
input n_1134;
input n_2830;
input n_2781;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_1696;
input n_2829;
input n_1995;
input n_1594;
input n_2181;
input n_664;
input n_1869;
input n_171;
input n_2911;
input n_1764;
input n_169;
input n_1429;
input n_2826;
input n_1610;
input n_1889;
input n_2379;
input n_435;
input n_1905;
input n_2016;
input n_2343;
input n_793;
input n_326;
input n_587;
input n_1593;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_1937;
input n_465;
input n_1790;
input n_1778;
input n_1635;
input n_1079;
input n_341;
input n_2515;
input n_1744;
input n_828;
input n_2139;
input n_2142;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_2448;
input n_1103;
input n_2875;
input n_2555;
input n_144;
input n_2219;
input n_1203;
input n_2851;
input n_820;
input n_2327;
input n_951;
input n_106;
input n_2201;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_2841;
input n_2420;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_2263;
input n_2304;
input n_1508;
input n_2487;
input n_732;
input n_974;
input n_2240;
input n_392;
input n_2278;
input n_2656;
input n_2538;
input n_724;
input n_2597;
input n_2375;
input n_1934;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_1728;
input n_557;
input n_2756;
input n_1871;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1661;
input n_1275;
input n_2884;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_421;
input n_1468;
input n_2855;
input n_1859;
input n_2102;
input n_2563;
input n_238;
input n_1095;
input n_2024;
input n_1595;
input n_202;
input n_2156;
input n_1718;
input n_1749;
input n_1683;
input n_1916;
input n_2598;
input n_597;
input n_280;
input n_1270;
input n_2549;
input n_1187;
input n_610;
input n_1403;
input n_1669;
input n_1852;
input n_1024;
input n_1768;
input n_2153;
input n_2544;
input n_2381;
input n_198;
input n_1847;
input n_2052;
input n_179;
input n_248;
input n_2302;
input n_517;
input n_1667;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1397;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_468;
input n_2755;
input n_923;
input n_504;
input n_1409;
input n_1841;
input n_2637;
input n_2823;
input n_1639;
input n_1623;
input n_183;
input n_1015;
input n_1503;
input n_2819;
input n_466;
input n_2526;
input n_2423;
input n_1057;
input n_2548;
input n_603;
input n_991;
input n_2785;
input n_1657;
input n_235;
input n_1126;
input n_2412;
input n_1997;
input n_2636;
input n_340;
input n_710;
input n_1108;
input n_1818;
input n_2439;
input n_2404;
input n_1182;
input n_1298;
input n_2559;
input n_2177;
input n_39;
input n_2595;
input n_2088;
input n_73;
input n_1611;
input n_785;
input n_2740;
input n_746;
input n_609;
input n_1601;
input n_1960;
input n_2694;
input n_2061;
input n_1686;
input n_2757;
input n_2337;
input n_2401;
input n_101;
input n_167;
input n_1356;
input n_1589;
input n_127;
input n_2309;
input n_2900;
input n_2607;
input n_1740;
input n_2737;
input n_1497;
input n_2890;
input n_1168;
input n_1216;
input n_1943;
input n_133;
input n_1320;
input n_2716;
input n_96;
input n_2452;
input n_1430;
input n_1316;
input n_1287;
input n_2722;
input n_1452;
input n_2854;
input n_2499;
input n_1622;
input n_1586;
input n_2543;
input n_2264;
input n_302;
input n_1694;
input n_380;
input n_1535;
input n_2486;
input n_137;
input n_2571;
input n_1596;
input n_20;
input n_1190;
input n_1734;
input n_397;
input n_2902;
input n_1983;
input n_1938;
input n_2498;
input n_122;
input n_2220;
input n_2577;
input n_34;
input n_1262;
input n_2472;
input n_218;
input n_1891;
input n_2171;
input n_1213;
input n_70;
input n_2235;
input n_1350;
input n_1673;
input n_2232;
input n_1715;
input n_172;
input n_1443;
input n_1272;
input n_2392;
input n_2894;
input n_2790;
input n_239;
input n_2037;
input n_97;
input n_2808;
input n_2298;
input n_782;
input n_2326;
input n_1539;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_1797;
input n_1608;
input n_986;
input n_2305;
input n_2120;
input n_80;
input n_1472;
input n_2050;
input n_2373;
input n_2164;
input n_2402;
input n_2225;
input n_1081;
input n_402;
input n_1870;
input n_352;
input n_1692;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_2169;
input n_2371;
input n_1827;
input n_1361;
input n_1864;
input n_2006;
input n_1491;
input n_2187;
input n_662;
input n_374;
input n_1152;
input n_1840;
input n_1705;
input n_450;
input n_2904;
input n_2244;
input n_2586;
input n_1684;
input n_921;
input n_2446;
input n_1346;
input n_711;
input n_1642;
input n_579;
input n_1352;
input n_2789;
input n_2872;
input n_937;
input n_2257;
input n_1682;
input n_2017;
input n_370;
input n_1695;
input n_1828;
input n_2046;
input n_2272;
input n_2699;
input n_2200;
input n_650;
input n_1046;
input n_2560;
input n_1940;
input n_1979;
input n_2760;
input n_2704;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_1963;
input n_2738;
input n_972;
input n_1405;
input n_2376;
input n_258;
input n_1406;
input n_456;
input n_2766;
input n_1332;
input n_260;
input n_2670;
input n_313;
input n_2700;
input n_624;
input n_962;
input n_1041;
input n_2346;
input n_565;
input n_356;
input n_1569;
input n_936;
input n_1883;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_2342;
input n_2167;
input n_2084;
input n_2882;
input n_2541;
input n_654;
input n_411;
input n_2518;
input n_2458;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_1823;
input n_2479;
input n_105;
input n_2782;
input n_227;
input n_1974;
input n_2673;
input n_2456;
input n_1720;
input n_2527;
input n_204;
input n_482;
input n_934;
input n_1637;
input n_2635;
input n_1407;
input n_1795;
input n_2768;
input n_2871;
input n_420;
input n_2688;
input n_1341;
input n_394;
input n_1456;
input n_1845;
input n_1489;
input n_164;
input n_2314;
input n_23;
input n_942;
input n_2798;
input n_2852;
input n_1524;
input n_543;
input n_2229;
input n_1964;
input n_2288;
input n_1920;
input n_2753;
input n_2099;
input n_1496;
input n_1271;
input n_1545;
input n_2007;
input n_2039;
input n_1946;
input n_1355;
input n_1225;
input n_1544;
input n_1485;
input n_2258;
input n_325;
input n_1640;
input n_804;
input n_464;
input n_1846;
input n_2406;
input n_533;
input n_2390;
input n_806;
input n_879;
input n_959;
input n_2310;
input n_2506;
input n_584;
input n_2141;
input n_2562;
input n_244;
input n_2642;
input n_1343;
input n_1522;
input n_76;
input n_2734;
input n_548;
input n_1782;
input n_94;
input n_282;
input n_2383;
input n_2626;
input n_1676;
input n_833;
input n_1830;
input n_2351;
input n_1567;
input n_523;
input n_1319;
input n_707;
input n_345;
input n_1900;
input n_799;
input n_1548;
input n_1155;
input n_2536;
input n_139;
input n_2196;
input n_41;
input n_2629;
input n_273;
input n_1633;
input n_2195;
input n_2809;
input n_787;
input n_2172;
input n_2835;
input n_1416;
input n_1528;
input n_2820;
input n_2293;
input n_1146;
input n_2021;
input n_2454;
input n_2114;
input n_159;
input n_1086;
input n_1066;
input n_1948;
input n_157;
input n_2125;
input n_2026;
input n_1282;
input n_2561;
input n_550;
input n_2567;
input n_2322;
input n_275;
input n_652;
input n_2154;
input n_2727;
input n_560;
input n_1906;
input n_1484;
input n_1241;
input n_1321;
input n_1672;
input n_569;
input n_2533;
input n_1758;
input n_2283;
input n_2869;
input n_2422;
input n_1925;
input n_737;
input n_1318;
input n_1914;
input n_1235;
input n_1229;
input n_2759;
input n_2361;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_2266;
input n_346;
input n_3;
input n_2427;
input n_1029;
input n_1447;
input n_2388;
input n_2056;
input n_790;
input n_2611;
input n_2901;
input n_138;
input n_1706;
input n_1498;
input n_2653;
input n_2417;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_2189;
input n_2680;
input n_2246;
input n_1047;
input n_1984;
input n_2236;
input n_1385;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_1931;
input n_2083;
input n_2834;
input n_502;
input n_2668;
input n_672;
input n_2441;
input n_1257;
input n_1751;
input n_2840;
input n_285;
input n_1375;
input n_1941;
input n_85;
input n_2128;
input n_655;
input n_706;
input n_1045;
input n_1650;
input n_786;
input n_1794;
input n_1236;
input n_1962;
input n_1559;
input n_1725;
input n_1928;
input n_2398;
input n_1872;
input n_834;
input n_19;
input n_29;
input n_2695;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1741;
input n_1325;
input n_1002;
input n_1746;
input n_1949;
input n_545;
input n_2671;
input n_489;
input n_2761;
input n_2885;
input n_2793;
input n_2715;
input n_2888;
input n_1804;
input n_1727;
input n_251;
input n_2508;
input n_1019;
input n_636;
input n_2054;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_2845;
input n_1337;
input n_660;
input n_2062;
input n_2041;
input n_438;
input n_1477;
input n_1360;
input n_2839;
input n_1860;
input n_2856;
input n_1904;
input n_2874;
input n_1200;
input n_2070;
input n_2588;
input n_479;
input n_1607;
input n_1353;
input n_1777;
input n_1908;
input n_1454;
input n_2484;
input n_2348;
input n_2614;
input n_2126;
input n_869;
input n_1154;
input n_1113;
input n_1600;
input n_2833;
input n_2253;
input n_2758;
input n_2366;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_1329;
input n_2045;
input n_817;
input n_2261;
input n_2216;
input n_2210;
input n_262;
input n_187;
input n_897;
input n_846;
input n_2066;
input n_841;
input n_1476;
input n_2516;
input n_1001;
input n_508;
input n_1800;
input n_2241;
input n_1050;
input n_1411;
input n_1463;
input n_2903;
input n_2827;
input n_1177;
input n_332;
input n_1150;
input n_1742;
input n_1562;
input n_1690;
input n_398;
input n_1191;
input n_1826;
input n_566;
input n_1023;
input n_1882;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_1807;
input n_1929;
input n_1378;
input n_2369;
input n_855;
input n_1592;
input n_1759;
input n_2719;
input n_1814;
input n_1631;
input n_52;
input n_591;
input n_1377;
input n_1879;
input n_256;
input n_853;
input n_440;
input n_695;
input n_1542;
input n_2587;
input n_875;
input n_209;
input n_367;
input n_680;
input n_1678;
input n_2569;
input n_661;
input n_2400;
input n_1716;
input n_278;
input n_1256;
input n_671;
input n_1953;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_2752;
input n_384;
input n_1976;
input n_2905;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_1824;
input n_310;
input n_1628;
input n_1324;
input n_1399;
input n_2122;
input n_2109;
input n_1435;
input n_969;
input n_988;
input n_2140;
input n_1065;
input n_2796;
input n_2507;
input n_84;
input n_1401;
input n_2358;
input n_1255;
input n_568;
input n_1516;
input n_143;
input n_1536;
input n_180;
input n_2163;
input n_2186;
input n_2029;
input n_2815;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_2528;
input n_2814;
input n_214;
input n_246;
input n_2787;
input n_1338;
input n_1097;
input n_2395;
input n_935;
input n_781;
input n_789;
input n_1554;
input n_1130;
input n_181;
input n_1810;
input n_182;
input n_573;
input n_769;
input n_2380;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_1583;
input n_1730;
input n_2295;
input n_555;
input n_389;
input n_814;
input n_2746;
input n_1643;
input n_2020;
input n_2500;
input n_2269;
input n_1729;
input n_669;
input n_2290;
input n_2048;
input n_176;
input n_114;
input n_300;
input n_222;
input n_2005;
input n_747;
input n_74;
input n_2565;
input n_1389;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_535;
input n_691;
input n_372;
input n_2076;
input n_2736;
input n_111;
input n_2883;
input n_314;
input n_1408;
input n_378;
input n_1196;
input n_377;
input n_1598;
input n_863;
input n_2175;
input n_601;
input n_2182;
input n_338;
input n_2910;
input n_1283;
input n_2385;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_1785;
input n_56;
input n_763;
input n_1147;
input n_1848;
input n_360;
input n_1754;
input n_2149;
input n_2396;
input n_1506;
input n_119;
input n_2584;
input n_1652;
input n_1812;
input n_957;
input n_1994;
input n_895;
input n_866;
input n_1227;
input n_2450;
input n_2485;
input n_2284;
input n_191;
input n_2566;
input n_387;
input n_2287;
input n_452;
input n_744;
input n_971;
input n_2702;
input n_946;
input n_344;
input n_2906;
input n_761;
input n_1303;
input n_2769;
input n_1205;
input n_2492;
input n_1258;
input n_2438;
input n_2914;
input n_1392;
input n_174;
input n_1173;
input n_1924;
input n_525;
input n_2463;
input n_2881;
input n_1677;
input n_1116;
input n_611;
input n_1570;
input n_1702;
input n_1219;
input n_1780;
input n_1689;
input n_8;
input n_2180;
input n_2858;
input n_2679;
input n_1174;
input n_1944;
input n_1016;
input n_1347;
input n_795;
input n_1501;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_2117;
input n_2234;
input n_2779;
input n_2685;
input n_1083;
input n_109;
input n_445;
input n_1561;
input n_2741;
input n_930;
input n_888;
input n_2275;
input n_1112;
input n_2465;
input n_2620;
input n_2081;
input n_2168;
input n_2568;
input n_234;
input n_2022;
input n_1945;
input n_2203;
input n_910;
input n_1656;
input n_1721;
input n_1460;
input n_911;
input n_2112;
input n_2255;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1737;
input n_2430;
input n_1414;
input n_752;
input n_908;
input n_2649;
input n_2721;
input n_944;
input n_2034;
input n_576;
input n_1028;
input n_2106;
input n_472;
input n_2862;
input n_270;
input n_2265;
input n_2615;
input n_414;
input n_2683;
input n_1922;
input n_563;
input n_2032;
input n_2744;
input n_1011;
input n_2474;
input n_1566;
input n_1215;
input n_2437;
input n_25;
input n_93;
input n_839;
input n_2444;
input n_2743;
input n_708;
input n_1973;
input n_2267;
input n_668;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1821;
input n_2205;
input n_1104;
input n_854;
input n_1058;
input n_2312;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_2242;
input n_1509;
input n_103;
input n_1693;
input n_1109;
input n_185;
input n_2222;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_2015;
input n_2118;
input n_2111;
input n_2466;
input n_390;
input n_2915;
input n_2530;
input n_1148;
input n_31;
input n_2188;
input n_2505;
input n_334;
input n_1989;
input n_1161;
input n_2609;
input n_1085;
input n_232;
input n_2802;
input n_2014;
input n_2042;
input n_46;
input n_1239;
input n_771;
input n_1584;
input n_2425;
input n_470;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_2318;
input n_2408;
input n_1149;
input n_265;
input n_1184;
input n_2483;
input n_228;
input n_719;
input n_1972;
input n_2592;
input n_1525;
input n_2594;
input n_455;
input n_2666;
input n_1585;
input n_1851;
input n_363;
input n_1799;
input n_1090;
input n_2147;
input n_2564;
input n_592;
input n_1816;
input n_2503;
input n_2433;
input n_1518;
input n_829;
input n_1156;
input n_1362;
input n_393;
input n_984;
input n_2600;
input n_1829;
input n_503;
input n_2035;
input n_1450;
input n_1638;
input n_132;
input n_868;
input n_570;
input n_859;
input n_2033;
input n_406;
input n_735;
input n_1789;
input n_2531;
input n_1770;
input n_878;
input n_620;
input n_130;
input n_519;
input n_2523;
input n_307;
input n_469;
input n_1218;
input n_2413;
input n_500;
input n_1482;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_2071;
input n_357;
input n_2429;
input n_985;
input n_2233;
input n_2440;
input n_2723;
input n_481;
input n_997;
input n_1710;
input n_2800;
input n_2161;
input n_1301;
input n_2805;
input n_802;
input n_561;
input n_33;
input n_980;
input n_2681;
input n_1306;
input n_2010;
input n_2282;
input n_1651;
input n_1198;
input n_2360;
input n_2047;
input n_2651;
input n_2095;
input n_1609;
input n_2174;
input n_2799;
input n_436;
input n_116;
input n_2334;
input n_409;
input n_1244;
input n_1685;
input n_1763;
input n_1998;
input n_1574;
input n_2426;
input n_2490;
input n_2844;
input n_240;
input n_756;
input n_2303;
input n_1619;
input n_2478;
input n_1981;
input n_2285;
input n_1606;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_2742;
input n_2640;
input n_1051;
input n_253;
input n_1552;
input n_2918;
input n_583;
input n_1996;
input n_2367;
input n_249;
input n_201;
input n_2867;
input n_1039;
input n_1442;
input n_2726;
input n_1034;
input n_2043;
input n_1480;
input n_1158;
input n_2909;
input n_2248;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_1305;
input n_2363;
input n_2578;
input n_553;
input n_43;
input n_849;
input n_2662;
input n_753;
input n_1753;
input n_2795;
input n_2471;
input n_467;
input n_2540;
input n_269;
input n_359;
input n_973;
input n_2807;
input n_1921;
input n_1479;
input n_1055;
input n_1675;
input n_2197;
input n_2217;
input n_582;
input n_2065;
input n_2879;
input n_861;
input n_857;
input n_967;
input n_571;
input n_2215;
input n_2461;
input n_271;
input n_404;
input n_2001;
input n_158;
input n_2107;
input n_1884;
input n_206;
input n_2040;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_1629;
input n_2221;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1819;
input n_2055;
input n_1010;
input n_2553;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_2038;
input n_812;
input n_2891;
input n_1131;
input n_2634;
input n_1761;
input n_2709;
input n_534;
input n_1578;
input n_1006;
input n_1861;
input n_373;
input n_87;
input n_1632;
input n_1890;
input n_1805;
input n_2477;
input n_257;
input n_1557;
input n_1888;
input n_2280;
input n_1833;
input n_730;
input n_1311;
input n_1494;
input n_2325;
input n_670;
input n_203;
input n_1850;
input n_1898;
input n_2443;
input n_2697;
input n_2308;
input n_2162;
input n_1868;
input n_207;
input n_2333;
input n_2079;
input n_1089;
input n_1887;
input n_1587;
input n_2512;
input n_1365;
input n_1417;
input n_205;
input n_1242;
input n_2086;
input n_2185;
input n_1836;
input n_2774;
input n_681;
input n_1226;
input n_1274;
input n_1486;
input n_2166;
input n_412;
input n_2899;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_1899;
input n_1428;
input n_1616;
input n_1576;
input n_1856;
input n_1862;
input n_1958;
input n_2077;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_2632;
input n_422;
input n_2579;
input n_722;
input n_862;
input n_2105;
input n_135;
input n_165;
input n_2098;
input n_540;
input n_1423;
input n_2813;
input n_1935;
input n_2027;
input n_457;
input n_2223;
input n_2091;
input n_364;
input n_1915;
input n_629;
input n_1621;
input n_1748;
input n_2547;
input n_2415;
input n_900;
input n_1449;
input n_531;
input n_827;
input n_2912;
input n_60;
input n_361;
input n_2659;
input n_1025;
input n_2419;
input n_2116;
input n_336;
input n_2320;
input n_12;
input n_1885;
input n_2677;
input n_1013;
input n_1259;
input n_192;
input n_2183;
input n_1538;
input n_51;
input n_649;
input n_1612;
input n_1240;

output n_13275;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_4452;
wire n_6566;
wire n_13045;
wire n_5172;
wire n_11173;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_6872;
wire n_5254;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_13146;
wire n_13235;
wire n_10587;
wire n_5019;
wire n_8713;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_3849;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_5138;
wire n_10931;
wire n_4388;
wire n_4395;
wire n_6960;
wire n_3089;
wire n_8169;
wire n_12265;
wire n_9002;
wire n_9130;
wire n_7180;
wire n_5653;
wire n_11574;
wire n_4978;
wire n_8604;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_13125;
wire n_3088;
wire n_8168;
wire n_3257;
wire n_4829;
wire n_5393;
wire n_3222;
wire n_7190;
wire n_7504;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_4686;
wire n_12322;
wire n_8899;
wire n_5524;
wire n_10236;
wire n_5345;
wire n_11205;
wire n_11678;
wire n_11776;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_11650;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_8534;
wire n_5963;
wire n_12179;
wire n_5055;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_11905;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_4249;
wire n_11536;
wire n_5950;
wire n_3564;
wire n_9104;
wire n_6999;
wire n_11046;
wire n_11079;
wire n_10283;
wire n_5548;
wire n_5057;
wire n_11065;
wire n_8339;
wire n_8272;
wire n_7161;
wire n_3030;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_3427;
wire n_11214;
wire n_5101;
wire n_3071;
wire n_7000;
wire n_8561;
wire n_11954;
wire n_7398;
wire n_2926;
wire n_10392;
wire n_12882;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_12617;
wire n_8411;
wire n_8499;
wire n_8236;
wire n_5102;
wire n_13137;
wire n_3345;
wire n_13221;
wire n_6882;
wire n_10775;
wire n_4501;
wire n_9626;
wire n_11163;
wire n_9526;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_5598;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_7389;
wire n_4997;
wire n_10719;
wire n_11419;
wire n_9018;
wire n_4843;
wire n_12095;
wire n_8070;
wire n_4696;
wire n_6660;
wire n_9055;
wire n_4347;
wire n_11740;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_7008;
wire n_3877;
wire n_12392;
wire n_3929;
wire n_8366;
wire n_3048;
wire n_8102;
wire n_9362;
wire n_11979;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_5894;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_10239;
wire n_5332;
wire n_9962;
wire n_4814;
wire n_5908;
wire n_3979;
wire n_10373;
wire n_3077;
wire n_11104;
wire n_3452;
wire n_8913;
wire n_9525;
wire n_3107;
wire n_10816;
wire n_9725;
wire n_4956;
wire n_11537;
wire n_12707;
wire n_7686;
wire n_3664;
wire n_6914;
wire n_10335;
wire n_5337;
wire n_5129;
wire n_11301;
wire n_12424;
wire n_5420;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_11703;
wire n_11699;
wire n_4646;
wire n_6374;
wire n_7651;
wire n_11543;
wire n_10947;
wire n_6628;
wire n_8125;
wire n_3760;
wire n_6015;
wire n_11261;
wire n_10226;
wire n_13247;
wire n_4262;
wire n_6526;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_3347;
wire n_10767;
wire n_5136;
wire n_8040;
wire n_11821;
wire n_5638;
wire n_13121;
wire n_9100;
wire n_4110;
wire n_6784;
wire n_12107;
wire n_10755;
wire n_4950;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_6323;
wire n_9614;
wire n_10682;
wire n_6110;
wire n_11684;
wire n_3999;
wire n_12652;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_10699;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_9400;
wire n_5151;
wire n_8142;
wire n_11627;
wire n_5684;
wire n_8598;
wire n_13139;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_7856;
wire n_7774;
wire n_5680;
wire n_6674;
wire n_6148;
wire n_6951;
wire n_11659;
wire n_7625;
wire n_4102;
wire n_3871;
wire n_9106;
wire n_12775;
wire n_4662;
wire n_8869;
wire n_6989;
wire n_4671;
wire n_7863;
wire n_3959;
wire n_8381;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_9520;
wire n_8958;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_12371;
wire n_4296;
wire n_10114;
wire n_12203;
wire n_10357;
wire n_7147;
wire n_8115;
wire n_4507;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_11497;
wire n_3484;
wire n_12359;
wire n_4677;
wire n_12915;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_13149;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_12742;
wire n_3923;
wire n_9042;
wire n_11768;
wire n_3900;
wire n_8412;
wire n_9267;
wire n_3488;
wire n_3732;
wire n_6485;
wire n_8987;
wire n_11805;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_4226;
wire n_5493;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_12770;
wire n_10012;
wire n_4294;
wire n_12985;
wire n_4698;
wire n_4445;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_7564;
wire n_11635;
wire n_3859;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_4456;
wire n_3914;
wire n_8119;
wire n_10296;
wire n_3397;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_9718;
wire n_9128;
wire n_10281;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_8748;
wire n_3927;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_6794;
wire n_6151;
wire n_3888;
wire n_8718;
wire n_7110;
wire n_5476;
wire n_12831;
wire n_9935;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_2922;
wire n_8223;
wire n_3882;
wire n_4856;
wire n_10097;
wire n_3492;
wire n_4369;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_4331;
wire n_7297;
wire n_9866;
wire n_10018;
wire n_4972;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_12427;
wire n_7533;
wire n_7221;
wire n_4375;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_11295;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_11662;
wire n_5532;
wire n_5897;
wire n_8246;
wire n_8952;
wire n_4613;
wire n_13014;
wire n_9070;
wire n_11708;
wire n_3012;
wire n_3875;
wire n_10266;
wire n_5609;
wire n_4717;
wire n_10897;
wire n_10827;
wire n_4877;
wire n_3247;
wire n_5922;
wire n_10449;
wire n_7569;
wire n_7823;
wire n_7734;
wire n_7062;
wire n_7861;
wire n_8955;
wire n_9477;
wire n_5658;
wire n_4731;
wire n_9680;
wire n_12172;
wire n_12147;
wire n_12923;
wire n_3052;
wire n_7039;
wire n_8577;
wire n_12384;
wire n_11349;
wire n_8594;
wire n_5046;
wire n_13227;
wire n_8428;
wire n_9829;
wire n_11260;
wire n_3298;
wire n_8848;
wire n_12825;
wire n_5058;
wire n_10685;
wire n_11351;
wire n_3273;
wire n_4467;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_5667;
wire n_8259;
wire n_12540;
wire n_10607;
wire n_5865;
wire n_12249;
wire n_8349;
wire n_6836;
wire n_5042;
wire n_5305;
wire n_11998;
wire n_4681;
wire n_8164;
wire n_13239;
wire n_4072;
wire n_10628;
wire n_4752;
wire n_4220;
wire n_7905;
wire n_5281;
wire n_8776;
wire n_11775;
wire n_9143;
wire n_8287;
wire n_10256;
wire n_10769;
wire n_7753;
wire n_10368;
wire n_6771;
wire n_7950;
wire n_9947;
wire n_9088;
wire n_8607;
wire n_10138;
wire n_12117;
wire n_11706;
wire n_6248;
wire n_11800;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_6795;
wire n_5314;
wire n_10452;
wire n_11464;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_12960;
wire n_13033;
wire n_11642;
wire n_4381;
wire n_11143;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_3968;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_12131;
wire n_12851;
wire n_5795;
wire n_11934;
wire n_12349;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_8416;
wire n_10396;
wire n_4518;
wire n_10724;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_9988;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_12740;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_10363;
wire n_13240;
wire n_3237;
wire n_8949;
wire n_10831;
wire n_3500;
wire n_3834;
wire n_9131;
wire n_11553;
wire n_10517;
wire n_12578;
wire n_12795;
wire n_4589;
wire n_10323;
wire n_12194;
wire n_2972;
wire n_10842;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_10876;
wire n_11511;
wire n_9137;
wire n_11180;
wire n_9724;
wire n_11146;
wire n_9281;
wire n_3192;
wire n_8995;
wire n_10883;
wire n_10101;
wire n_9393;
wire n_4394;
wire n_6581;
wire n_12709;
wire n_6010;
wire n_3352;
wire n_8711;
wire n_3073;
wire n_7013;
wire n_12771;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_3696;
wire n_4082;
wire n_7290;
wire n_12278;
wire n_10820;
wire n_4921;
wire n_9687;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_7315;
wire n_13194;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_4697;
wire n_13244;
wire n_4289;
wire n_4288;
wire n_11866;
wire n_3763;
wire n_6185;
wire n_11450;
wire n_12522;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_9102;
wire n_11526;
wire n_9578;
wire n_3614;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_7438;
wire n_7268;
wire n_7337;
wire n_11851;
wire n_4964;
wire n_9489;
wire n_12804;
wire n_5957;
wire n_6965;
wire n_12116;
wire n_10728;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_10094;
wire n_9144;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_7461;
wire n_8285;
wire n_4322;
wire n_10655;
wire n_3644;
wire n_9797;
wire n_6955;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_4287;
wire n_4137;
wire n_9521;
wire n_8332;
wire n_9478;
wire n_9932;
wire n_13040;
wire n_7278;
wire n_6509;
wire n_11370;
wire n_4576;
wire n_7454;
wire n_11253;
wire n_11379;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_11981;
wire n_3179;
wire n_3400;
wire n_9895;
wire n_8741;
wire n_12918;
wire n_4000;
wire n_9351;
wire n_11585;
wire n_5445;
wire n_13140;
wire n_4389;
wire n_5342;
wire n_5501;
wire n_6839;
wire n_3970;
wire n_7377;
wire n_4345;
wire n_7232;
wire n_6646;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_9189;
wire n_4664;
wire n_4156;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_7904;
wire n_11691;
wire n_6033;
wire n_11541;
wire n_3158;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_5748;
wire n_3782;
wire n_9356;
wire n_12865;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_3700;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_10959;
wire n_3104;
wire n_6809;
wire n_11233;
wire n_3435;
wire n_5636;
wire n_7840;
wire n_10972;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_13213;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_7080;
wire n_6636;
wire n_5286;
wire n_8229;
wire n_4528;
wire n_8410;
wire n_5811;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_7624;
wire n_4914;
wire n_4939;
wire n_7629;
wire n_3418;
wire n_9735;
wire n_9186;
wire n_10818;
wire n_5530;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_12552;
wire n_11069;
wire n_4096;
wire n_5595;
wire n_4123;
wire n_9941;
wire n_11951;
wire n_7003;
wire n_12222;
wire n_11900;
wire n_3119;
wire n_5427;
wire n_10788;
wire n_3735;
wire n_11369;
wire n_4379;
wire n_10563;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_5901;
wire n_6538;
wire n_5962;
wire n_5599;
wire n_3631;
wire n_7010;
wire n_8107;
wire n_11108;
wire n_9728;
wire n_12883;
wire n_11004;
wire n_12992;
wire n_5324;
wire n_6519;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_3770;
wire n_9818;
wire n_6530;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_4440;
wire n_8774;
wire n_4402;
wire n_10566;
wire n_10178;
wire n_5052;
wire n_7299;
wire n_12367;
wire n_4541;
wire n_12104;
wire n_5009;
wire n_4872;
wire n_6402;
wire n_12469;
wire n_9936;
wire n_12563;
wire n_4551;
wire n_6195;
wire n_13132;
wire n_7243;
wire n_6609;
wire n_7326;
wire n_9530;
wire n_10115;
wire n_5326;
wire n_7471;
wire n_7067;
wire n_10455;
wire n_11778;
wire n_12793;
wire n_4627;
wire n_4079;
wire n_5300;
wire n_9909;
wire n_11393;
wire n_8691;
wire n_8620;
wire n_12406;
wire n_3342;
wire n_6748;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_13270;
wire n_7790;
wire n_11719;
wire n_6149;
wire n_10052;
wire n_10109;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_11963;
wire n_12428;
wire n_8424;
wire n_9571;
wire n_3025;
wire n_8026;
wire n_9638;
wire n_7528;
wire n_9470;
wire n_4798;
wire n_3810;
wire n_3006;
wire n_10265;
wire n_8174;
wire n_12655;
wire n_7941;
wire n_11175;
wire n_5010;
wire n_11483;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_5089;
wire n_11371;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_6264;
wire n_8861;
wire n_5359;
wire n_8644;
wire n_8907;
wire n_12304;
wire n_11080;
wire n_10984;
wire n_5137;
wire n_6902;
wire n_3331;
wire n_5104;
wire n_10100;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7913;
wire n_7478;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_3606;
wire n_12692;
wire n_3591;
wire n_7939;
wire n_8503;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_6449;
wire n_6723;
wire n_7458;
wire n_9108;
wire n_9787;
wire n_6440;
wire n_7436;
wire n_10846;
wire n_4746;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_8446;
wire n_5194;
wire n_9376;
wire n_9786;
wire n_9033;
wire n_12933;
wire n_7435;
wire n_12908;
wire n_3441;
wire n_9537;
wire n_11297;
wire n_3534;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_12996;
wire n_5947;
wire n_8923;
wire n_12643;
wire n_6736;
wire n_6124;
wire n_3944;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_5985;
wire n_8197;
wire n_3605;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_3306;
wire n_12827;
wire n_12678;
wire n_9115;
wire n_3026;
wire n_12235;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_11833;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_5001;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_9938;
wire n_11285;
wire n_8082;
wire n_12098;
wire n_4428;
wire n_8730;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_9203;
wire n_9977;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_5761;
wire n_9242;
wire n_6773;
wire n_4618;
wire n_12611;
wire n_13269;
wire n_7375;
wire n_4679;
wire n_3479;
wire n_11262;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_12713;
wire n_12880;
wire n_13144;
wire n_4805;
wire n_8651;
wire n_3454;
wire n_9141;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_6531;
wire n_10952;
wire n_10851;
wire n_11027;
wire n_11852;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_10221;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_11803;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_5100;
wire n_9286;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_8281;
wire n_10819;
wire n_3816;
wire n_4807;
wire n_8842;
wire n_4411;
wire n_9184;
wire n_3214;
wire n_9704;
wire n_2928;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_8024;
wire n_7730;
wire n_12562;
wire n_8814;
wire n_8530;
wire n_11428;
wire n_11592;
wire n_4180;
wire n_9193;
wire n_8467;
wire n_11677;
wire n_7281;
wire n_3109;
wire n_9717;
wire n_3354;
wire n_7711;
wire n_3126;
wire n_11090;
wire n_8984;
wire n_3663;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_9290;
wire n_5740;
wire n_5820;
wire n_5648;
wire n_13266;
wire n_5745;
wire n_4707;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_9875;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_8676;
wire n_5534;
wire n_8003;
wire n_4880;
wire n_8785;
wire n_9853;
wire n_13192;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_4126;
wire n_3845;
wire n_6556;
wire n_8692;
wire n_6889;
wire n_7230;
wire n_9183;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_9778;
wire n_5196;
wire n_6199;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_10852;
wire n_4470;
wire n_6726;
wire n_12374;
wire n_13200;
wire n_9529;
wire n_4813;
wire n_5542;
wire n_3901;
wire n_7011;
wire n_8998;
wire n_10538;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_4014;
wire n_4704;
wire n_11066;
wire n_10315;
wire n_4252;
wire n_9123;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_4048;
wire n_4596;
wire n_12368;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_3406;
wire n_13193;
wire n_6100;
wire n_12796;
wire n_6516;
wire n_3919;
wire n_8462;
wire n_6977;
wire n_9380;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_12529;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_8979;
wire n_6522;
wire n_4952;
wire n_5023;
wire n_5906;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_5660;
wire n_3981;
wire n_7890;
wire n_12785;
wire n_3973;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_12461;
wire n_6808;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_6207;
wire n_7006;
wire n_6931;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_9082;
wire n_10925;
wire n_4770;
wire n_9879;
wire n_11158;
wire n_3474;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_4690;
wire n_11669;
wire n_3864;
wire n_8264;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_12078;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_10618;
wire n_8135;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_3592;
wire n_11739;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_10497;
wire n_9445;
wire n_7627;
wire n_9803;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_3195;
wire n_6346;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_8408;
wire n_12639;
wire n_3277;
wire n_5386;
wire n_10661;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_3817;
wire n_10028;
wire n_7811;
wire n_13158;
wire n_11676;
wire n_11044;
wire n_11771;
wire n_12266;
wire n_3659;
wire n_12175;
wire n_5003;
wire n_10512;
wire n_11384;
wire n_4827;
wire n_12287;
wire n_11679;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_12353;
wire n_3042;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_12398;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_9087;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_9043;
wire n_6075;
wire n_12991;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_10789;
wire n_11134;
wire n_12705;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_11828;
wire n_12326;
wire n_7847;
wire n_8506;
wire n_3464;
wire n_6494;
wire n_13178;
wire n_6133;
wire n_3723;
wire n_11548;
wire n_13041;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_7822;
wire n_6453;
wire n_4380;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_6127;
wire n_10762;
wire n_11342;
wire n_4398;
wire n_11452;
wire n_11362;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_5031;
wire n_6006;
wire n_10797;
wire n_7289;
wire n_4193;
wire n_11266;
wire n_3570;
wire n_12309;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_5338;
wire n_3828;
wire n_12479;
wire n_7354;
wire n_8352;
wire n_12502;
wire n_3424;
wire n_4131;
wire n_10360;
wire n_7960;
wire n_9450;
wire n_3594;
wire n_5689;
wire n_7482;
wire n_12912;
wire n_10312;
wire n_4090;
wire n_12211;
wire n_6115;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_9223;
wire n_13191;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_10131;
wire n_12537;
wire n_6838;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_11988;
wire n_12600;
wire n_12921;
wire n_13226;
wire n_3485;
wire n_5931;
wire n_6139;
wire n_4077;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_6256;
wire n_7965;
wire n_3262;
wire n_6613;
wire n_11438;
wire n_11244;
wire n_4008;
wire n_12919;
wire n_3356;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_3210;
wire n_6361;
wire n_9880;
wire n_13253;
wire n_4689;
wire n_8183;
wire n_11348;
wire n_4547;
wire n_11245;
wire n_9685;
wire n_6085;
wire n_7474;
wire n_11169;
wire n_11685;
wire n_5731;
wire n_12422;
wire n_6329;
wire n_11607;
wire n_8650;
wire n_6678;
wire n_11546;
wire n_3329;
wire n_8662;
wire n_10503;
wire n_9694;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_13215;
wire n_4601;
wire n_9905;
wire n_9948;
wire n_10465;
wire n_12429;
wire n_10590;
wire n_3647;
wire n_3681;
wire n_4300;
wire n_8526;
wire n_4623;
wire n_7325;
wire n_10887;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_5883;
wire n_7166;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_6560;
wire n_11319;
wire n_3476;
wire n_7028;
wire n_4842;
wire n_7838;
wire n_9890;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_11492;
wire n_7873;
wire n_6535;
wire n_12731;
wire n_12399;
wire n_7518;
wire n_12342;
wire n_7414;
wire n_9817;
wire n_9744;
wire n_6147;
wire n_9199;
wire n_10063;
wire n_12640;
wire n_9548;
wire n_8973;
wire n_11160;
wire n_6448;
wire n_7791;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_12533;
wire n_3292;
wire n_9862;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_12616;
wire n_11385;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_12535;
wire n_3437;
wire n_12178;
wire n_4111;
wire n_12653;
wire n_6643;
wire n_12327;
wire n_7146;
wire n_9471;
wire n_4608;
wire n_3712;
wire n_11346;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_9069;
wire n_13110;
wire n_5852;
wire n_3562;
wire n_2973;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_8249;
wire n_7052;
wire n_11343;
wire n_12348;
wire n_3665;
wire n_10496;
wire n_3007;
wire n_12257;
wire n_3528;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_4571;
wire n_10843;
wire n_3698;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_3355;
wire n_8234;
wire n_3174;
wire n_5321;
wire n_9960;
wire n_10997;
wire n_4215;
wire n_9010;
wire n_10998;
wire n_9003;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_12418;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_7312;
wire n_13263;
wire n_7919;
wire n_5145;
wire n_4219;
wire n_11269;
wire n_10800;
wire n_7085;
wire n_11491;
wire n_12065;
wire n_3958;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_11408;
wire n_3985;
wire n_11772;
wire n_4196;
wire n_4774;
wire n_5210;
wire n_13183;
wire n_6689;
wire n_10993;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12519;
wire n_9172;
wire n_12769;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_5149;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_11311;
wire n_10112;
wire n_10765;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_11792;
wire n_7304;
wire n_3713;
wire n_9734;
wire n_7288;
wire n_8558;
wire n_13242;
wire n_10489;
wire n_7707;
wire n_3197;
wire n_7223;
wire n_12421;
wire n_7833;
wire n_12113;
wire n_4987;
wire n_5512;
wire n_7274;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_4736;
wire n_3743;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_3124;
wire n_10612;
wire n_11086;
wire n_7466;
wire n_6529;
wire n_10260;
wire n_11293;
wire n_3759;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_12285;
wire n_11710;
wire n_8619;
wire n_11568;
wire n_3511;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_9150;
wire n_10134;
wire n_11603;
wire n_7277;
wire n_6455;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_13099;
wire n_12015;
wire n_8146;
wire n_4492;
wire n_8813;
wire n_5607;
wire n_11562;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_10194;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_12157;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_8910;
wire n_12311;
wire n_4376;
wire n_6203;
wire n_6408;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_13064;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_4708;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_12031;
wire n_5341;
wire n_8643;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_11718;
wire n_8565;
wire n_10821;
wire n_11170;
wire n_11758;
wire n_12126;
wire n_8550;
wire n_4081;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_7322;
wire n_9053;
wire n_11658;
wire n_11893;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_4536;
wire n_9480;
wire n_5562;
wire n_3303;
wire n_4324;
wire n_7051;
wire n_10850;
wire n_8477;
wire n_9185;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_4382;
wire n_12195;
wire n_13115;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_5911;
wire n_3954;
wire n_11601;
wire n_11971;
wire n_13182;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_5622;
wire n_3503;
wire n_9919;
wire n_3160;
wire n_12135;
wire n_6574;
wire n_11116;
wire n_12604;
wire n_6571;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_8876;
wire n_5124;
wire n_9151;
wire n_3951;
wire n_8829;
wire n_7824;
wire n_9359;
wire n_13236;
wire n_3569;
wire n_7094;
wire n_3874;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8140;
wire n_8971;
wire n_8060;
wire n_10558;
wire n_3027;
wire n_7036;
wire n_4083;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_6392;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_9049;
wire n_7351;
wire n_4480;
wire n_9352;
wire n_7608;
wire n_5779;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_13202;
wire n_7909;
wire n_7413;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_11340;
wire n_10734;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_11903;
wire n_7027;
wire n_7992;
wire n_6912;
wire n_11560;
wire n_10395;
wire n_7175;
wire n_8276;
wire n_3617;
wire n_10330;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_3567;
wire n_11465;
wire n_7524;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_11564;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_11265;
wire n_9370;
wire n_11125;
wire n_9670;
wire n_13136;
wire n_4027;
wire n_12916;
wire n_3154;
wire n_9334;
wire n_7783;
wire n_13220;
wire n_6692;
wire n_3898;
wire n_10276;
wire n_12331;
wire n_3520;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_12531;
wire n_8245;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_12521;
wire n_11302;
wire n_12910;
wire n_9956;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_10991;
wire n_10098;
wire n_11745;
wire n_8891;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_11690;
wire n_9487;
wire n_3897;
wire n_11707;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_7697;
wire n_6403;
wire n_7306;
wire n_7947;
wire n_10118;
wire n_7470;
wire n_7547;
wire n_6013;
wire n_7733;
wire n_7693;
wire n_9557;
wire n_3215;
wire n_6491;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_13039;
wire n_13130;
wire n_8582;
wire n_10441;
wire n_5518;
wire n_6982;
wire n_10002;
wire n_5068;
wire n_6293;
wire n_9124;
wire n_6661;
wire n_5847;
wire n_7345;
wire n_6049;
wire n_9762;
wire n_8847;
wire n_11242;
wire n_8957;
wire n_7385;
wire n_10923;
wire n_5159;
wire n_4068;
wire n_6558;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_3703;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_12313;
wire n_3962;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_9543;
wire n_3035;
wire n_4166;
wire n_11396;
wire n_8356;
wire n_6136;
wire n_9660;
wire n_11443;
wire n_9483;
wire n_3378;
wire n_6855;
wire n_3745;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_6091;
wire n_3667;
wire n_3523;
wire n_13093;
wire n_13062;
wire n_9328;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_6312;
wire n_8747;
wire n_11532;
wire n_9539;
wire n_4817;
wire n_6668;
wire n_9415;
wire n_4115;
wire n_2999;
wire n_9385;
wire n_3697;
wire n_9147;
wire n_11209;
wire n_7653;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_13185;
wire n_9027;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_4383;
wire n_6995;
wire n_10902;
wire n_4491;
wire n_12889;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_4486;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_11304;
wire n_9642;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_3024;
wire n_7475;
wire n_10485;
wire n_12105;
wire n_4612;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_13219;
wire n_5673;
wire n_5443;
wire n_6351;
wire n_9079;
wire n_9382;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_10444;
wire n_4529;
wire n_3361;
wire n_11377;
wire n_3478;
wire n_8018;
wire n_8653;
wire n_3936;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_5823;
wire n_7305;
wire n_3496;
wire n_13160;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_4390;
wire n_12248;
wire n_3096;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_8884;
wire n_8803;
wire n_3239;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_5537;
wire n_10978;
wire n_8222;
wire n_6822;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_11715;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_9706;
wire n_3101;
wire n_10642;
wire n_4233;
wire n_12181;
wire n_10187;
wire n_3374;
wire n_10387;
wire n_11014;
wire n_3288;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_11864;
wire n_3876;
wire n_11007;
wire n_11224;
wire n_11006;
wire n_9564;
wire n_3125;
wire n_7391;
wire n_8790;
wire n_9230;
wire n_6617;
wire n_4293;
wire n_10219;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_4684;
wire n_3116;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_10364;
wire n_10479;
wire n_11422;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_4412;
wire n_8178;
wire n_6801;
wire n_12489;
wire n_8491;
wire n_3618;
wire n_4580;
wire n_5630;
wire n_4758;
wire n_10065;
wire n_4781;
wire n_12046;
wire n_10212;
wire n_9283;
wire n_8700;
wire n_4148;
wire n_12030;
wire n_12738;
wire n_4057;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_10268;
wire n_3444;
wire n_3059;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_12601;
wire n_9425;
wire n_12917;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_3017;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_10559;
wire n_13173;
wire n_8439;
wire n_3001;
wire n_9641;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_12059;
wire n_12488;
wire n_3795;
wire n_7321;
wire n_5289;
wire n_3852;
wire n_4138;
wire n_8200;
wire n_11110;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_8304;
wire n_3815;
wire n_3896;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_3274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_4457;
wire n_7537;
wire n_10516;
wire n_4093;
wire n_8675;
wire n_10892;
wire n_6254;
wire n_5989;
wire n_10493;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_4794;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_9016;
wire n_13101;
wire n_11887;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_11545;
wire n_9729;
wire n_5073;
wire n_12691;
wire n_8846;
wire n_8315;
wire n_12471;
wire n_11033;
wire n_12451;
wire n_4834;
wire n_11040;
wire n_12665;
wire n_11754;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_4762;
wire n_5581;
wire n_9411;
wire n_9029;
wire n_11672;
wire n_3113;
wire n_6837;
wire n_10353;
wire n_3813;
wire n_3660;
wire n_10847;
wire n_12651;
wire n_3766;
wire n_10451;
wire n_11043;
wire n_5303;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_9414;
wire n_3266;
wire n_7023;
wire n_3574;
wire n_9615;
wire n_12003;
wire n_7496;
wire n_11277;
wire n_4154;
wire n_12165;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_10866;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_3844;
wire n_8777;
wire n_4975;
wire n_11061;
wire n_11763;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_8535;
wire n_10653;
wire n_11534;
wire n_6373;
wire n_5375;
wire n_11587;
wire n_12280;
wire n_9221;
wire n_12492;
wire n_12972;
wire n_5370;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_9811;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_13188;
wire n_4819;
wire n_7906;
wire n_5248;
wire n_9951;
wire n_7131;
wire n_6411;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_11032;
wire n_5112;
wire n_3332;
wire n_4134;
wire n_10507;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_11843;
wire n_4092;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_7797;
wire n_3668;
wire n_11335;
wire n_11629;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_7687;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_5635;
wire n_4087;
wire n_7582;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_4302;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_11698;
wire n_6534;
wire n_3340;
wire n_10614;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_2989;
wire n_5778;
wire n_8425;
wire n_11257;
wire n_8087;
wire n_9910;
wire n_3395;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_11801;
wire n_13217;
wire n_12073;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_10743;
wire n_5165;
wire n_4884;
wire n_10853;
wire n_7867;
wire n_9651;
wire n_3275;
wire n_10249;
wire n_8361;
wire n_6135;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_10270;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_3440;
wire n_11115;
wire n_8669;
wire n_12978;
wire n_8001;
wire n_7525;
wire n_7257;
wire n_12363;
wire n_9372;
wire n_7553;
wire n_7529;
wire n_4692;
wire n_6791;
wire n_8496;
wire n_3165;
wire n_11915;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_11788;
wire n_12544;
wire n_3890;
wire n_13036;
wire n_3750;
wire n_3607;
wire n_7650;
wire n_12476;
wire n_13199;
wire n_3316;
wire n_8568;
wire n_6903;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_4311;
wire n_12023;
wire n_8637;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_13002;
wire n_3261;
wire n_12632;
wire n_12620;
wire n_7520;
wire n_9831;
wire n_13203;
wire n_4187;
wire n_6309;
wire n_7903;
wire n_9697;
wire n_11303;
wire n_11877;
wire n_6733;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_5430;
wire n_8610;
wire n_5942;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_9902;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_3532;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_9039;
wire n_12598;
wire n_11854;
wire n_12416;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_8265;
wire n_4619;
wire n_7639;
wire n_8704;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_11609;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_13230;
wire n_9294;
wire n_5036;
wire n_12811;
wire n_4221;
wire n_3297;
wire n_12186;
wire n_11747;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_12494;
wire n_13032;
wire n_7054;
wire n_7605;
wire n_3067;
wire n_11556;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_11529;
wire n_5327;
wire n_10021;
wire n_9146;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_2996;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_3803;
wire n_8941;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_9073;
wire n_10075;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_8775;
wire n_12272;
wire n_9302;
wire n_5519;
wire n_11798;
wire n_9062;
wire n_11895;
wire n_6269;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_3412;
wire n_8279;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_12191;
wire n_9580;
wire n_8019;
wire n_9972;
wire n_3791;
wire n_13003;
wire n_6083;
wire n_13091;
wire n_12909;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_4320;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_3884;
wire n_9465;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_5231;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_3438;
wire n_4141;
wire n_10436;
wire n_8464;
wire n_6547;
wire n_8799;
wire n_12794;
wire n_5193;
wire n_6423;
wire n_9442;
wire n_6342;
wire n_6641;
wire n_6984;
wire n_12467;
wire n_3373;
wire n_5789;
wire n_10763;
wire n_7441;
wire n_9957;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_12112;
wire n_13060;
wire n_3883;
wire n_10245;
wire n_5961;
wire n_10905;
wire n_11235;
wire n_9449;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_6687;
wire n_9313;
wire n_5822;
wire n_9173;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_5726;
wire n_3949;
wire n_9563;
wire n_11015;
wire n_9160;
wire n_5364;
wire n_9974;
wire n_12129;
wire n_11166;
wire n_3315;
wire n_7031;
wire n_9285;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_9631;
wire n_8033;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_12032;
wire n_4720;
wire n_10784;
wire n_12202;
wire n_4893;
wire n_3857;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_12815;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_9945;
wire n_8661;
wire n_12431;
wire n_7424;
wire n_3714;
wire n_7523;
wire n_8654;
wire n_5039;
wire n_11855;
wire n_4772;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_3099;
wire n_11156;
wire n_8531;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6459;
wire n_6505;
wire n_12333;
wire n_12636;
wire n_8379;
wire n_8609;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_7626;
wire n_13100;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_12334;
wire n_3294;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_9209;
wire n_3686;
wire n_7669;
wire n_11218;
wire n_4502;
wire n_12119;
wire n_11787;
wire n_12618;
wire n_5958;
wire n_8793;
wire n_12355;
wire n_8103;
wire n_9767;
wire n_2971;
wire n_9838;
wire n_10195;
wire n_4277;
wire n_4526;
wire n_9300;
wire n_11500;
wire n_3490;
wire n_4849;
wire n_12943;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_8367;
wire n_11891;
wire n_7367;
wire n_5792;
wire n_11021;
wire n_3581;
wire n_12401;
wire n_8543;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_6905;
wire n_3715;
wire n_10243;
wire n_9700;
wire n_10564;
wire n_8682;
wire n_3725;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_3933;
wire n_8533;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_7244;
wire n_10745;
wire n_7368;
wire n_3691;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_7633;
wire n_4146;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_11509;
wire n_8640;
wire n_8063;
wire n_3961;
wire n_11960;
wire n_4855;
wire n_12599;
wire n_3917;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_12411;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_12465;
wire n_7427;
wire n_10605;
wire n_4004;
wire n_11029;
wire n_2967;
wire n_13250;
wire n_13118;
wire n_5404;
wire n_9933;
wire n_11449;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_4292;
wire n_9892;
wire n_8570;
wire n_6163;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_5549;
wire n_9408;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_10163;
wire n_10454;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_12568;
wire n_3280;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_12970;
wire n_8902;
wire n_8916;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_3510;
wire n_8843;
wire n_9891;
wire n_10146;
wire n_7128;
wire n_9946;
wire n_12959;
wire n_9885;
wire n_6849;
wire n_12330;
wire n_7594;
wire n_8129;
wire n_8162;
wire n_7457;
wire n_10643;
wire n_8744;
wire n_3009;
wire n_10504;
wire n_5824;
wire n_3719;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_6760;
wire n_10701;
wire n_3827;
wire n_5154;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_3889;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_12798;
wire n_5329;
wire n_9015;
wire n_9925;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_10874;
wire n_6825;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_11831;
wire n_9628;
wire n_7767;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_12243;
wire n_6611;
wire n_8562;
wire n_4560;
wire n_12614;
wire n_11378;
wire n_4899;
wire n_10250;
wire n_5728;
wire n_5471;
wire n_10032;
wire n_10592;
wire n_11433;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_7744;
wire n_7021;
wire n_2932;
wire n_3431;
wire n_10595;
wire n_7748;
wire n_8537;
wire n_3450;
wire n_6827;
wire n_10126;
wire n_12041;
wire n_4663;
wire n_11713;
wire n_11073;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_12566;
wire n_12931;
wire n_6227;
wire n_7215;
wire n_7485;
wire n_3421;
wire n_13074;
wire n_9066;
wire n_3183;
wire n_4802;
wire n_5523;
wire n_10302;
wire n_11974;
wire n_12881;
wire n_3405;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_10645;
wire n_13058;
wire n_10604;
wire n_5074;
wire n_11096;
wire n_12036;
wire n_12876;
wire n_6564;
wire n_4044;
wire n_3436;
wire n_11161;
wire n_9671;
wire n_8782;
wire n_8709;
wire n_3442;
wire n_3366;
wire n_12911;
wire n_6468;
wire n_12491;
wire n_3937;
wire n_10080;
wire n_11216;
wire n_12228;
wire n_10570;
wire n_9857;
wire n_3159;
wire n_4701;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_12929;
wire n_10882;
wire n_9338;
wire n_13071;
wire n_6857;
wire n_3240;
wire n_8144;
wire n_12261;
wire n_3576;
wire n_10435;
wire n_9542;
wire n_12536;
wire n_3385;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_12106;
wire n_12061;
wire n_3293;
wire n_3922;
wire n_11085;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_10609;
wire n_11157;
wire n_4991;
wire n_5594;
wire n_12291;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_12124;
wire n_11755;
wire n_9783;
wire n_9510;
wire n_9389;
wire n_12074;
wire n_4934;
wire n_9404;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5087;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_13234;
wire n_5292;
wire n_9314;
wire n_11918;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5000;
wire n_5403;
wire n_12887;
wire n_5551;
wire n_7652;
wire n_3150;
wire n_10220;
wire n_8701;
wire n_10341;
wire n_11347;
wire n_4479;
wire n_6499;
wire n_10550;
wire n_7830;
wire n_4011;
wire n_5131;
wire n_12217;
wire n_12365;
wire n_3133;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_9679;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_13272;
wire n_4688;
wire n_4753;
wire n_8712;
wire n_10232;
wire n_4058;
wire n_10461;
wire n_8289;
wire n_11178;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_7966;
wire n_8591;
wire n_5059;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_8824;
wire n_11673;
wire n_11432;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_10412;
wire n_4475;
wire n_5242;
wire n_10326;
wire n_12650;
wire n_5219;
wire n_8417;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_3537;
wire n_10499;
wire n_8340;
wire n_4443;
wire n_6008;
wire n_3887;
wire n_12487;
wire n_12658;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_5460;
wire n_4587;
wire n_4114;
wire n_2948;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_9210;
wire n_12185;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_6893;
wire n_5686;
wire n_5899;
wire n_7406;
wire n_8681;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_3223;
wire n_10617;
wire n_12271;
wire n_12704;
wire n_3140;
wire n_7807;
wire n_4749;
wire n_3185;
wire n_9592;
wire n_5155;
wire n_7680;
wire n_9180;
wire n_10922;
wire n_10544;
wire n_12958;
wire n_13030;
wire n_3654;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_12056;
wire n_8106;
wire n_9502;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_3788;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_6422;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_3837;
wire n_11087;
wire n_11477;
wire n_3325;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_4085;
wire n_13243;
wire n_4464;
wire n_8612;
wire n_13042;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_10095;
wire n_4659;
wire n_10309;
wire n_3600;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_3324;
wire n_6160;
wire n_9871;
wire n_10050;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_7066;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_7789;
wire n_13197;
wire n_10306;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_7193;
wire n_3987;
wire n_6039;
wire n_4487;
wire n_11919;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_10450;
wire n_5721;
wire n_11414;
wire n_11472;
wire n_3638;
wire n_9114;
wire n_11978;
wire n_4816;
wire n_12520;
wire n_8515;
wire n_10529;
wire n_5719;
wire n_5773;
wire n_5482;
wire n_3393;
wire n_8812;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_3451;
wire n_9392;
wire n_13148;
wire n_10429;
wire n_4937;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_3615;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_11538;
wire n_3072;
wire n_3087;
wire n_10037;
wire n_12808;
wire n_4222;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_4401;
wire n_12744;
wire n_6064;
wire n_11136;
wire n_9903;
wire n_3142;
wire n_4015;
wire n_5793;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_4709;
wire n_9228;
wire n_10179;
wire n_11539;
wire n_4976;
wire n_7710;
wire n_12143;
wire n_9499;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_9522;
wire n_5578;
wire n_11215;
wire n_4658;
wire n_5296;
wire n_11076;
wire n_9366;
wire n_11890;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_9148;
wire n_11054;
wire n_11806;
wire n_8406;
wire n_6277;
wire n_10754;
wire n_5742;
wire n_5207;
wire n_11050;
wire n_3705;
wire n_3211;
wire n_12443;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_11683;
wire n_8554;
wire n_10920;
wire n_9275;
wire n_10223;
wire n_6051;
wire n_8896;
wire n_4665;
wire n_3582;
wire n_11484;
wire n_7206;
wire n_4223;
wire n_11126;
wire n_7538;
wire n_5674;
wire n_12934;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_5282;
wire n_10295;
wire n_9409;
wire n_5464;
wire n_6799;
wire n_10336;
wire n_10228;
wire n_12555;
wire n_4362;
wire n_3913;
wire n_3311;
wire n_7716;
wire n_6487;
wire n_11646;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_8818;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_4348;
wire n_12980;
wire n_9881;
wire n_12530;
wire n_5013;
wire n_8954;
wire n_6807;
wire n_9463;
wire n_7251;
wire n_4489;
wire n_4839;
wire n_7254;
wire n_12212;
wire n_10466;
wire n_12973;
wire n_3163;
wire n_7540;
wire n_11953;
wire n_4404;
wire n_13123;
wire n_5589;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_13231;
wire n_12624;
wire n_7882;
wire n_8552;
wire n_10425;
wire n_7554;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_8373;
wire n_10848;
wire n_13165;
wire n_6481;
wire n_5628;
wire n_4825;
wire n_7765;
wire n_11482;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_12151;
wire n_4006;
wire n_11089;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_6384;
wire n_3869;
wire n_7421;
wire n_10166;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_13179;
wire n_5251;
wire n_3753;
wire n_12033;
wire n_11839;
wire n_3742;
wire n_9844;
wire n_3683;
wire n_8318;
wire n_4801;
wire n_12826;
wire n_3260;
wire n_10366;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_11365;
wire n_3175;
wire n_9595;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_11217;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_9287;
wire n_7991;
wire n_13051;
wire n_6233;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_3284;
wire n_12214;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_8926;
wire n_6257;
wire n_4386;
wire n_4132;
wire n_10361;
wire n_11228;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_4955;
wire n_8965;
wire n_11290;
wire n_5936;
wire n_4149;
wire n_12518;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_3234;
wire n_9052;
wire n_8817;
wire n_8190;
wire n_11488;
wire n_12162;
wire n_3202;
wire n_3220;
wire n_6587;
wire n_6987;
wire n_7781;
wire n_7360;
wire n_11037;
wire n_11702;
wire n_6069;
wire n_7497;
wire n_4655;
wire n_11372;
wire n_5706;
wire n_7665;
wire n_9354;
wire n_3429;
wire n_10501;
wire n_10817;
wire n_11829;
wire n_11517;
wire n_7793;
wire n_8355;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_12741;
wire n_7101;
wire n_7671;
wire n_9436;
wire n_7530;
wire n_8489;
wire n_13150;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_11551;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_7654;
wire n_13152;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_8369;
wire n_9022;
wire n_9238;
wire n_8059;
wire n_6633;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_6579;
wire n_11665;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_11138;
wire n_11731;
wire n_5187;
wire n_5875;
wire n_9839;
wire n_12821;
wire n_4024;
wire n_8831;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_7120;
wire n_8728;
wire n_10807;
wire n_12478;
wire n_12233;
wire n_3250;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_8853;
wire n_4582;
wire n_6252;
wire n_4860;
wire n_6211;
wire n_10511;
wire n_5844;
wire n_8862;
wire n_3414;
wire n_10580;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_9675;
wire n_7786;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_10058;
wire n_10873;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_11454;
wire n_3449;
wire n_8900;
wire n_12523;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_10484;
wire n_4304;
wire n_4558;
wire n_6737;
wire n_11744;
wire n_4488;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_8478;
wire n_6606;
wire n_6695;
wire n_3550;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_4211;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_11626;
wire n_12148;
wire n_4016;
wire n_11072;
wire n_5867;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_12907;
wire n_3839;
wire n_8497;
wire n_10770;
wire n_8820;
wire n_6410;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_5597;
wire n_9028;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_9374;
wire n_7419;
wire n_6506;
wire n_5515;
wire n_5662;
wire n_3131;
wire n_12132;
wire n_3730;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_10593;
wire n_13019;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_4397;
wire n_3399;
wire n_12182;
wire n_12670;
wire n_5050;
wire n_10636;
wire n_12043;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_10203;
wire n_3498;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_8992;
wire n_12708;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_6234;
wire n_2957;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_9983;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_6608;
wire n_10467;
wire n_3533;
wire n_9109;
wire n_9849;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_11207;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_12493;
wire n_3138;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_9237;
wire n_11668;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_8466;
wire n_6753;
wire n_12137;
wire n_6527;
wire n_7341;
wire n_11328;
wire n_2988;
wire n_9349;
wire n_12306;
wire n_4908;
wire n_3136;
wire n_11200;
wire n_12088;
wire n_11091;
wire n_8094;
wire n_4109;
wire n_4192;
wire n_10940;
wire n_6639;
wire n_4824;
wire n_12096;
wire n_4567;
wire n_6430;
wire n_12508;
wire n_5150;
wire n_8832;
wire n_10987;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_4595;
wire n_4174;
wire n_12891;
wire n_11098;
wire n_11615;
wire n_10533;
wire n_11059;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_11965;
wire n_4904;
wire n_10938;
wire n_10176;
wire n_7517;
wire n_6627;
wire n_8080;
wire n_3544;
wire n_5988;
wire n_4150;
wire n_5585;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_7745;
wire n_12941;
wire n_3105;
wire n_6666;
wire n_3692;
wire n_10927;
wire n_12200;
wire n_4616;
wire n_8321;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_4982;
wire n_11722;
wire n_8786;
wire n_8592;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_4643;
wire n_6249;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_9805;
wire n_5480;
wire n_10155;
wire n_4323;
wire n_8157;
wire n_4831;
wire n_7095;
wire n_3045;
wire n_3821;
wire n_11461;
wire n_10714;
wire n_11701;
wire n_6969;
wire n_6615;
wire n_6161;
wire n_7459;
wire n_2970;
wire n_7294;
wire n_8206;
wire n_3676;
wire n_4896;
wire n_3666;
wire n_4916;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_9110;
wire n_11811;
wire n_10569;
wire n_8622;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_9335;
wire n_6062;
wire n_7908;
wire n_12550;
wire n_4122;
wire n_9452;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_10051;
wire n_4209;
wire n_8104;
wire n_10414;
wire n_11255;
wire n_8344;
wire n_3858;
wire n_5284;
wire n_11720;
wire n_4298;
wire n_12673;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_4128;
wire n_10746;
wire n_12225;
wire n_9188;
wire n_6294;
wire n_5147;
wire n_9611;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_8779;
wire n_9810;
wire n_8621;
wire n_5503;
wire n_5845;
wire n_9250;
wire n_5945;
wire n_9550;
wire n_11212;
wire n_12884;
wire n_13145;
wire n_10697;
wire n_11714;
wire n_11263;
wire n_10641;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_12207;
wire n_9975;
wire n_7250;
wire n_5600;
wire n_5755;
wire n_8762;
wire n_12011;
wire n_13195;
wire n_8043;
wire n_8694;
wire n_5048;
wire n_6053;
wire n_11994;
wire n_7252;
wire n_3246;
wire n_3381;
wire n_9207;
wire n_3208;
wire n_4944;
wire n_11860;
wire n_11990;
wire n_12837;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_10926;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_10626;
wire n_6901;
wire n_4935;
wire n_13273;
wire n_4694;
wire n_11503;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_2962;
wire n_8376;
wire n_8171;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_6774;
wire n_12854;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_8710;
wire n_12806;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_8599;
wire n_2960;
wire n_8549;
wire n_10172;
wire n_5993;
wire n_8054;
wire n_11273;
wire n_10400;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_3258;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_13218;
wire n_9096;
wire n_9081;
wire n_11697;
wire n_13076;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_9236;
wire n_11762;
wire n_11969;
wire n_12950;
wire n_7914;
wire n_8628;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_13028;
wire n_8857;
wire n_8517;
wire n_4850;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_3008;
wire n_6162;
wire n_10433;
wire n_6779;
wire n_8010;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_9116;
wire n_10774;
wire n_3972;
wire n_12332;
wire n_4153;
wire n_11034;
wire n_10901;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_3506;
wire n_7216;
wire n_3855;
wire n_12762;
wire n_11499;
wire n_10825;
wire n_3091;
wire n_4317;
wire n_8275;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_10761;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_9035;
wire n_11579;
wire n_10398;
wire n_8291;
wire n_4143;
wire n_4170;
wire n_11535;
wire n_3642;
wire n_12558;
wire n_4650;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_5016;
wire n_12975;
wire n_11402;
wire n_6458;
wire n_7642;
wire n_4967;
wire n_9678;
wire n_11401;
wire n_8247;
wire n_6577;
wire n_12506;
wire n_6740;
wire n_3308;
wire n_12718;
wire n_12956;
wire n_11510;
wire n_6315;
wire n_10581;
wire n_12638;
wire n_4912;
wire n_4799;
wire n_9284;
wire n_12736;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_12086;
wire n_5170;
wire n_6910;
wire n_7604;
wire n_6262;
wire n_7703;
wire n_3515;
wire n_9606;
wire n_6319;
wire n_2951;
wire n_10470;
wire n_11589;
wire n_2949;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_12350;
wire n_12542;
wire n_5028;
wire n_5839;
wire n_6536;
wire n_12747;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_8827;
wire n_10625;
wire n_8280;
wire n_12561;
wire n_12390;
wire n_5514;
wire n_13216;
wire n_2931;
wire n_8388;
wire n_12849;
wire n_10235;
wire n_11312;
wire n_3866;
wire n_6978;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_4543;
wire n_10445;
wire n_7378;
wire n_10738;
wire n_12866;
wire n_4157;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_9190;
wire n_6947;
wire n_11612;
wire n_4229;
wire n_9482;
wire n_5293;
wire n_12447;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_12900;
wire n_3865;
wire n_4073;
wire n_8569;
wire n_3629;
wire n_5400;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_8877;
wire n_9412;
wire n_7498;
wire n_10679;
wire n_11323;
wire n_10799;
wire n_3846;
wire n_6321;
wire n_12914;
wire n_11916;
wire n_3512;
wire n_6819;
wire n_7501;
wire n_5201;
wire n_9506;
wire n_10136;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_10585;
wire n_12764;
wire n_4783;
wire n_11356;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_9092;
wire n_10034;
wire n_9451;
wire n_4910;
wire n_11148;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_3083;
wire n_6899;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_6592;
wire n_11280;
wire n_12337;
wire n_13254;
wire n_3049;
wire n_8686;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_7613;
wire n_3541;
wire n_11493;
wire n_6101;
wire n_9220;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_10528;
wire n_10860;
wire n_12763;
wire n_4930;
wire n_8588;
wire n_11339;
wire n_5623;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_4112;
wire n_12712;
wire n_11220;
wire n_9012;
wire n_4557;
wire n_13012;
wire n_4917;
wire n_8698;
wire n_8924;
wire n_12584;
wire n_4432;
wire n_3739;
wire n_10376;
wire n_12752;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_4593;
wire n_7238;
wire n_9994;
wire n_4465;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_11596;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_11885;
wire n_5117;
wire n_5663;
wire n_7572;
wire n_3363;
wire n_8214;
wire n_10224;
wire n_11955;
wire n_12777;
wire n_5990;
wire n_7043;
wire n_10777;
wire n_3721;
wire n_11462;
wire n_3062;
wire n_11732;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_12819;
wire n_8722;
wire n_11654;
wire n_12268;
wire n_10214;
wire n_8241;
wire n_8589;
wire n_12077;
wire n_3969;
wire n_12982;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_4231;
wire n_6281;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_13133;
wire n_4256;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_6311;
wire n_10469;
wire n_9229;
wire n_11194;
wire n_11480;
wire n_7590;
wire n_9342;
wire n_12237;
wire n_13271;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_5426;
wire n_10175;
wire n_5803;
wire n_11481;
wire n_9868;
wire n_11375;
wire n_5285;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_4335;
wire n_9311;
wire n_12275;
wire n_6593;
wire n_8630;
wire n_12376;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_4521;
wire n_8405;
wire n_8145;
wire n_10447;
wire n_9260;
wire n_7176;
wire n_8928;
wire n_7682;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_11925;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_10406;
wire n_3204;
wire n_5715;
wire n_12509;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_11985;
wire n_8447;
wire n_7901;
wire n_5395;
wire n_10522;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_11782;
wire n_6446;
wire n_10278;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_3802;
wire n_3256;
wire n_6996;
wire n_7218;
wire n_8828;
wire n_9430;
wire n_11407;
wire n_9750;
wire n_9749;
wire n_12710;
wire n_6749;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_7005;
wire n_10408;
wire n_8572;
wire n_10965;
wire n_10798;
wire n_7732;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_9776;
wire n_11911;
wire n_6777;
wire n_4265;
wire n_11987;
wire n_11442;
wire n_8227;
wire n_12936;
wire n_12721;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_8475;
wire n_3060;
wire n_11730;
wire n_10482;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_4105;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_12039;
wire n_4926;
wire n_11388;
wire n_11651;
wire n_3123;
wire n_8314;
wire n_3380;
wire n_9386;
wire n_10154;
wire n_5617;
wire n_7922;
wire n_13089;
wire n_10377;
wire n_5580;
wire n_5266;
wire n_4828;
wire n_10033;
wire n_9926;
wire n_3038;
wire n_11121;
wire n_13167;
wire n_11270;
wire n_12329;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_8311;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_3769;
wire n_12253;
wire n_11147;
wire n_12928;
wire n_5310;
wire n_9661;
wire n_9843;
wire n_9877;
wire n_8764;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_13001;
wire n_5390;
wire n_13232;
wire n_9901;
wire n_5593;
wire n_12990;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_8567;
wire n_11817;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_5237;
wire n_3344;
wire n_5133;
wire n_11042;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_3989;
wire n_7144;
wire n_7089;
wire n_7286;
wire n_11479;
wire n_11737;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_12028;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_13016;
wire n_11272;
wire n_13095;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_6332;
wire n_4303;
wire n_5853;
wire n_12048;
wire n_8283;
wire n_5982;
wire n_10930;
wire n_11600;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_3147;
wire n_4909;
wire n_12057;
wire n_6696;
wire n_3925;
wire n_13251;
wire n_9882;
wire n_9527;
wire n_3180;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_3472;
wire n_8516;
wire n_8302;
wire n_10637;
wire n_8317;
wire n_5376;
wire n_12229;
wire n_5106;
wire n_6116;
wire n_9205;
wire n_9511;
wire n_8167;
wire n_7859;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_7972;
wire n_11254;
wire n_4768;
wire n_11617;
wire n_9071;
wire n_7916;
wire n_3717;
wire n_9368;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_10415;
wire n_13069;
wire n_11711;
wire n_5410;
wire n_12362;
wire n_8944;
wire n_6167;
wire n_13233;
wire n_11931;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_8109;
wire n_9459;
wire n_5156;
wire n_12780;
wire n_13267;
wire n_6307;
wire n_10410;
wire n_6094;
wire n_9098;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_9133;
wire n_12664;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_9504;
wire n_8975;
wire n_6267;
wire n_9063;
wire n_7787;
wire n_3903;
wire n_12360;
wire n_5998;
wire n_9268;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_10456;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_13186;
wire n_5916;
wire n_11907;
wire n_4648;
wire n_10096;
wire n_3094;
wire n_10025;
wire n_10627;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_6299;
wire n_6813;
wire n_8825;
wire n_12969;
wire n_11753;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_8266;
wire n_5691;
wire n_12457;
wire n_4951;
wire n_8981;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_3079;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_12939;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_10404;
wire n_8639;
wire n_8138;
wire n_8058;
wire n_9308;
wire n_3504;
wire n_6638;
wire n_12779;
wire n_11838;
wire n_10508;
wire n_7719;
wire n_4272;
wire n_10811;
wire n_8333;
wire n_2930;
wire n_5615;
wire n_6220;
wire n_7562;
wire n_3111;
wire n_12816;
wire n_6985;
wire n_7619;
wire n_12783;
wire n_7170;
wire n_9211;
wire n_12019;
wire n_8176;
wire n_8124;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_10891;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_3054;
wire n_10803;
wire n_8147;
wire n_13190;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_5262;
wire n_10700;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_11695;
wire n_4620;
wire n_3152;
wire n_7935;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_8458;
wire n_6772;
wire n_8113;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_3178;
wire n_11453;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_6318;
wire n_11970;
wire n_4099;
wire n_7918;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_6916;
wire n_4490;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_10783;
wire n_11862;
wire n_10147;
wire n_12163;
wire n_10725;
wire n_3952;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_12944;
wire n_3911;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_11660;
wire n_4285;
wire n_3465;
wire n_10812;
wire n_12297;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_6604;
wire n_5161;
wire n_5373;
wire n_10001;
wire n_3708;
wire n_11107;
wire n_4078;
wire n_9301;
wire n_12145;
wire n_3046;
wire n_11088;
wire n_2956;
wire n_5573;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_8160;
wire n_10284;
wire n_12757;
wire n_12054;
wire n_5659;
wire n_8099;
wire n_11595;
wire n_8840;
wire n_3619;
wire n_11405;
wire n_13189;
wire n_5881;
wire n_8522;
wire n_12971;
wire n_7222;
wire n_7942;
wire n_8578;
wire n_6473;
wire n_13103;
wire n_4198;
wire n_3754;
wire n_10046;
wire n_12328;
wire n_11318;
wire n_9083;
wire n_7725;
wire n_10977;
wire n_2974;
wire n_4213;
wire n_11299;
wire n_10397;
wire n_2982;
wire n_6483;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_4065;
wire n_5863;
wire n_7647;
wire n_8626;
wire n_10385;
wire n_10936;
wire n_12442;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_9835;
wire n_7300;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_4446;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_4733;
wire n_6729;
wire n_6728;
wire n_4764;
wire n_3879;
wire n_11240;
wire n_4743;
wire n_10207;
wire n_3080;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_11487;
wire n_8441;
wire n_11441;
wire n_6076;
wire n_8933;
wire n_3023;
wire n_3232;
wire n_7778;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_11287;
wire n_4060;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_4879;
wire n_6390;
wire n_10139;
wire n_13246;
wire n_5796;
wire n_10104;
wire n_8726;
wire n_12986;
wire n_11381;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_9117;
wire n_9720;
wire n_3028;
wire n_7746;
wire n_3662;
wire n_9381;
wire n_2981;
wire n_6958;
wire n_3076;
wire n_10169;
wire n_12049;
wire n_12690;
wire n_7563;
wire n_12475;
wire n_3624;
wire n_4556;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_8414;
wire n_6297;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_12526;
wire n_4687;
wire n_7531;
wire n_12377;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_13214;
wire n_8615;
wire n_11062;
wire n_7721;
wire n_7192;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_9887;
wire n_9149;
wire n_4600;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_13211;
wire n_8316;
wire n_4250;
wire n_9990;
wire n_5829;
wire n_3906;
wire n_10005;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_4954;
wire n_5191;
wire n_8505;
wire n_9273;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_13061;
wire n_9682;
wire n_4881;
wire n_12513;
wire n_4253;
wire n_10640;
wire n_6582;
wire n_5734;
wire n_4255;
wire n_4071;
wire n_10729;
wire n_12545;
wire n_7388;
wire n_3568;
wire n_3850;
wire n_11657;
wire n_9924;
wire n_8717;
wire n_5770;
wire n_5705;
wire n_3313;
wire n_13176;
wire n_4605;
wire n_9064;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_13102;
wire n_11268;
wire n_12753;
wire n_4691;
wire n_7090;
wire n_9254;
wire n_12894;
wire n_3943;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_4305;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_4297;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_12010;
wire n_9738;
wire n_5675;
wire n_9570;
wire n_12026;
wire n_4227;
wire n_12356;
wire n_11857;
wire n_11077;
wire n_6240;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_9593;
wire n_7689;
wire n_9846;
wire n_13262;
wire n_6511;
wire n_5297;
wire n_7121;
wire n_9469;
wire n_10764;
wire n_9677;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_8449;
wire n_6358;
wire n_13204;
wire n_4094;
wire n_6603;
wire n_4765;
wire n_3193;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_6986;
wire n_4732;
wire n_3912;
wire n_8801;
wire n_9322;
wire n_3118;
wire n_10438;
wire n_5959;
wire n_11201;
wire n_3720;
wire n_10531;
wire n_8918;
wire n_8031;
wire n_12878;
wire n_9348;
wire n_12188;
wire n_8219;
wire n_8696;
wire n_4745;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_12630;
wire n_4581;
wire n_6890;
wire n_11028;
wire n_12171;
wire n_4377;
wire n_12299;
wire n_12022;
wire n_9249;
wire n_12935;
wire n_7827;
wire n_8180;
wire n_10741;
wire n_6109;
wire n_10760;
wire n_4792;
wire n_12425;
wire n_9444;
wire n_7731;
wire n_3842;
wire n_10772;
wire n_11527;
wire n_7114;
wire n_4878;
wire n_3514;
wire n_11327;
wire n_10915;
wire n_4979;
wire n_9535;
wire n_6770;
wire n_3036;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_5302;
wire n_12000;
wire n_4511;
wire n_9707;
wire n_12490;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_3895;
wire n_8943;
wire n_8486;
wire n_10279;
wire n_4520;
wire n_5299;
wire n_12829;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_10680;
wire n_10127;
wire n_3599;
wire n_5543;
wire n_5361;
wire n_11610;
wire n_7132;
wire n_7081;
wire n_11814;
wire n_12255;
wire n_12739;
wire n_13015;
wire n_5885;
wire n_6663;
wire n_4199;
wire n_9723;
wire n_5356;
wire n_12609;
wire n_4441;
wire n_7319;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_11176;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_11360;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5038;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_10039;
wire n_11726;
wire n_10854;
wire n_11358;
wire n_5463;
wire n_3022;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_12904;
wire n_8833;
wire n_9191;
wire n_5489;
wire n_5892;
wire n_7828;
wire n_10142;
wire n_4773;
wire n_7940;
wire n_9918;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_6009;
wire n_3281;
wire n_9034;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_9390;
wire n_5113;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_5714;
wire n_3549;
wire n_8541;
wire n_8074;
wire n_8485;
wire n_8860;
wire n_5510;
wire n_3940;
wire n_6621;
wire n_11958;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_13070;
wire n_8271;
wire n_5692;
wire n_8473;
wire n_4800;
wire n_9266;
wire n_3453;
wire n_12728;
wire n_5555;
wire n_3410;
wire n_10027;
wire n_12784;
wire n_3768;
wire n_4958;
wire n_4043;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_8699;
wire n_3785;
wire n_6897;
wire n_2963;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_5366;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_2980;
wire n_4886;
wire n_9931;
wire n_13198;
wire n_3227;
wire n_3289;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_4055;
wire n_12610;
wire n_11671;
wire n_10328;
wire n_5968;
wire n_11251;
wire n_12293;
wire n_11063;
wire n_3326;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_13174;
wire n_4200;
wire n_3460;
wire n_7108;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_8368;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_11879;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_8546;
wire n_10963;
wire n_8300;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_8148;
wire n_11400;
wire n_8150;
wire n_3578;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_10483;
wire n_12160;
wire n_4737;
wire n_11563;
wire n_4925;
wire n_9620;
wire n_4116;
wire n_5415;
wire n_8986;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_5419;
wire n_11243;
wire n_3805;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_6409;
wire n_11939;
wire n_3252;
wire n_3253;
wire n_7954;
wire n_9824;
wire n_11119;
wire n_7951;
wire n_7552;
wire n_8096;
wire n_11468;
wire n_12166;
wire n_8233;
wire n_6130;
wire n_4603;
wire n_7273;
wire n_9683;
wire n_10646;
wire n_7231;
wire n_5080;
wire n_5976;
wire n_11704;
wire n_3128;
wire n_5732;
wire n_5372;
wire n_11878;
wire n_4471;
wire n_7772;
wire n_7449;
wire n_8763;
wire n_12800;
wire n_5208;
wire n_8679;
wire n_7239;
wire n_9848;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_6623;
wire n_9561;
wire n_10378;
wire n_12070;
wire n_9714;
wire n_9740;
wire n_3078;
wire n_9773;
wire n_10313;
wire n_3838;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_3941;
wire n_3793;
wire n_10216;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_12354;
wire n_12666;
wire n_6047;
wire n_12581;
wire n_8292;
wire n_12631;
wire n_3037;
wire n_10133;
wire n_3729;
wire n_8601;
wire n_10773;
wire n_4994;
wire n_6652;
wire n_9377;
wire n_11932;
wire n_10971;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_6921;
wire n_6970;
wire n_5168;
wire n_4661;
wire n_13027;
wire n_12867;
wire n_4988;
wire n_7674;
wire n_9826;
wire n_3171;
wire n_12607;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_12075;
wire n_4540;
wire n_11942;
wire n_6344;
wire n_12305;
wire n_12123;
wire n_3459;
wire n_9772;
wire n_12170;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_6624;
wire n_9630;
wire n_6956;
wire n_4284;
wire n_12966;
wire n_6305;
wire n_9255;
wire n_6209;
wire n_8310;
wire n_10231;
wire n_12547;
wire n_9758;
wire n_3426;
wire n_11922;
wire n_4971;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_5125;
wire n_5857;
wire n_12358;
wire n_7329;
wire n_8646;
wire n_7408;
wire n_9691;
wire n_12997;
wire n_10259;
wire n_7107;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_7690;
wire n_8969;
wire n_7123;
wire n_10752;
wire n_11577;
wire n_5499;
wire n_8117;
wire n_10067;
wire n_3229;
wire n_3348;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_12498;
wire n_11475;
wire n_6950;
wire n_8208;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_11010;
wire n_2933;
wire n_10274;
wire n_9590;
wire n_11588;
wire n_6694;
wire n_3497;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_9168;
wire n_3580;
wire n_11221;
wire n_12387;
wire n_9497;
wire n_8536;
wire n_13255;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_3704;
wire n_11448;
wire n_9219;
wire n_5507;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_8914;
wire n_12576;
wire n_7258;
wire n_5190;
wire n_8391;
wire n_10579;
wire n_10832;
wire n_3173;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_6466;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_10584;
wire n_4218;
wire n_5392;
wire n_12862;
wire n_11445;
wire n_13151;
wire n_3880;
wire n_3685;
wire n_8216;
wire n_11552;
wire n_10332;
wire n_7709;
wire n_11874;
wire n_3609;
wire n_9982;
wire n_10171;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_12656;
wire n_9852;
wire n_6820;
wire n_11623;
wire n_8313;
wire n_3019;
wire n_3471;
wire n_5511;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_4175;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_10540;
wire n_11936;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_3200;
wire n_4771;
wire n_10200;
wire n_7332;
wire n_12734;
wire n_3259;
wire n_10382;
wire n_13164;
wire n_3167;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_3867;
wire n_10269;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_12262;
wire n_13223;
wire n_9169;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_4140;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_7766;
wire n_11018;
wire n_8738;
wire n_10981;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_12797;
wire n_3032;
wire n_6223;
wire n_11376;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_9481;
wire n_9600;
wire n_9122;
wire n_8085;
wire n_11274;
wire n_5098;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_5707;
wire n_12012;
wire n_5140;
wire n_4992;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_9927;
wire n_5497;
wire n_10076;
wire n_11515;
wire n_8721;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_11554;
wire n_7637;
wire n_10148;
wire n_10318;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_7127;
wire n_4533;
wire n_9635;
wire n_5481;
wire n_12890;
wire n_3590;
wire n_8666;
wire n_5344;
wire n_9264;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_5408;
wire n_7801;
wire n_9155;
wire n_4053;
wire n_10234;
wire n_8460;
wire n_3848;
wire n_10416;
wire n_3327;
wire n_8836;
wire n_7959;
wire n_7019;
wire n_8181;
wire n_11325;
wire n_8254;
wire n_4167;
wire n_8071;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_10731;
wire n_10735;
wire n_10583;
wire n_9878;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_9825;
wire n_5494;
wire n_7444;
wire n_11628;
wire n_5234;
wire n_4431;
wire n_7546;
wire n_6272;
wire n_4387;
wire n_6588;
wire n_3265;
wire n_11549;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_12286;
wire n_9001;
wire n_10393;
wire n_11498;
wire n_13081;
wire n_10513;
wire n_12252;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_12627;
wire n_4890;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_12281;
wire n_11237;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_9373;
wire n_6268;
wire n_5827;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_12347;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_11181;
wire n_9967;
wire n_7521;
wire n_3407;
wire n_5992;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_3856;
wire n_4236;
wire n_9971;
wire n_7187;
wire n_3425;
wire n_10894;
wire n_3894;
wire n_9524;
wire n_12277;
wire n_3127;
wire n_12698;
wire n_5312;
wire n_3623;
wire n_6467;
wire n_9182;
wire n_9243;
wire n_9282;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_9224;
wire n_3646;
wire n_10347;
wire n_5513;
wire n_5614;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_12410;
wire n_4830;
wire n_4706;
wire n_13225;
wire n_5225;
wire n_4570;
wire n_10208;
wire n_7722;
wire n_3188;
wire n_3243;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_8141;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_12957;
wire n_4693;
wire n_13141;
wire n_4206;
wire n_11616;
wire n_8791;
wire n_11920;
wire n_10793;
wire n_8288;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_12786;
wire n_5049;
wire n_12711;
wire n_11675;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_5846;
wire n_8323;
wire n_10440;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_10391;
wire n_7636;
wire n_9799;
wire n_9695;
wire n_2955;
wire n_11083;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_7866;
wire n_4609;
wire n_11306;
wire n_3051;
wire n_9784;
wire n_11198;
wire n_3367;
wire n_7205;
wire n_8757;
wire n_7990;
wire n_7020;
wire n_10036;
wire n_13035;
wire n_13021;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_8596;
wire n_3525;
wire n_5157;
wire n_3314;
wire n_11840;
wire n_2993;
wire n_4754;
wire n_3016;
wire n_4647;
wire n_9556;
wire n_3688;
wire n_11292;
wire n_8720;
wire n_8590;
wire n_10261;
wire n_13157;
wire n_5708;
wire n_4003;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_4894;
wire n_5474;
wire n_12289;
wire n_4113;
wire n_10813;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_11326;
wire n_13046;
wire n_6421;
wire n_11870;
wire n_7407;
wire n_9827;
wire n_3466;
wire n_10907;
wire n_5704;
wire n_11431;
wire n_4983;
wire n_7148;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_6236;
wire n_9417;
wire n_11834;
wire n_12020;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_3907;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_3338;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_6835;
wire n_8834;
wire n_3636;
wire n_11624;
wire n_8826;
wire n_11352;
wire n_5516;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_10822;
wire n_11234;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_12099;
wire n_12858;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_7799;
wire n_8364;
wire n_5698;
wire n_11092;
wire n_3276;
wire n_9534;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_3572;
wire n_11836;
wire n_6602;
wire n_10924;
wire n_3886;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_9647;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_10885;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_13201;
wire n_3637;
wire n_6242;
wire n_12527;
wire n_4574;
wire n_13274;
wire n_12379;
wire n_9312;
wire n_9019;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_4234;
wire n_12477;
wire n_7469;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_10895;
wire n_3974;
wire n_10875;
wire n_3634;
wire n_11736;
wire n_11977;
wire n_7560;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_3236;
wire n_11696;
wire n_12400;
wire n_5096;
wire n_3141;
wire n_11734;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_12114;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_11507;
wire n_9145;
wire n_7082;
wire n_12092;
wire n_3112;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_4270;
wire n_11837;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_3417;
wire n_9000;
wire n_5677;
wire n_9454;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_8307;
wire n_5153;
wire n_11967;
wire n_9383;
wire n_9253;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_5927;
wire n_7392;
wire n_7495;
wire n_9566;
wire n_11338;
wire n_11996;
wire n_5435;
wire n_12174;
wire n_9765;
wire n_3213;
wire n_9807;
wire n_4333;
wire n_5200;
wire n_3820;
wire n_8706;
wire n_9057;
wire n_6400;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_6941;
wire n_5115;
wire n_12053;
wire n_5566;
wire n_11250;
wire n_7829;
wire n_12619;
wire n_3249;
wire n_7543;
wire n_8680;
wire n_11289;
wire n_13169;
wire n_7877;
wire n_7963;
wire n_9672;
wire n_12582;
wire n_4152;
wire n_5487;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_5486;
wire n_9503;
wire n_12423;
wire n_11391;
wire n_5092;
wire n_5244;
wire n_3172;
wire n_13265;
wire n_8270;
wire n_4832;
wire n_12714;
wire n_5889;
wire n_11738;
wire n_3217;
wire n_7284;
wire n_12153;
wire n_7264;
wire n_5391;
wire n_11522;
wire n_9763;
wire n_7737;
wire n_6537;
wire n_8614;
wire n_7328;
wire n_10702;
wire n_11070;
wire n_10958;
wire n_9479;
wire n_3394;
wire n_9162;
wire n_9568;
wire n_3536;
wire n_12405;
wire n_8816;
wire n_3957;
wire n_3710;
wire n_9119;
wire n_4195;
wire n_10319;
wire n_5849;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_6224;
wire n_6578;
wire n_3040;
wire n_8802;
wire n_9859;
wire n_3279;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_6092;
wire n_10879;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_10639;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_8121;
wire n_3905;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_12554;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_10491;
wire n_12037;
wire n_5152;
wire n_5265;
wire n_12792;
wire n_11717;
wire n_9943;
wire n_4927;
wire n_5574;
wire n_12391;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_7152;
wire n_11723;
wire n_9575;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_11830;
wire n_12438;
wire n_5469;
wire n_8766;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_12838;
wire n_6567;
wire n_9165;
wire n_12323;
wire n_5910;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_3134;
wire n_5965;
wire n_9596;
wire n_3115;
wire n_7240;
wire n_7570;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_10476;
wire n_4875;
wire n_9966;
wire n_13156;
wire n_7817;
wire n_5682;
wire n_10710;
wire n_5387;
wire n_5557;
wire n_11394;
wire n_8850;
wire n_11906;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_8002;
wire n_9741;
wire n_3307;
wire n_11486;
wire n_12677;
wire n_4321;
wire n_10180;
wire n_4183;
wire n_8370;
wire n_7237;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_9090;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_4145;
wire n_4901;
wire n_4821;
wire n_3121;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_12901;
wire n_4040;
wire n_10518;
wire n_8301;
wire n_12895;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_9771;
wire n_5316;
wire n_7718;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_7396;
wire n_10942;
wire n_12726;
wire n_12668;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_13010;
wire n_6320;
wire n_8126;
wire n_11239;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4943;
wire n_10953;
wire n_12432;
wire n_3044;
wire n_4757;
wire n_7561;
wire n_6810;
wire n_7842;
wire n_12352;
wire n_6202;
wire n_10099;
wire n_9969;
wire n_11437;
wire n_4682;
wire n_9961;
wire n_12898;
wire n_12879;
wire n_5564;
wire n_11869;
wire n_12559;
wire n_5620;
wire n_7163;
wire n_4530;
wire n_10343;
wire n_10836;
wire n_4942;
wire n_9899;
wire n_9258;
wire n_13004;
wire n_10181;
wire n_10286;
wire n_5406;
wire n_8072;
wire n_10371;
wire n_8277;
wire n_7236;
wire n_4604;
wire n_13117;
wire n_10257;
wire n_3305;
wire n_7130;
wire n_2992;
wire n_5724;
wire n_7201;
wire n_11219;
wire n_3157;
wire n_4841;
wire n_10047;
wire n_3221;
wire n_3267;
wire n_5806;
wire n_10949;
wire n_4338;
wire n_3457;
wire n_10486;
wire n_11226;
wire n_11282;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_3005;
wire n_11413;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_5355;
wire n_5320;
wire n_3984;
wire n_7491;
wire n_5353;
wire n_9995;
wire n_5186;
wire n_5710;
wire n_9076;
wire n_11232;
wire n_12351;
wire n_12693;
wire n_9105;
wire n_6792;
wire n_12080;
wire n_5093;
wire n_4052;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_9668;
wire n_3558;
wire n_10372;
wire n_7559;
wire n_5438;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_13259;
wire n_4326;
wire n_12702;
wire n_5517;
wire n_13175;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_3401;
wire n_10744;
wire n_12648;
wire n_3242;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_5907;
wire n_11334;
wire n_6045;
wire n_13075;
wire n_13129;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_7526;
wire n_5040;
wire n_6063;
wire n_10736;
wire n_10917;
wire n_6504;
wire n_3761;
wire n_11575;
wire n_4315;
wire n_2923;
wire n_7004;
wire n_7821;
wire n_12407;
wire n_8308;
wire n_6154;
wire n_11284;
wire n_6943;
wire n_4301;
wire n_10597;
wire n_11827;
wire n_13049;
wire n_3744;
wire n_8165;
wire n_12038;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_8210;
wire n_11656;
wire n_12644;
wire n_5977;
wire n_10446;
wire n_13134;
wire n_11826;
wire n_7879;
wire n_10271;
wire n_3814;
wire n_3781;
wire n_10888;
wire n_10116;
wire n_7696;
wire n_11570;
wire n_6003;
wire n_12952;
wire n_6684;
wire n_3843;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_5451;
wire n_9323;
wire n_3687;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_9331;
wire n_3621;
wire n_6031;
wire n_10170;
wire n_9922;
wire n_13252;
wire n_11909;
wire n_8331;
wire n_12024;
wire n_13084;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_12004;
wire n_3216;
wire n_12830;
wire n_12637;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_4365;
wire n_6060;
wire n_7929;
wire n_10255;
wire n_10572;
wire n_3726;
wire n_12009;
wire n_7270;
wire n_11490;
wire n_3758;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_10113;
wire n_7550;
wire n_3199;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_3339;
wire n_6853;
wire n_6742;
wire n_10188;
wire n_4923;
wire n_5864;
wire n_10686;
wire n_9841;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_12681;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_6172;
wire n_3343;
wire n_12634;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_8627;
wire n_9513;
wire n_9863;
wire n_12680;
wire n_11613;
wire n_4885;
wire n_10233;
wire n_12034;
wire n_10500;
wire n_10555;
wire n_5432;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_11929;
wire n_10810;
wire n_11075;
wire n_7851;
wire n_6894;
wire n_12176;
wire n_9791;
wire n_10311;
wire n_9179;
wire n_5453;
wire n_3658;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_3034;
wire n_11177;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_6817;
wire n_5842;
wire n_10937;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_12449;
wire n_5814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_11310;
wire n_12094;
wire n_6215;
wire n_3231;
wire n_11165;
wire n_4212;
wire n_9736;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_12823;
wire n_2953;
wire n_12517;
wire n_6517;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_10167;
wire n_7862;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_2946;
wire n_11923;
wire n_12071;
wire n_3430;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_8808;
wire n_10061;
wire n_12963;
wire n_10428;
wire n_13087;
wire n_11865;
wire n_12366;
wire n_8528;
wire n_8204;
wire n_13024;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_5495;
wire n_10694;
wire n_12339;
wire n_10602;
wire n_7100;
wire n_12729;
wire n_3583;
wire n_12198;
wire n_3860;
wire n_11041;
wire n_9420;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_9708;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_8154;
wire n_6966;
wire n_8889;
wire n_3015;
wire n_9790;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_4009;
wire n_5002;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_13258;
wire n_6035;
wire n_3473;
wire n_7874;
wire n_8490;
wire n_7622;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_13166;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_6364;
wire n_8635;
wire n_3241;
wire n_7420;
wire n_7102;
wire n_4342;
wire n_12605;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_7831;
wire n_6253;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_8532;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_3100;
wire n_11140;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_8796;
wire n_12218;
wire n_4106;
wire n_5737;
wire n_3604;
wire n_12343;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_12597;
wire n_12316;
wire n_4711;
wire n_11478;
wire n_12834;
wire n_3068;
wire n_10066;
wire n_13017;
wire n_12236;
wire n_12902;
wire n_6419;
wire n_8372;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_3553;
wire n_10088;
wire n_13038;
wire n_7225;
wire n_8077;
wire n_12892;
wire n_3811;
wire n_11294;
wire n_3494;
wire n_6244;
wire n_9812;
wire n_6900;
wire n_9337;
wire n_3486;
wire n_4086;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_9432;
wire n_9949;
wire n_10289;
wire n_6942;
wire n_7705;
wire n_11819;
wire n_7228;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_7932;
wire n_4812;
wire n_11573;
wire n_4409;
wire n_9576;
wire n_7509;
wire n_10145;
wire n_5872;
wire n_6862;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_6840;
wire n_13005;
wire n_3181;
wire n_6338;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_6037;
wire n_7981;
wire n_9577;
wire n_9874;
wire n_3699;
wire n_12588;
wire n_4913;
wire n_12589;
wire n_6266;
wire n_5874;
wire n_6488;
wire n_8337;
wire n_7164;
wire n_9231;
wire n_11844;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_11364;
wire n_3868;
wire n_9569;
wire n_13184;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_8358;
wire n_10009;
wire n_9552;
wire n_12927;
wire n_11100;
wire n_9279;
wire n_11902;
wire n_6317;
wire n_8199;
wire n_5588;
wire n_11993;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_10443;
wire n_8656;
wire n_7167;
wire n_10756;
wire n_12813;
wire n_6480;
wire n_3645;
wire n_10918;
wire n_13122;
wire n_5075;
wire n_11797;
wire n_3682;
wire n_3304;
wire n_4968;
wire n_3771;
wire n_12765;
wire n_7865;
wire n_12663;
wire n_10384;
wire n_9289;
wire n_5085;
wire n_11315;
wire n_5736;
wire n_4259;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_7134;
wire n_9633;
wire n_11153;
wire n_12312;
wire n_3422;
wire n_10074;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_4104;
wire n_9547;
wire n_13097;
wire n_6875;
wire n_10934;
wire n_10197;
wire n_8346;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_8761;
wire n_13112;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_8226;
wire n_11949;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_9084;
wire n_5928;
wire n_12256;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_11746;
wire n_11812;
wire n_3219;
wire n_9371;
wire n_13163;
wire n_3702;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_4779;
wire n_7267;
wire n_10367;
wire n_4599;
wire n_3233;
wire n_12315;
wire n_11505;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_12375;
wire n_12556;
wire n_3310;
wire n_3264;
wire n_12998;
wire n_7812;
wire n_7103;
wire n_13143;
wire n_9080;
wire n_4061;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_9519;
wire n_6367;
wire n_3881;
wire n_11363;
wire n_12156;
wire n_13128;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_11530;
wire n_12671;
wire n_10621;
wire n_7056;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_13260;
wire n_4642;
wire n_4051;
wire n_7813;
wire n_10085;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_6080;
wire n_4865;
wire n_8182;
wire n_8387;
wire n_12525;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_12076;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_7200;
wire n_11359;
wire n_3206;
wire n_7688;
wire n_4562;
wire n_3383;
wire n_8707;
wire n_12357;
wire n_4903;
wire n_3709;
wire n_10561;
wire n_11434;
wire n_3738;
wire n_9208;
wire n_11791;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_13212;
wire n_8494;
wire n_5812;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_11848;
wire n_3610;
wire n_11152;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_11632;
wire n_7795;
wire n_12180;
wire n_8788;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_7723;
wire n_4341;
wire n_11621;
wire n_10160;
wire n_9327;
wire n_10560;
wire n_7404;
wire n_12857;
wire n_13171;
wire n_5368;
wire n_4263;
wire n_8177;
wire n_3555;
wire n_9854;
wire n_7059;
wire n_7450;
wire n_11667;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_12208;
wire n_6145;
wire n_11964;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_3110;
wire n_7271;
wire n_7826;
wire n_9713;
wire n_11298;
wire n_5933;
wire n_8993;
wire n_6204;
wire n_7076;
wire n_4780;
wire n_10300;
wire n_9588;
wire n_11403;
wire n_11741;
wire n_12383;
wire n_11912;
wire n_4973;
wire n_3908;
wire n_6842;
wire n_3467;
wire n_12773;
wire n_6866;
wire n_9044;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_3950;
wire n_9423;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_2927;
wire n_4750;
wire n_12962;
wire n_6451;
wire n_9813;
wire n_3039;
wire n_9127;
wire n_6514;
wire n_3740;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_3186;
wire n_7105;
wire n_10140;
wire n_12612;
wire n_9244;
wire n_9869;
wire n_11142;
wire n_7049;
wire n_5903;
wire n_5986;
wire n_3065;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_12885;
wire n_11644;
wire n_6345;
wire n_9715;
wire n_8618;
wire n_3387;
wire n_12108;
wire n_9094;
wire n_13108;
wire n_5782;
wire n_7535;
wire n_3420;
wire n_5041;
wire n_13170;
wire n_4275;
wire n_10862;
wire n_11531;
wire n_4283;
wire n_4959;
wire n_8248;
wire n_8911;
wire n_9056;
wire n_11357;
wire n_4426;
wire n_9407;
wire n_11476;
wire n_4425;
wire n_3409;
wire n_9985;
wire n_4449;
wire n_12089;
wire n_12496;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_11959;
wire n_11367;
wire n_3002;
wire n_6957;
wire n_9361;
wire n_11921;
wire n_4809;
wire n_8495;
wire n_12676;
wire n_8783;
wire n_12987;
wire n_11566;
wire n_3392;
wire n_8529;
wire n_8733;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_10254;
wire n_7944;
wire n_13080;
wire n_11208;
wire n_7262;
wire n_3773;
wire n_8647;
wire n_11374;
wire n_12967;
wire n_12452;
wire n_8574;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_12232;
wire n_3301;
wire n_4241;
wire n_11859;
wire n_12818;
wire n_10386;
wire n_12128;
wire n_6379;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_5563;
wire n_11026;
wire n_8044;
wire n_2977;
wire n_5840;
wire n_6719;
wire n_7178;
wire n_9439;
wire n_9553;
wire n_11633;
wire n_11467;
wire n_7506;
wire n_12672;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_8330;
wire n_12760;
wire n_4050;
wire n_6232;
wire n_9132;
wire n_13172;
wire n_5717;
wire n_6017;
wire n_9696;
wire n_10861;
wire n_9120;
wire n_8879;
wire n_11203;
wire n_11159;
wire n_8052;
wire n_12168;
wire n_4578;
wire n_6362;
wire n_4777;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_8903;
wire n_11030;
wire n_4702;
wire n_12590;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_12924;
wire n_7142;
wire n_12577;
wire n_10182;
wire n_12732;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_10073;
wire n_4531;
wire n_3282;
wire n_11655;
wire n_5072;
wire n_3626;
wire n_11017;
wire n_7241;
wire n_7247;
wire n_12843;
wire n_12069;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_10333;
wire n_12430;
wire n_10317;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_7235;
wire n_8540;
wire n_11248;
wire n_12613;
wire n_6239;
wire n_12270;
wire n_9915;
wire n_4617;
wire n_9325;
wire n_9196;
wire n_4010;
wire n_5896;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_11141;
wire n_5105;
wire n_12695;
wire n_10893;
wire n_4308;
wire n_11093;
wire n_5021;
wire n_9251;
wire n_3463;
wire n_11576;
wire n_8939;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_8468;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_13181;
wire n_5134;
wire n_7096;
wire n_3063;
wire n_12210;
wire n_8778;
wire n_11197;
wire n_3998;
wire n_7442;
wire n_3632;
wire n_10093;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_6174;
wire n_12006;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_6087;
wire n_7593;
wire n_12246;
wire n_5249;
wire n_8068;
wire n_9955;
wire n_3829;
wire n_10539;
wire n_4164;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_4919;
wire n_3737;
wire n_10107;
wire n_5969;
wire n_3655;
wire n_10121;
wire n_10196;
wire n_8198;
wire n_3825;
wire n_3225;
wire n_13085;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_13224;
wire n_11469;
wire n_6454;
wire n_5022;
wire n_12625;
wire n_9270;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_8557;
wire n_6041;
wire n_6918;
wire n_9099;
wire n_12389;
wire n_9309;
wire n_3296;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_10814;
wire n_5276;
wire n_9627;
wire n_11252;
wire n_8012;
wire n_7672;
wire n_11494;
wire n_6664;
wire n_5047;
wire n_7318;
wire n_2985;
wire n_6472;
wire n_10218;
wire n_8114;
wire n_13131;
wire n_3792;
wire n_4202;
wire n_12995;
wire n_3938;
wire n_13209;
wire n_4791;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_5879;
wire n_8062;
wire n_4403;
wire n_11883;
wire n_5238;
wire n_11256;
wire n_11832;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_12370;
wire n_3531;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_10975;
wire n_11901;
wire n_6352;
wire n_12974;
wire n_9460;
wire n_8542;
wire n_12136;
wire n_10859;
wire n_13078;
wire n_7063;
wire n_7047;
wire n_11652;
wire n_4139;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_6238;
wire n_10542;
wire n_8038;
wire n_3931;
wire n_4349;
wire n_10681;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_11572;
wire n_5141;
wire n_11894;
wire n_3603;
wire n_10222;
wire n_6724;
wire n_13113;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_8716;
wire n_11336;
wire n_6705;
wire n_3822;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_4163;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_7074;
wire n_3812;
wire n_3910;
wire n_8734;
wire n_9204;
wire n_9476;
wire n_9689;
wire n_11849;
wire n_12142;
wire n_10659;
wire n_6591;
wire n_7585;
wire n_4948;
wire n_12564;
wire n_5268;
wire n_9780;
wire n_6946;
wire n_3482;
wire n_6002;
wire n_4080;
wire n_3319;
wire n_10403;
wire n_12983;
wire n_7037;
wire n_6289;
wire n_3748;
wire n_3272;
wire n_11784;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_3396;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_12886;
wire n_6532;
wire n_4372;
wire n_7293;
wire n_13000;
wire n_12035;
wire n_13006;
wire n_5640;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_6721;
wire n_5560;
wire n_13205;
wire n_6644;
wire n_6512;
wire n_5544;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_12810;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_4918;
wire n_3824;
wire n_9597;
wire n_5067;
wire n_11322;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_11892;
wire n_12122;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_12241;
wire n_12396;
wire n_7614;
wire n_9343;
wire n_2941;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_4032;
wire n_6086;
wire n_9837;
wire n_11421;
wire n_11057;
wire n_4147;
wire n_10896;
wire n_10969;
wire n_4477;
wire n_11966;
wire n_12748;
wire n_3168;
wire n_7383;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_10562;
wire n_5941;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_5611;
wire n_3601;
wire n_6340;
wire n_10054;
wire n_3092;
wire n_6219;
wire n_10355;
wire n_3055;
wire n_6706;
wire n_7479;
wire n_3966;
wire n_11853;
wire n_12571;
wire n_9692;
wire n_7395;
wire n_10598;
wire n_13034;
wire n_8947;
wire n_4742;
wire n_3734;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_7078;
wire n_8188;
wire n_6761;
wire n_8972;
wire n_10007;
wire n_3649;
wire n_11751;
wire n_11423;
wire n_11725;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_12674;
wire n_8510;
wire n_11410;
wire n_3384;
wire n_12230;
wire n_9567;
wire n_6811;
wire n_9061;
wire n_11495;
wire n_3419;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_4478;
wire n_7372;
wire n_5367;
wire n_3794;
wire n_12220;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_10704;
wire n_11520;
wire n_11622;
wire n_4838;
wire n_5970;
wire n_12169;
wire n_12283;
wire n_12336;
wire n_7174;
wire n_13268;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_10457;
wire n_12543;
wire n_4965;
wire n_8021;
wire n_3346;
wire n_9705;
wire n_7803;
wire n_11012;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_12595;
wire n_9624;
wire n_3861;
wire n_9701;
wire n_11502;
wire n_11429;
wire n_10389;
wire n_11631;
wire n_3891;
wire n_6659;
wire n_4523;
wire n_9709;
wire n_6011;
wire n_9295;
wire n_9416;
wire n_4371;
wire n_6225;
wire n_11842;
wire n_12463;
wire n_10990;
wire n_2994;
wire n_11640;
wire n_5502;
wire n_12263;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_9929;
wire n_12920;
wire n_10264;
wire n_5850;
wire n_4673;
wire n_9953;
wire n_7086;
wire n_3415;
wire n_6648;
wire n_4607;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_12717;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_12141;
wire n_8584;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_13196;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_11904;
wire n_8480;
wire n_10301;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_13018;
wire n_7025;
wire n_9364;
wire n_8228;
wire n_2976;
wire n_8076;
wire n_6826;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_9836;
wire n_10929;
wire n_9107;
wire n_3809;
wire n_11279;
wire n_11724;
wire n_13044;
wire n_11789;
wire n_3139;
wire n_13228;
wire n_11525;
wire n_8100;
wire n_4070;
wire n_11999;
wire n_13086;
wire n_10837;
wire n_3545;
wire n_3885;
wire n_10554;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_12746;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_10149;
wire n_10970;
wire n_7768;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_5496;
wire n_3780;
wire n_5802;
wire n_7982;
wire n_12190;
wire n_12787;
wire n_8804;
wire n_3337;
wire n_11383;
wire n_12799;
wire n_4002;
wire n_11847;
wire n_11976;
wire n_3209;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_5547;
wire n_8158;
wire n_12511;
wire n_11167;
wire n_6879;
wire n_12532;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_3477;
wire n_8433;
wire n_10102;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_5983;
wire n_8213;
wire n_3146;
wire n_3953;
wire n_4588;
wire n_10534;
wire n_11825;
wire n_4653;
wire n_4435;
wire n_11049;
wire n_10619;
wire n_7684;
wire n_10932;
wire n_5604;
wire n_8451;
wire n_5411;
wire n_8334;
wire n_12743;
wire n_4019;
wire n_8731;
wire n_10589;
wire n_11681;
wire n_11611;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_11202;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_5815;
wire n_3616;
wire n_7370;
wire n_9748;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_8539;
wire n_10205;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_9226;
wire n_3727;
wire n_5235;
wire n_10110;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_11688;
wire n_6888;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_12715;
wire n_11709;
wire n_12434;
wire n_12628;
wire n_8122;
wire n_6095;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_11331;
wire n_5311;
wire n_12979;
wire n_9528;
wire n_6590;
wire n_10638;
wire n_7583;
wire n_12201;
wire n_3522;
wire n_6559;
wire n_12499;
wire n_3924;
wire n_9112;
wire n_12448;
wire n_4621;
wire n_4216;
wire n_11876;
wire n_5797;
wire n_9235;
wire n_10610;
wire n_11187;
wire n_4240;
wire n_12761;
wire n_5572;
wire n_3491;
wire n_9333;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_8950;
wire n_10758;
wire n_10190;
wire n_5520;
wire n_3353;
wire n_11804;
wire n_3975;
wire n_3018;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_6287;
wire n_12809;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_7353;
wire n_9330;
wire n_12538;
wire n_7758;
wire n_4021;
wire n_12446;
wire n_9490;
wire n_3014;
wire n_12029;
wire n_4103;
wire n_9355;
wire n_11052;
wire n_5060;
wire n_9523;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_9582;
wire n_4775;
wire n_5884;
wire n_10060;
wire n_6671;
wire n_11009;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_9288;
wire n_9686;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_13068;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_11446;
wire n_10910;
wire n_10162;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_13248;
wire n_7792;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_2958;
wire n_8703;
wire n_10014;
wire n_7109;
wire n_12642;
wire n_3731;
wire n_2936;
wire n_3224;
wire n_12484;
wire n_6128;
wire n_8822;
wire n_6029;
wire n_10677;
wire n_12187;
wire n_5751;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_12321;
wire n_5924;
wire n_9992;
wire n_11247;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_12669;
wire n_13106;
wire n_3129;
wire n_8476;
wire n_6702;
wire n_11927;
wire n_3620;
wire n_11179;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_3693;
wire n_8545;
wire n_8736;
wire n_9051;
wire n_4497;
wire n_7749;
wire n_10105;
wire n_10078;
wire n_11514;
wire n_12470;
wire n_12994;
wire n_11321;
wire n_9500;
wire n_8705;
wire n_10215;
wire n_11779;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_5694;
wire n_3203;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_10834;
wire n_7574;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_4306;
wire n_11882;
wire n_11647;
wire n_4224;
wire n_12064;
wire n_10706;
wire n_12462;
wire n_3341;
wire n_6005;
wire n_8872;
wire n_12696;
wire n_4453;
wire n_9555;
wire n_11133;
wire n_5449;
wire n_3559;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_3546;
wire n_3661;
wire n_12735;
wire n_7713;
wire n_4564;
wire n_11222;
wire n_9200;
wire n_5146;
wire n_10709;
wire n_3056;
wire n_12646;
wire n_3201;
wire n_10871;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_3103;
wire n_10304;
wire n_5398;
wire n_4573;
wire n_5860;
wire n_6936;
wire n_4535;
wire n_10244;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_7641;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_7203;
wire n_12999;
wire n_9397;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_12682;
wire n_3612;
wire n_9673;
wire n_4695;
wire n_6848;
wire n_8642;
wire n_3509;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11941;
wire n_11875;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_12111;
wire n_8912;
wire n_2966;
wire n_7439;
wire n_9496;
wire n_3196;
wire n_8110;
wire n_5319;
wire n_10796;
wire n_10016;
wire n_9008;
wire n_12903;
wire n_12079;
wire n_6343;
wire n_12593;
wire n_5270;
wire n_10030;
wire n_8805;
wire n_6850;
wire n_12864;
wire n_5005;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_11307;
wire n_5181;
wire n_6979;
wire n_7815;
wire n_13222;
wire n_7934;
wire n_9545;
wire n_3144;
wire n_8111;
wire n_3244;
wire n_9603;
wire n_9629;
wire n_11578;
wire n_6865;
wire n_10432;
wire n_12719;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_3287;
wire n_3322;
wire n_5043;
wire n_8739;
wire n_6747;
wire n_9674;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_10462;
wire n_12725;
wire n_3640;
wire n_3481;
wire n_6640;
wire n_11769;
wire n_8856;
wire n_3033;
wire n_6142;
wire n_9930;
wire n_11908;
wire n_12925;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_6034;
wire n_9781;
wire n_10291;
wire n_13159;
wire n_4597;
wire n_9659;
wire n_3364;
wire n_3226;
wire n_4020;
wire n_7233;
wire n_8732;
wire n_11913;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_11341;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_13256;
wire n_10669;
wire n_6870;
wire n_6221;
wire n_8231;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_4063;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_4237;
wire n_5029;
wire n_5127;
wire n_12317;
wire n_6071;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_8908;
wire n_10185;
wire n_11182;
wire n_3212;
wire n_10092;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_12782;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_11231;
wire n_3093;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_12875;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_8137;
wire n_7045;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_3169;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_11727;
wire n_6788;
wire n_7014;
wire n_12192;
wire n_12633;
wire n_10430;
wire n_8305;
wire n_4614;
wire n_3360;
wire n_10277;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_6709;
wire n_4422;
wire n_10948;
wire n_11749;
wire n_6550;
wire n_6712;
wire n_10525;
wire n_9507;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_3004;
wire n_8841;
wire n_3870;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_6743;
wire n_12497;
wire n_4632;
wire n_10354;
wire n_12412;
wire n_3084;
wire n_11880;
wire n_5785;
wire n_7465;
wire n_13177;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_12724;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_9485;
wire n_4966;
wire n_2942;
wire n_9457;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_7936;
wire n_8966;
wire n_6084;
wire n_11249;
wire n_4847;
wire n_10287;
wire n_4054;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_12101;
wire n_10119;
wire n_11145;
wire n_3586;
wire n_12606;
wire n_11986;
wire n_3653;
wire n_8395;
wire n_10900;
wire n_5966;
wire n_10349;
wire n_6634;
wire n_4668;
wire n_3349;
wire n_5213;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_13229;
wire n_5735;
wire n_12118;
wire n_7490;
wire n_11380;
wire n_7545;
wire n_10792;
wire n_11513;
wire n_8625;
wire n_7160;
wire n_7464;
wire n_9809;
wire n_8937;
wire n_4214;
wire n_6919;
wire n_10750;
wire n_3448;
wire n_7805;
wire n_10995;
wire n_13092;
wire n_7115;
wire n_7295;
wire n_2924;
wire n_12087;
wire n_9192;
wire n_3595;
wire n_7348;
wire n_5752;
wire n_11618;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_10537;
wire n_11861;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_10426;
wire n_4405;
wire n_4413;
wire n_9558;
wire n_11594;
wire n_7453;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_4036;
wire n_10684;
wire n_4759;
wire n_7162;
wire n_3670;
wire n_11436;
wire n_12346;
wire n_4667;
wire n_5081;
wire n_11729;
wire n_4182;
wire n_3230;
wire n_8371;
wire n_8702;
wire n_8116;
wire n_8195;
wire n_7946;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_12244;
wire n_5877;
wire n_9991;
wire n_11670;
wire n_11366;
wire n_11872;
wire n_7681;
wire n_8845;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_5189;
wire n_7702;
wire n_6676;
wire n_8149;
wire n_10823;
wire n_3041;
wire n_4637;
wire n_9976;
wire n_8042;
wire n_11516;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_8392;
wire n_9560;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_10830;
wire n_11132;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_6854;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_4977;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_6032;
wire n_9047;
wire n_12953;
wire n_12842;
wire n_3650;
wire n_8968;
wire n_12481;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_5446;
wire n_11316;
wire n_3010;
wire n_7855;
wire n_3043;
wire n_11047;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_4590;
wire n_8399;
wire n_5090;
wire n_3137;
wire n_9599;
wire n_11767;
wire n_3560;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_3177;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_12435;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_11586;
wire n_6981;
wire n_7065;
wire n_12149;
wire n_9216;
wire n_3238;
wire n_3529;
wire n_12002;
wire n_12836;
wire n_4835;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_11229;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_4038;
wire n_6122;
wire n_11225;
wire n_11397;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_12840;
wire n_3784;
wire n_7330;
wire n_5437;
wire n_8883;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_10577;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_7357;
wire n_8756;
wire n_11324;
wire n_8737;
wire n_10334;
wire n_4434;
wire n_12945;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_10151;
wire n_6439;
wire n_11614;
wire n_4290;
wire n_8602;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_5407;
wire n_10411;
wire n_13249;
wire n_9484;
wire n_12984;
wire n_10989;
wire n_8422;
wire n_3029;
wire n_10939;
wire n_12224;
wire n_5913;
wire n_3597;
wire n_7088;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_8878;
wire n_11144;
wire n_10090;
wire n_6406;
wire n_7440;
wire n_11361;
wire n_6945;
wire n_8112;
wire n_11567;
wire n_3790;
wire n_10962;
wire n_7029;
wire n_11128;
wire n_9292;
wire n_9622;
wire n_10721;
wire n_8593;
wire n_12197;
wire n_10186;
wire n_3318;
wire n_4833;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_6618;
wire n_6474;
wire n_13082;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_13094;
wire n_7317;
wire n_10856;
wire n_12403;
wire n_6000;
wire n_3350;
wire n_12679;
wire n_9584;
wire n_3977;
wire n_8194;
wire n_9461;
wire n_8055;
wire n_11168;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_8360;
wire n_3588;
wire n_5008;
wire n_4279;
wire n_12018;
wire n_6425;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_9845;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_11937;
wire n_12872;
wire n_7522;
wire n_6492;
wire n_10071;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_6046;
wire n_11460;
wire n_8251;
wire n_5323;
wire n_11565;
wire n_3388;
wire n_4790;
wire n_4181;
wire n_3184;
wire n_12372;
wire n_9618;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_11192;
wire n_11808;
wire n_4007;
wire n_13257;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_4239;
wire n_8677;
wire n_13052;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_5991;
wire n_4184;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_2986;
wire n_5702;
wire n_10035;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_9699;
wire n_12340;
wire n_3489;
wire n_8108;
wire n_5243;
wire n_5914;
wire n_12955;
wire n_12068;
wire n_10252;
wire n_5250;
wire n_11555;
wire n_3074;
wire n_6869;
wire n_3102;
wire n_10041;
wire n_9321;
wire n_5590;
wire n_10345;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_3321;
wire n_5809;
wire n_10543;
wire n_3377;
wire n_7924;
wire n_4782;
wire n_12394;
wire n_7659;
wire n_9005;
wire n_3530;
wire n_9161;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_12954;
wire n_7836;
wire n_10737;
wire n_12662;
wire n_4876;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_7280;
wire n_10644;
wire n_12801;
wire n_5813;
wire n_9293;
wire n_12503;
wire n_10365;
wire n_5833;
wire n_11781;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_12965;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_10809;
wire n_8927;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_6228;
wire n_6711;
wire n_11997;
wire n_3483;
wire n_11884;
wire n_5416;
wire n_8946;
wire n_13090;
wire n_12822;
wire n_11863;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_9646;
wire n_8017;
wire n_12264;
wire n_11761;
wire n_8474;
wire n_9984;
wire n_3524;
wire n_7275;
wire n_8232;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_9649;
wire n_8904;
wire n_11199;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_10629;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_8382;
wire n_4421;
wire n_13023;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_4793;
wire n_4498;
wire n_10006;
wire n_11757;
wire n_7259;
wire n_12320;
wire n_12274;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_12622;
wire n_6992;
wire n_11185;
wire n_2944;
wire n_8128;
wire n_12659;
wire n_6818;
wire n_3831;
wire n_10206;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5932;
wire n_5830;
wire n_3589;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_7539;
wire n_12586;
wire n_3391;
wire n_12629;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_10275;
wire n_11081;
wire n_3458;
wire n_7775;
wire n_13011;
wire n_4505;
wire n_11392;
wire n_9981;
wire n_3190;
wire n_7930;
wire n_5558;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_8205;
wire n_5051;
wire n_9907;
wire n_13088;
wire n_5587;
wire n_6976;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_12269;
wire n_7640;
wire n_9816;
wire n_10498;
wire n_11424;
wire n_12585;
wire n_5012;
wire n_11463;
wire n_10292;
wire n_6864;
wire n_7969;
wire n_8605;
wire n_11278;
wire n_10358;
wire n_3787;
wire n_7548;
wire n_3585;
wire n_10635;
wire n_3565;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_12832;
wire n_12913;
wire n_5025;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_12301;
wire n_3135;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_7197;
wire n_9676;
wire n_5645;
wire n_3990;
wire n_11881;
wire n_7393;
wire n_11332;
wire n_6917;
wire n_6937;
wire n_7591;
wire n_13207;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_7727;
wire n_7358;
wire n_7324;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_11935;
wire n_4534;
wire n_6301;
wire n_9788;
wire n_6929;
wire n_11309;
wire n_8719;
wire n_8045;
wire n_10785;
wire n_7729;
wire n_2969;
wire n_12341;
wire n_12615;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_8209;
wire n_10802;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_6699;
wire n_12926;
wire n_9213;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_8784;
wire n_7382;
wire n_4811;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_12167;
wire n_9473;
wire n_4857;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_6677;
wire n_12161;
wire n_3432;
wire n_12085;
wire n_11735;
wire n_7618;
wire n_4282;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_6764;
wire n_8575;
wire n_12298;
wire n_10081;
wire n_5733;
wire n_3774;
wire n_10324;
wire n_6780;
wire n_11189;
wire n_8815;
wire n_11582;
wire n_12569;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_3268;
wire n_9303;
wire n_11105;
wire n_3057;
wire n_11705;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_7673;
wire n_6830;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_7282;
wire n_6586;
wire n_9968;
wire n_10808;
wire n_11474;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_7953;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_9722;
wire n_12042;
wire n_12155;
wire n_5657;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_8695;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_4911;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_4436;
wire n_8363;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_8665;
wire n_13098;
wire n_6510;
wire n_8282;
wire n_3334;
wire n_9388;
wire n_5938;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_12654;
wire n_5602;
wire n_9379;
wire n_11992;
wire n_5097;
wire n_4985;
wire n_7751;
wire n_10869;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_13142;
wire n_7581;
wire n_13180;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_3584;
wire n_5246;
wire n_10453;
wire n_12386;
wire n_4858;
wire n_4678;
wire n_9952;
wire n_3556;
wire n_9911;
wire n_12183;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_12419;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_12964;
wire n_10473;
wire n_5107;
wire n_5095;
wire n_3456;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_11439;
wire n_10957;
wire n_4243;
wire n_7579;
wire n_12863;
wire n_10352;
wire n_4025;
wire n_11188;
wire n_7428;
wire n_3404;
wire n_5666;
wire n_12221;
wire n_4059;
wire n_9195;
wire n_10442;
wire n_11687;
wire n_4121;
wire n_3290;
wire n_8870;
wire n_7155;
wire n_7150;
wire n_8252;
wire n_11774;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_6475;
wire n_4142;
wire n_7283;
wire n_7015;
wire n_3982;
wire n_7699;
wire n_8507;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_13206;
wire n_9623;
wire n_6103;
wire n_5546;
wire n_7249;
wire n_10713;
wire n_3796;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_10954;
wire n_4246;
wire n_12267;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_4532;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_11329;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_9516;
wire n_4244;
wire n_13241;
wire n_13187;
wire n_13162;
wire n_4049;
wire n_6752;
wire n_12768;
wire n_8976;
wire n_6426;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_8156;
wire n_11661;
wire n_7494;
wire n_4353;
wire n_11120;
wire n_9222;
wire n_13031;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_4787;
wire n_7736;
wire n_10622;
wire n_5633;
wire n_13155;
wire n_9546;
wire n_5664;
wire n_7589;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_13066;
wire n_8660;
wire n_11296;
wire n_8479;
wire n_12993;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_3521;
wire n_11314;
wire n_8723;
wire n_11019;
wire n_8606;
wire n_9663;
wire n_6235;
wire n_7843;
wire n_8235;
wire n_13083;
wire n_3764;
wire n_12647;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_9820;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_9743;
wire n_6496;
wire n_3066;
wire n_7756;
wire n_12749;
wire n_8342;
wire n_8940;
wire n_13048;
wire n_11584;
wire n_5280;
wire n_8448;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_4332;
wire n_7555;
wire n_10000;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_10582;
wire n_12066;
wire n_12812;
wire n_3695;
wire n_10427;
wire n_11816;
wire n_12060;
wire n_3976;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_3563;
wire n_6513;
wire n_7500;
wire n_10246;
wire n_11910;
wire n_3198;
wire n_11693;
wire n_3495;
wire n_5925;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_9822;
wire n_10835;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_3359;
wire n_12164;
wire n_5272;
wire n_11368;
wire n_10125;
wire n_12824;
wire n_13111;
wire n_6330;
wire n_10117;
wire n_9065;
wire n_3187;
wire n_12716;
wire n_10844;
wire n_3218;
wire n_8457;
wire n_6802;
wire n_10654;
wire n_9153;
wire n_9086;
wire n_10505;
wire n_9339;
wire n_10198;
wire n_6909;
wire n_7157;
wire n_11064;
wire n_13237;
wire n_6908;
wire n_8237;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_11409;
wire n_4201;
wire n_2968;
wire n_4336;
wire n_7266;
wire n_8046;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_12437;
wire n_5624;
wire n_4852;
wire n_4981;
wire n_4210;
wire n_10840;
wire n_12052;
wire n_6477;
wire n_9746;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_5440;
wire n_6490;
wire n_11533;
wire n_11605;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_7198;
wire n_8335;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_9440;
wire n_10144;
wire n_3955;
wire n_9684;
wire n_6184;
wire n_3945;
wire n_5817;
wire n_5214;
wire n_10973;
wire n_4936;
wire n_4205;
wire n_9493;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_3433;
wire n_11330;
wire n_12720;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_6038;
wire n_10551;
wire n_5861;
wire n_3833;
wire n_10553;
wire n_13127;
wire n_3162;
wire n_8309;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_12687;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_9032;
wire n_9814;
wire n_6313;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_13208;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_5859;
wire n_12325;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_5776;
wire n_8166;
wire n_5606;
wire n_4433;
wire n_3085;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_5826;
wire n_10108;
wire n_8960;
wire n_12789;
wire n_5920;
wire n_2991;
wire n_10307;
wire n_5030;
wire n_4194;
wire n_7994;
wire n_4703;
wire n_8443;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_6180;
wire n_8683;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_12127;
wire n_12382;
wire n_12504;
wire n_3182;
wire n_5756;
wire n_12602;
wire n_5527;
wire n_3283;
wire n_6476;
wire n_8037;
wire n_12062;
wire n_4030;
wire n_12573;

CKINVDCx5p33_ASAP7_75t_R g2921 ( 
.A(n_2269),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2812),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2674),
.Y(n_2923)
);

CKINVDCx5p33_ASAP7_75t_R g2924 ( 
.A(n_2441),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_1986),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_1093),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2759),
.Y(n_2927)
);

CKINVDCx20_ASAP7_75t_R g2928 ( 
.A(n_1894),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_1099),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_1893),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_899),
.Y(n_2931)
);

CKINVDCx5p33_ASAP7_75t_R g2932 ( 
.A(n_2729),
.Y(n_2932)
);

INVx1_ASAP7_75t_SL g2933 ( 
.A(n_1537),
.Y(n_2933)
);

CKINVDCx20_ASAP7_75t_R g2934 ( 
.A(n_1743),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_1239),
.Y(n_2935)
);

CKINVDCx5p33_ASAP7_75t_R g2936 ( 
.A(n_1752),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_570),
.Y(n_2937)
);

BUFx10_ASAP7_75t_L g2938 ( 
.A(n_2355),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_323),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_2742),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2807),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_1899),
.Y(n_2942)
);

CKINVDCx20_ASAP7_75t_R g2943 ( 
.A(n_1329),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_1582),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_1266),
.Y(n_2945)
);

CKINVDCx5p33_ASAP7_75t_R g2946 ( 
.A(n_2050),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_290),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_1090),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2497),
.Y(n_2949)
);

CKINVDCx20_ASAP7_75t_R g2950 ( 
.A(n_2756),
.Y(n_2950)
);

INVx1_ASAP7_75t_SL g2951 ( 
.A(n_598),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_1733),
.Y(n_2952)
);

CKINVDCx16_ASAP7_75t_R g2953 ( 
.A(n_2750),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_1900),
.Y(n_2954)
);

CKINVDCx5p33_ASAP7_75t_R g2955 ( 
.A(n_527),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_625),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_550),
.Y(n_2957)
);

CKINVDCx16_ASAP7_75t_R g2958 ( 
.A(n_1630),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2239),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2876),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_1809),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2644),
.Y(n_2962)
);

CKINVDCx5p33_ASAP7_75t_R g2963 ( 
.A(n_1422),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_1167),
.Y(n_2964)
);

INVx1_ASAP7_75t_SL g2965 ( 
.A(n_2873),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_2668),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_1680),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_555),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_1767),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_1873),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_1780),
.Y(n_2971)
);

CKINVDCx20_ASAP7_75t_R g2972 ( 
.A(n_2016),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_954),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_105),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2866),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_1419),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2920),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_152),
.Y(n_2978)
);

CKINVDCx5p33_ASAP7_75t_R g2979 ( 
.A(n_1089),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_1867),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2109),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2044),
.Y(n_2982)
);

INVx1_ASAP7_75t_SL g2983 ( 
.A(n_1568),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_885),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2675),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_988),
.Y(n_2986)
);

CKINVDCx16_ASAP7_75t_R g2987 ( 
.A(n_2850),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_470),
.Y(n_2988)
);

INVx1_ASAP7_75t_SL g2989 ( 
.A(n_1728),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2099),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_723),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_861),
.Y(n_2992)
);

CKINVDCx5p33_ASAP7_75t_R g2993 ( 
.A(n_1015),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_1252),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_1074),
.Y(n_2995)
);

CKINVDCx5p33_ASAP7_75t_R g2996 ( 
.A(n_1400),
.Y(n_2996)
);

CKINVDCx5p33_ASAP7_75t_R g2997 ( 
.A(n_1604),
.Y(n_2997)
);

BUFx3_ASAP7_75t_L g2998 ( 
.A(n_545),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2330),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_1784),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2617),
.Y(n_3001)
);

CKINVDCx5p33_ASAP7_75t_R g3002 ( 
.A(n_1567),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_1505),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_1350),
.Y(n_3004)
);

CKINVDCx20_ASAP7_75t_R g3005 ( 
.A(n_2173),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_789),
.Y(n_3006)
);

CKINVDCx5p33_ASAP7_75t_R g3007 ( 
.A(n_233),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_1346),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_1730),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_1723),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2725),
.Y(n_3011)
);

INVx4_ASAP7_75t_R g3012 ( 
.A(n_2854),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2181),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_153),
.Y(n_3014)
);

BUFx10_ASAP7_75t_L g3015 ( 
.A(n_1413),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_509),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2113),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_47),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_1875),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_399),
.Y(n_3020)
);

CKINVDCx20_ASAP7_75t_R g3021 ( 
.A(n_2137),
.Y(n_3021)
);

CKINVDCx5p33_ASAP7_75t_R g3022 ( 
.A(n_2692),
.Y(n_3022)
);

INVx2_ASAP7_75t_SL g3023 ( 
.A(n_2328),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_2687),
.Y(n_3024)
);

CKINVDCx5p33_ASAP7_75t_R g3025 ( 
.A(n_1425),
.Y(n_3025)
);

CKINVDCx5p33_ASAP7_75t_R g3026 ( 
.A(n_1708),
.Y(n_3026)
);

CKINVDCx20_ASAP7_75t_R g3027 ( 
.A(n_2139),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_1512),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_1148),
.Y(n_3029)
);

BUFx2_ASAP7_75t_SL g3030 ( 
.A(n_1433),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_1889),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_38),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_336),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_1544),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2803),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_1832),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_2849),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2902),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2663),
.Y(n_3039)
);

CKINVDCx5p33_ASAP7_75t_R g3040 ( 
.A(n_2262),
.Y(n_3040)
);

CKINVDCx5p33_ASAP7_75t_R g3041 ( 
.A(n_1641),
.Y(n_3041)
);

CKINVDCx5p33_ASAP7_75t_R g3042 ( 
.A(n_113),
.Y(n_3042)
);

CKINVDCx5p33_ASAP7_75t_R g3043 ( 
.A(n_438),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_342),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_1246),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_575),
.Y(n_3046)
);

CKINVDCx5p33_ASAP7_75t_R g3047 ( 
.A(n_2177),
.Y(n_3047)
);

INVx1_ASAP7_75t_SL g3048 ( 
.A(n_2748),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2648),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2625),
.Y(n_3050)
);

CKINVDCx20_ASAP7_75t_R g3051 ( 
.A(n_215),
.Y(n_3051)
);

INVx1_ASAP7_75t_SL g3052 ( 
.A(n_2378),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2395),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2149),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_1968),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_1300),
.Y(n_3056)
);

HB1xp67_ASAP7_75t_L g3057 ( 
.A(n_2471),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2051),
.Y(n_3058)
);

CKINVDCx5p33_ASAP7_75t_R g3059 ( 
.A(n_2227),
.Y(n_3059)
);

INVx3_ASAP7_75t_L g3060 ( 
.A(n_1613),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2194),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_2871),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_1095),
.Y(n_3063)
);

CKINVDCx5p33_ASAP7_75t_R g3064 ( 
.A(n_2652),
.Y(n_3064)
);

CKINVDCx5p33_ASAP7_75t_R g3065 ( 
.A(n_2758),
.Y(n_3065)
);

CKINVDCx5p33_ASAP7_75t_R g3066 ( 
.A(n_1678),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2658),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_1859),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2123),
.Y(n_3069)
);

HB1xp67_ASAP7_75t_L g3070 ( 
.A(n_2193),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_754),
.Y(n_3071)
);

BUFx10_ASAP7_75t_L g3072 ( 
.A(n_878),
.Y(n_3072)
);

CKINVDCx5p33_ASAP7_75t_R g3073 ( 
.A(n_2697),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2007),
.Y(n_3074)
);

CKINVDCx20_ASAP7_75t_R g3075 ( 
.A(n_1868),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_1170),
.Y(n_3076)
);

CKINVDCx5p33_ASAP7_75t_R g3077 ( 
.A(n_1680),
.Y(n_3077)
);

CKINVDCx5p33_ASAP7_75t_R g3078 ( 
.A(n_984),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_2531),
.Y(n_3079)
);

INVx1_ASAP7_75t_SL g3080 ( 
.A(n_2383),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_1821),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_1284),
.Y(n_3082)
);

BUFx6f_ASAP7_75t_L g3083 ( 
.A(n_284),
.Y(n_3083)
);

CKINVDCx5p33_ASAP7_75t_R g3084 ( 
.A(n_236),
.Y(n_3084)
);

CKINVDCx5p33_ASAP7_75t_R g3085 ( 
.A(n_1928),
.Y(n_3085)
);

BUFx10_ASAP7_75t_L g3086 ( 
.A(n_2604),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_1737),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_1684),
.Y(n_3088)
);

INVx1_ASAP7_75t_SL g3089 ( 
.A(n_2186),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_1935),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2875),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_2219),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_1749),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2748),
.Y(n_3094)
);

CKINVDCx5p33_ASAP7_75t_R g3095 ( 
.A(n_1879),
.Y(n_3095)
);

INVx1_ASAP7_75t_SL g3096 ( 
.A(n_2833),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2883),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2567),
.Y(n_3098)
);

CKINVDCx5p33_ASAP7_75t_R g3099 ( 
.A(n_1049),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_824),
.Y(n_3100)
);

CKINVDCx5p33_ASAP7_75t_R g3101 ( 
.A(n_794),
.Y(n_3101)
);

BUFx2_ASAP7_75t_SL g3102 ( 
.A(n_1234),
.Y(n_3102)
);

CKINVDCx5p33_ASAP7_75t_R g3103 ( 
.A(n_1073),
.Y(n_3103)
);

CKINVDCx16_ASAP7_75t_R g3104 ( 
.A(n_2831),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_2212),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_1857),
.Y(n_3106)
);

BUFx2_ASAP7_75t_L g3107 ( 
.A(n_607),
.Y(n_3107)
);

INVx1_ASAP7_75t_SL g3108 ( 
.A(n_1193),
.Y(n_3108)
);

CKINVDCx20_ASAP7_75t_R g3109 ( 
.A(n_2674),
.Y(n_3109)
);

BUFx5_ASAP7_75t_L g3110 ( 
.A(n_2594),
.Y(n_3110)
);

CKINVDCx5p33_ASAP7_75t_R g3111 ( 
.A(n_2744),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_2666),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2843),
.Y(n_3113)
);

CKINVDCx5p33_ASAP7_75t_R g3114 ( 
.A(n_1220),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2546),
.Y(n_3115)
);

CKINVDCx20_ASAP7_75t_R g3116 ( 
.A(n_1288),
.Y(n_3116)
);

CKINVDCx5p33_ASAP7_75t_R g3117 ( 
.A(n_2062),
.Y(n_3117)
);

CKINVDCx5p33_ASAP7_75t_R g3118 ( 
.A(n_871),
.Y(n_3118)
);

CKINVDCx20_ASAP7_75t_R g3119 ( 
.A(n_2743),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2823),
.Y(n_3120)
);

CKINVDCx5p33_ASAP7_75t_R g3121 ( 
.A(n_92),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_2112),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_324),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_598),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2230),
.Y(n_3125)
);

BUFx3_ASAP7_75t_L g3126 ( 
.A(n_2569),
.Y(n_3126)
);

INVx2_ASAP7_75t_SL g3127 ( 
.A(n_2291),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_2057),
.Y(n_3128)
);

CKINVDCx20_ASAP7_75t_R g3129 ( 
.A(n_1831),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_2299),
.Y(n_3130)
);

CKINVDCx5p33_ASAP7_75t_R g3131 ( 
.A(n_1208),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_2690),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_1275),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_576),
.Y(n_3134)
);

CKINVDCx5p33_ASAP7_75t_R g3135 ( 
.A(n_2042),
.Y(n_3135)
);

CKINVDCx5p33_ASAP7_75t_R g3136 ( 
.A(n_248),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2802),
.Y(n_3137)
);

CKINVDCx5p33_ASAP7_75t_R g3138 ( 
.A(n_2784),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_975),
.Y(n_3139)
);

BUFx6f_ASAP7_75t_L g3140 ( 
.A(n_2673),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2285),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_1883),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2203),
.Y(n_3143)
);

CKINVDCx5p33_ASAP7_75t_R g3144 ( 
.A(n_1149),
.Y(n_3144)
);

CKINVDCx20_ASAP7_75t_R g3145 ( 
.A(n_742),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2788),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_1152),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2552),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_2863),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2706),
.Y(n_3150)
);

BUFx2_ASAP7_75t_L g3151 ( 
.A(n_2132),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_2649),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_640),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2861),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_1676),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2827),
.Y(n_3156)
);

CKINVDCx5p33_ASAP7_75t_R g3157 ( 
.A(n_241),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_1651),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_996),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_259),
.Y(n_3160)
);

INVx1_ASAP7_75t_SL g3161 ( 
.A(n_2491),
.Y(n_3161)
);

HB1xp67_ASAP7_75t_L g3162 ( 
.A(n_1171),
.Y(n_3162)
);

CKINVDCx5p33_ASAP7_75t_R g3163 ( 
.A(n_2856),
.Y(n_3163)
);

CKINVDCx5p33_ASAP7_75t_R g3164 ( 
.A(n_2372),
.Y(n_3164)
);

CKINVDCx5p33_ASAP7_75t_R g3165 ( 
.A(n_2026),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_1085),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_274),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2464),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_422),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_2905),
.Y(n_3170)
);

CKINVDCx20_ASAP7_75t_R g3171 ( 
.A(n_1003),
.Y(n_3171)
);

CKINVDCx5p33_ASAP7_75t_R g3172 ( 
.A(n_1897),
.Y(n_3172)
);

CKINVDCx5p33_ASAP7_75t_R g3173 ( 
.A(n_2670),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2772),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2126),
.Y(n_3175)
);

CKINVDCx20_ASAP7_75t_R g3176 ( 
.A(n_2717),
.Y(n_3176)
);

BUFx3_ASAP7_75t_L g3177 ( 
.A(n_1987),
.Y(n_3177)
);

BUFx10_ASAP7_75t_L g3178 ( 
.A(n_1580),
.Y(n_3178)
);

CKINVDCx5p33_ASAP7_75t_R g3179 ( 
.A(n_278),
.Y(n_3179)
);

CKINVDCx5p33_ASAP7_75t_R g3180 ( 
.A(n_1653),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_675),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_1015),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2604),
.Y(n_3183)
);

CKINVDCx5p33_ASAP7_75t_R g3184 ( 
.A(n_2704),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_629),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_1170),
.Y(n_3186)
);

CKINVDCx5p33_ASAP7_75t_R g3187 ( 
.A(n_1332),
.Y(n_3187)
);

CKINVDCx16_ASAP7_75t_R g3188 ( 
.A(n_396),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_765),
.Y(n_3189)
);

INVx4_ASAP7_75t_R g3190 ( 
.A(n_2775),
.Y(n_3190)
);

CKINVDCx5p33_ASAP7_75t_R g3191 ( 
.A(n_2581),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_89),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_897),
.Y(n_3193)
);

CKINVDCx5p33_ASAP7_75t_R g3194 ( 
.A(n_2760),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_685),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_371),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2865),
.Y(n_3197)
);

CKINVDCx5p33_ASAP7_75t_R g3198 ( 
.A(n_2766),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_2480),
.Y(n_3199)
);

INVx1_ASAP7_75t_SL g3200 ( 
.A(n_1522),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_1552),
.Y(n_3201)
);

CKINVDCx20_ASAP7_75t_R g3202 ( 
.A(n_460),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_579),
.Y(n_3203)
);

CKINVDCx20_ASAP7_75t_R g3204 ( 
.A(n_2863),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_892),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_310),
.Y(n_3206)
);

CKINVDCx5p33_ASAP7_75t_R g3207 ( 
.A(n_388),
.Y(n_3207)
);

CKINVDCx5p33_ASAP7_75t_R g3208 ( 
.A(n_309),
.Y(n_3208)
);

CKINVDCx20_ASAP7_75t_R g3209 ( 
.A(n_188),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_1533),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_2867),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_2485),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_1367),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_432),
.Y(n_3214)
);

CKINVDCx20_ASAP7_75t_R g3215 ( 
.A(n_1991),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_1978),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_2054),
.Y(n_3217)
);

BUFx3_ASAP7_75t_L g3218 ( 
.A(n_872),
.Y(n_3218)
);

CKINVDCx16_ASAP7_75t_R g3219 ( 
.A(n_401),
.Y(n_3219)
);

BUFx10_ASAP7_75t_L g3220 ( 
.A(n_2038),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2708),
.Y(n_3221)
);

CKINVDCx5p33_ASAP7_75t_R g3222 ( 
.A(n_866),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_710),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_1523),
.Y(n_3224)
);

BUFx3_ASAP7_75t_L g3225 ( 
.A(n_2559),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_2896),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_150),
.Y(n_3227)
);

CKINVDCx5p33_ASAP7_75t_R g3228 ( 
.A(n_360),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2402),
.Y(n_3229)
);

INVxp67_ASAP7_75t_L g3230 ( 
.A(n_2274),
.Y(n_3230)
);

BUFx3_ASAP7_75t_L g3231 ( 
.A(n_1214),
.Y(n_3231)
);

CKINVDCx5p33_ASAP7_75t_R g3232 ( 
.A(n_1491),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_1498),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2730),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2463),
.Y(n_3235)
);

CKINVDCx5p33_ASAP7_75t_R g3236 ( 
.A(n_769),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_625),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_1642),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_2825),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_480),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_651),
.Y(n_3241)
);

CKINVDCx20_ASAP7_75t_R g3242 ( 
.A(n_1531),
.Y(n_3242)
);

CKINVDCx20_ASAP7_75t_R g3243 ( 
.A(n_313),
.Y(n_3243)
);

BUFx6f_ASAP7_75t_L g3244 ( 
.A(n_2806),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2582),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_2798),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_39),
.Y(n_3247)
);

CKINVDCx20_ASAP7_75t_R g3248 ( 
.A(n_2756),
.Y(n_3248)
);

CKINVDCx20_ASAP7_75t_R g3249 ( 
.A(n_2796),
.Y(n_3249)
);

BUFx3_ASAP7_75t_L g3250 ( 
.A(n_2734),
.Y(n_3250)
);

CKINVDCx5p33_ASAP7_75t_R g3251 ( 
.A(n_539),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_633),
.Y(n_3252)
);

CKINVDCx5p33_ASAP7_75t_R g3253 ( 
.A(n_173),
.Y(n_3253)
);

CKINVDCx5p33_ASAP7_75t_R g3254 ( 
.A(n_10),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2773),
.Y(n_3255)
);

CKINVDCx5p33_ASAP7_75t_R g3256 ( 
.A(n_2400),
.Y(n_3256)
);

CKINVDCx5p33_ASAP7_75t_R g3257 ( 
.A(n_688),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_1917),
.Y(n_3258)
);

CKINVDCx5p33_ASAP7_75t_R g3259 ( 
.A(n_1346),
.Y(n_3259)
);

CKINVDCx5p33_ASAP7_75t_R g3260 ( 
.A(n_2759),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_432),
.Y(n_3261)
);

BUFx8_ASAP7_75t_SL g3262 ( 
.A(n_2195),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_1242),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_1591),
.Y(n_3264)
);

BUFx8_ASAP7_75t_SL g3265 ( 
.A(n_1249),
.Y(n_3265)
);

BUFx3_ASAP7_75t_L g3266 ( 
.A(n_41),
.Y(n_3266)
);

CKINVDCx5p33_ASAP7_75t_R g3267 ( 
.A(n_2523),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_1358),
.Y(n_3268)
);

CKINVDCx5p33_ASAP7_75t_R g3269 ( 
.A(n_1278),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2535),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_1445),
.Y(n_3271)
);

CKINVDCx5p33_ASAP7_75t_R g3272 ( 
.A(n_1488),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_1297),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_1304),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_850),
.Y(n_3275)
);

CKINVDCx5p33_ASAP7_75t_R g3276 ( 
.A(n_960),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2357),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_719),
.Y(n_3278)
);

CKINVDCx20_ASAP7_75t_R g3279 ( 
.A(n_690),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2785),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_752),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_2792),
.Y(n_3282)
);

CKINVDCx5p33_ASAP7_75t_R g3283 ( 
.A(n_2284),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2749),
.Y(n_3284)
);

CKINVDCx5p33_ASAP7_75t_R g3285 ( 
.A(n_2795),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2216),
.Y(n_3286)
);

CKINVDCx5p33_ASAP7_75t_R g3287 ( 
.A(n_847),
.Y(n_3287)
);

CKINVDCx5p33_ASAP7_75t_R g3288 ( 
.A(n_2398),
.Y(n_3288)
);

CKINVDCx5p33_ASAP7_75t_R g3289 ( 
.A(n_2699),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_675),
.Y(n_3290)
);

CKINVDCx5p33_ASAP7_75t_R g3291 ( 
.A(n_733),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_2702),
.Y(n_3292)
);

BUFx10_ASAP7_75t_L g3293 ( 
.A(n_2771),
.Y(n_3293)
);

CKINVDCx5p33_ASAP7_75t_R g3294 ( 
.A(n_2755),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_1270),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_2100),
.Y(n_3296)
);

CKINVDCx5p33_ASAP7_75t_R g3297 ( 
.A(n_2325),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2754),
.Y(n_3298)
);

CKINVDCx5p33_ASAP7_75t_R g3299 ( 
.A(n_2712),
.Y(n_3299)
);

CKINVDCx14_ASAP7_75t_R g3300 ( 
.A(n_1452),
.Y(n_3300)
);

CKINVDCx5p33_ASAP7_75t_R g3301 ( 
.A(n_1234),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_792),
.Y(n_3302)
);

CKINVDCx5p33_ASAP7_75t_R g3303 ( 
.A(n_2607),
.Y(n_3303)
);

CKINVDCx5p33_ASAP7_75t_R g3304 ( 
.A(n_2782),
.Y(n_3304)
);

INVxp67_ASAP7_75t_L g3305 ( 
.A(n_2841),
.Y(n_3305)
);

CKINVDCx5p33_ASAP7_75t_R g3306 ( 
.A(n_2768),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_1809),
.Y(n_3307)
);

BUFx10_ASAP7_75t_L g3308 ( 
.A(n_2804),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_1779),
.Y(n_3309)
);

CKINVDCx5p33_ASAP7_75t_R g3310 ( 
.A(n_287),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_1201),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_451),
.Y(n_3312)
);

CKINVDCx5p33_ASAP7_75t_R g3313 ( 
.A(n_1967),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2582),
.Y(n_3314)
);

CKINVDCx5p33_ASAP7_75t_R g3315 ( 
.A(n_2767),
.Y(n_3315)
);

BUFx3_ASAP7_75t_L g3316 ( 
.A(n_2215),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2680),
.Y(n_3317)
);

CKINVDCx5p33_ASAP7_75t_R g3318 ( 
.A(n_395),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_13),
.Y(n_3319)
);

CKINVDCx20_ASAP7_75t_R g3320 ( 
.A(n_2011),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2002),
.Y(n_3321)
);

CKINVDCx20_ASAP7_75t_R g3322 ( 
.A(n_2589),
.Y(n_3322)
);

CKINVDCx20_ASAP7_75t_R g3323 ( 
.A(n_2407),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2791),
.Y(n_3324)
);

CKINVDCx5p33_ASAP7_75t_R g3325 ( 
.A(n_707),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2916),
.Y(n_3326)
);

CKINVDCx5p33_ASAP7_75t_R g3327 ( 
.A(n_1870),
.Y(n_3327)
);

CKINVDCx5p33_ASAP7_75t_R g3328 ( 
.A(n_884),
.Y(n_3328)
);

CKINVDCx5p33_ASAP7_75t_R g3329 ( 
.A(n_1691),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_215),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_31),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_346),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_10),
.Y(n_3333)
);

CKINVDCx5p33_ASAP7_75t_R g3334 ( 
.A(n_1783),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_2332),
.Y(n_3335)
);

CKINVDCx5p33_ASAP7_75t_R g3336 ( 
.A(n_249),
.Y(n_3336)
);

CKINVDCx5p33_ASAP7_75t_R g3337 ( 
.A(n_547),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2415),
.Y(n_3338)
);

CKINVDCx5p33_ASAP7_75t_R g3339 ( 
.A(n_1850),
.Y(n_3339)
);

CKINVDCx5p33_ASAP7_75t_R g3340 ( 
.A(n_2187),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_900),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_2746),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_1037),
.Y(n_3343)
);

CKINVDCx5p33_ASAP7_75t_R g3344 ( 
.A(n_2389),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_616),
.Y(n_3345)
);

CKINVDCx5p33_ASAP7_75t_R g3346 ( 
.A(n_320),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2002),
.Y(n_3347)
);

CKINVDCx5p33_ASAP7_75t_R g3348 ( 
.A(n_2442),
.Y(n_3348)
);

INVx2_ASAP7_75t_SL g3349 ( 
.A(n_1141),
.Y(n_3349)
);

HB1xp67_ASAP7_75t_L g3350 ( 
.A(n_1112),
.Y(n_3350)
);

CKINVDCx5p33_ASAP7_75t_R g3351 ( 
.A(n_1350),
.Y(n_3351)
);

CKINVDCx5p33_ASAP7_75t_R g3352 ( 
.A(n_2552),
.Y(n_3352)
);

INVx1_ASAP7_75t_SL g3353 ( 
.A(n_2738),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2472),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_368),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_897),
.Y(n_3356)
);

CKINVDCx14_ASAP7_75t_R g3357 ( 
.A(n_2434),
.Y(n_3357)
);

CKINVDCx5p33_ASAP7_75t_R g3358 ( 
.A(n_2753),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_1256),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2851),
.Y(n_3360)
);

CKINVDCx20_ASAP7_75t_R g3361 ( 
.A(n_721),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_1159),
.Y(n_3362)
);

CKINVDCx5p33_ASAP7_75t_R g3363 ( 
.A(n_1825),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_1534),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_33),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_1491),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_1792),
.Y(n_3367)
);

CKINVDCx5p33_ASAP7_75t_R g3368 ( 
.A(n_1156),
.Y(n_3368)
);

CKINVDCx5p33_ASAP7_75t_R g3369 ( 
.A(n_2718),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_2794),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2814),
.Y(n_3371)
);

CKINVDCx5p33_ASAP7_75t_R g3372 ( 
.A(n_2366),
.Y(n_3372)
);

CKINVDCx5p33_ASAP7_75t_R g3373 ( 
.A(n_2297),
.Y(n_3373)
);

CKINVDCx5p33_ASAP7_75t_R g3374 ( 
.A(n_2540),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2400),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2728),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_293),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2870),
.Y(n_3378)
);

BUFx8_ASAP7_75t_SL g3379 ( 
.A(n_1609),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_2142),
.Y(n_3380)
);

CKINVDCx5p33_ASAP7_75t_R g3381 ( 
.A(n_2732),
.Y(n_3381)
);

CKINVDCx5p33_ASAP7_75t_R g3382 ( 
.A(n_1218),
.Y(n_3382)
);

CKINVDCx5p33_ASAP7_75t_R g3383 ( 
.A(n_2122),
.Y(n_3383)
);

CKINVDCx5p33_ASAP7_75t_R g3384 ( 
.A(n_732),
.Y(n_3384)
);

CKINVDCx5p33_ASAP7_75t_R g3385 ( 
.A(n_1947),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2723),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2235),
.Y(n_3387)
);

CKINVDCx5p33_ASAP7_75t_R g3388 ( 
.A(n_1166),
.Y(n_3388)
);

INVxp67_ASAP7_75t_L g3389 ( 
.A(n_2681),
.Y(n_3389)
);

CKINVDCx5p33_ASAP7_75t_R g3390 ( 
.A(n_596),
.Y(n_3390)
);

CKINVDCx5p33_ASAP7_75t_R g3391 ( 
.A(n_2891),
.Y(n_3391)
);

CKINVDCx5p33_ASAP7_75t_R g3392 ( 
.A(n_1978),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_2112),
.Y(n_3393)
);

CKINVDCx5p33_ASAP7_75t_R g3394 ( 
.A(n_2821),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2667),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2862),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_2075),
.Y(n_3397)
);

CKINVDCx5p33_ASAP7_75t_R g3398 ( 
.A(n_1793),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_248),
.Y(n_3399)
);

CKINVDCx5p33_ASAP7_75t_R g3400 ( 
.A(n_2817),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2682),
.Y(n_3401)
);

CKINVDCx20_ASAP7_75t_R g3402 ( 
.A(n_967),
.Y(n_3402)
);

CKINVDCx5p33_ASAP7_75t_R g3403 ( 
.A(n_1905),
.Y(n_3403)
);

CKINVDCx5p33_ASAP7_75t_R g3404 ( 
.A(n_1171),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2072),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2096),
.Y(n_3406)
);

INVx1_ASAP7_75t_SL g3407 ( 
.A(n_2846),
.Y(n_3407)
);

INVx1_ASAP7_75t_SL g3408 ( 
.A(n_2135),
.Y(n_3408)
);

CKINVDCx5p33_ASAP7_75t_R g3409 ( 
.A(n_225),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_925),
.Y(n_3410)
);

CKINVDCx5p33_ASAP7_75t_R g3411 ( 
.A(n_516),
.Y(n_3411)
);

CKINVDCx5p33_ASAP7_75t_R g3412 ( 
.A(n_389),
.Y(n_3412)
);

CKINVDCx5p33_ASAP7_75t_R g3413 ( 
.A(n_729),
.Y(n_3413)
);

CKINVDCx5p33_ASAP7_75t_R g3414 ( 
.A(n_474),
.Y(n_3414)
);

BUFx3_ASAP7_75t_L g3415 ( 
.A(n_2820),
.Y(n_3415)
);

CKINVDCx5p33_ASAP7_75t_R g3416 ( 
.A(n_2268),
.Y(n_3416)
);

CKINVDCx5p33_ASAP7_75t_R g3417 ( 
.A(n_1701),
.Y(n_3417)
);

CKINVDCx5p33_ASAP7_75t_R g3418 ( 
.A(n_2776),
.Y(n_3418)
);

CKINVDCx5p33_ASAP7_75t_R g3419 ( 
.A(n_2764),
.Y(n_3419)
);

BUFx6f_ASAP7_75t_L g3420 ( 
.A(n_334),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_415),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2033),
.Y(n_3422)
);

CKINVDCx5p33_ASAP7_75t_R g3423 ( 
.A(n_578),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_2104),
.Y(n_3424)
);

CKINVDCx5p33_ASAP7_75t_R g3425 ( 
.A(n_1096),
.Y(n_3425)
);

CKINVDCx14_ASAP7_75t_R g3426 ( 
.A(n_2876),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2703),
.Y(n_3427)
);

BUFx10_ASAP7_75t_L g3428 ( 
.A(n_2787),
.Y(n_3428)
);

CKINVDCx5p33_ASAP7_75t_R g3429 ( 
.A(n_2140),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_428),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_365),
.Y(n_3431)
);

CKINVDCx5p33_ASAP7_75t_R g3432 ( 
.A(n_431),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_1266),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_2657),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_226),
.Y(n_3435)
);

CKINVDCx5p33_ASAP7_75t_R g3436 ( 
.A(n_2395),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2287),
.Y(n_3437)
);

CKINVDCx5p33_ASAP7_75t_R g3438 ( 
.A(n_1580),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_579),
.Y(n_3439)
);

CKINVDCx5p33_ASAP7_75t_R g3440 ( 
.A(n_542),
.Y(n_3440)
);

INVx1_ASAP7_75t_SL g3441 ( 
.A(n_981),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_1099),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_229),
.Y(n_3443)
);

BUFx3_ASAP7_75t_L g3444 ( 
.A(n_1265),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_5),
.Y(n_3445)
);

CKINVDCx5p33_ASAP7_75t_R g3446 ( 
.A(n_345),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_1160),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_1297),
.Y(n_3448)
);

CKINVDCx5p33_ASAP7_75t_R g3449 ( 
.A(n_1256),
.Y(n_3449)
);

CKINVDCx5p33_ASAP7_75t_R g3450 ( 
.A(n_1226),
.Y(n_3450)
);

CKINVDCx20_ASAP7_75t_R g3451 ( 
.A(n_2662),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_1613),
.Y(n_3452)
);

BUFx2_ASAP7_75t_L g3453 ( 
.A(n_291),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_786),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_348),
.Y(n_3455)
);

CKINVDCx5p33_ASAP7_75t_R g3456 ( 
.A(n_2738),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_674),
.Y(n_3457)
);

INVx2_ASAP7_75t_SL g3458 ( 
.A(n_1177),
.Y(n_3458)
);

BUFx3_ASAP7_75t_L g3459 ( 
.A(n_1677),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_2673),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_2780),
.Y(n_3461)
);

CKINVDCx20_ASAP7_75t_R g3462 ( 
.A(n_148),
.Y(n_3462)
);

CKINVDCx5p33_ASAP7_75t_R g3463 ( 
.A(n_637),
.Y(n_3463)
);

CKINVDCx5p33_ASAP7_75t_R g3464 ( 
.A(n_1758),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2599),
.Y(n_3465)
);

CKINVDCx5p33_ASAP7_75t_R g3466 ( 
.A(n_2609),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_2487),
.Y(n_3467)
);

BUFx6f_ASAP7_75t_L g3468 ( 
.A(n_2506),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_729),
.Y(n_3469)
);

BUFx3_ASAP7_75t_L g3470 ( 
.A(n_1942),
.Y(n_3470)
);

CKINVDCx5p33_ASAP7_75t_R g3471 ( 
.A(n_1240),
.Y(n_3471)
);

CKINVDCx5p33_ASAP7_75t_R g3472 ( 
.A(n_56),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_2524),
.Y(n_3473)
);

CKINVDCx20_ASAP7_75t_R g3474 ( 
.A(n_2869),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_2829),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_672),
.Y(n_3476)
);

CKINVDCx5p33_ASAP7_75t_R g3477 ( 
.A(n_1561),
.Y(n_3477)
);

CKINVDCx20_ASAP7_75t_R g3478 ( 
.A(n_1605),
.Y(n_3478)
);

BUFx3_ASAP7_75t_L g3479 ( 
.A(n_2394),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_866),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_2801),
.Y(n_3481)
);

CKINVDCx16_ASAP7_75t_R g3482 ( 
.A(n_2864),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_2747),
.Y(n_3483)
);

CKINVDCx5p33_ASAP7_75t_R g3484 ( 
.A(n_702),
.Y(n_3484)
);

BUFx3_ASAP7_75t_L g3485 ( 
.A(n_1010),
.Y(n_3485)
);

INVx1_ASAP7_75t_SL g3486 ( 
.A(n_928),
.Y(n_3486)
);

CKINVDCx5p33_ASAP7_75t_R g3487 ( 
.A(n_278),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_219),
.Y(n_3488)
);

BUFx10_ASAP7_75t_L g3489 ( 
.A(n_2855),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_1599),
.Y(n_3490)
);

CKINVDCx5p33_ASAP7_75t_R g3491 ( 
.A(n_474),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_699),
.Y(n_3492)
);

CKINVDCx5p33_ASAP7_75t_R g3493 ( 
.A(n_1975),
.Y(n_3493)
);

CKINVDCx20_ASAP7_75t_R g3494 ( 
.A(n_331),
.Y(n_3494)
);

CKINVDCx20_ASAP7_75t_R g3495 ( 
.A(n_2135),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_2672),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_1236),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_1182),
.Y(n_3498)
);

INVx2_ASAP7_75t_SL g3499 ( 
.A(n_546),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_2745),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_778),
.Y(n_3501)
);

CKINVDCx5p33_ASAP7_75t_R g3502 ( 
.A(n_2203),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_857),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_145),
.Y(n_3504)
);

CKINVDCx5p33_ASAP7_75t_R g3505 ( 
.A(n_2632),
.Y(n_3505)
);

CKINVDCx5p33_ASAP7_75t_R g3506 ( 
.A(n_1516),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_2805),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_1683),
.Y(n_3508)
);

BUFx10_ASAP7_75t_L g3509 ( 
.A(n_1467),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_1211),
.Y(n_3510)
);

CKINVDCx5p33_ASAP7_75t_R g3511 ( 
.A(n_1554),
.Y(n_3511)
);

CKINVDCx5p33_ASAP7_75t_R g3512 ( 
.A(n_2779),
.Y(n_3512)
);

CKINVDCx16_ASAP7_75t_R g3513 ( 
.A(n_969),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_2797),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_693),
.Y(n_3515)
);

CKINVDCx5p33_ASAP7_75t_R g3516 ( 
.A(n_2715),
.Y(n_3516)
);

CKINVDCx5p33_ASAP7_75t_R g3517 ( 
.A(n_2822),
.Y(n_3517)
);

CKINVDCx5p33_ASAP7_75t_R g3518 ( 
.A(n_2381),
.Y(n_3518)
);

BUFx10_ASAP7_75t_L g3519 ( 
.A(n_540),
.Y(n_3519)
);

CKINVDCx5p33_ASAP7_75t_R g3520 ( 
.A(n_724),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_280),
.Y(n_3521)
);

CKINVDCx5p33_ASAP7_75t_R g3522 ( 
.A(n_75),
.Y(n_3522)
);

BUFx5_ASAP7_75t_L g3523 ( 
.A(n_1172),
.Y(n_3523)
);

CKINVDCx5p33_ASAP7_75t_R g3524 ( 
.A(n_1529),
.Y(n_3524)
);

BUFx10_ASAP7_75t_L g3525 ( 
.A(n_2456),
.Y(n_3525)
);

BUFx10_ASAP7_75t_L g3526 ( 
.A(n_2711),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_2860),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_126),
.Y(n_3528)
);

CKINVDCx5p33_ASAP7_75t_R g3529 ( 
.A(n_2352),
.Y(n_3529)
);

CKINVDCx5p33_ASAP7_75t_R g3530 ( 
.A(n_1371),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2161),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_2404),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2676),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_92),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_2252),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_159),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_1956),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_563),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_294),
.Y(n_3539)
);

BUFx6f_ASAP7_75t_L g3540 ( 
.A(n_2770),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_1561),
.Y(n_3541)
);

CKINVDCx5p33_ASAP7_75t_R g3542 ( 
.A(n_827),
.Y(n_3542)
);

BUFx3_ASAP7_75t_L g3543 ( 
.A(n_1544),
.Y(n_3543)
);

CKINVDCx5p33_ASAP7_75t_R g3544 ( 
.A(n_1506),
.Y(n_3544)
);

CKINVDCx5p33_ASAP7_75t_R g3545 ( 
.A(n_822),
.Y(n_3545)
);

CKINVDCx5p33_ASAP7_75t_R g3546 ( 
.A(n_575),
.Y(n_3546)
);

BUFx10_ASAP7_75t_L g3547 ( 
.A(n_438),
.Y(n_3547)
);

CKINVDCx5p33_ASAP7_75t_R g3548 ( 
.A(n_2369),
.Y(n_3548)
);

CKINVDCx5p33_ASAP7_75t_R g3549 ( 
.A(n_2562),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_1791),
.Y(n_3550)
);

BUFx6f_ASAP7_75t_L g3551 ( 
.A(n_1688),
.Y(n_3551)
);

CKINVDCx5p33_ASAP7_75t_R g3552 ( 
.A(n_2329),
.Y(n_3552)
);

CKINVDCx5p33_ASAP7_75t_R g3553 ( 
.A(n_2521),
.Y(n_3553)
);

BUFx3_ASAP7_75t_L g3554 ( 
.A(n_2783),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_2224),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_1018),
.Y(n_3556)
);

CKINVDCx5p33_ASAP7_75t_R g3557 ( 
.A(n_2687),
.Y(n_3557)
);

CKINVDCx5p33_ASAP7_75t_R g3558 ( 
.A(n_516),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_2630),
.Y(n_3559)
);

CKINVDCx5p33_ASAP7_75t_R g3560 ( 
.A(n_235),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_1794),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_2170),
.Y(n_3562)
);

CKINVDCx5p33_ASAP7_75t_R g3563 ( 
.A(n_400),
.Y(n_3563)
);

CKINVDCx5p33_ASAP7_75t_R g3564 ( 
.A(n_2487),
.Y(n_3564)
);

CKINVDCx5p33_ASAP7_75t_R g3565 ( 
.A(n_1433),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2764),
.Y(n_3566)
);

BUFx2_ASAP7_75t_L g3567 ( 
.A(n_2735),
.Y(n_3567)
);

CKINVDCx5p33_ASAP7_75t_R g3568 ( 
.A(n_1358),
.Y(n_3568)
);

CKINVDCx5p33_ASAP7_75t_R g3569 ( 
.A(n_1051),
.Y(n_3569)
);

CKINVDCx5p33_ASAP7_75t_R g3570 ( 
.A(n_603),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_607),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_76),
.Y(n_3572)
);

INVx2_ASAP7_75t_SL g3573 ( 
.A(n_277),
.Y(n_3573)
);

CKINVDCx5p33_ASAP7_75t_R g3574 ( 
.A(n_1332),
.Y(n_3574)
);

CKINVDCx5p33_ASAP7_75t_R g3575 ( 
.A(n_2508),
.Y(n_3575)
);

CKINVDCx5p33_ASAP7_75t_R g3576 ( 
.A(n_2263),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_2111),
.Y(n_3577)
);

CKINVDCx5p33_ASAP7_75t_R g3578 ( 
.A(n_2736),
.Y(n_3578)
);

CKINVDCx20_ASAP7_75t_R g3579 ( 
.A(n_1632),
.Y(n_3579)
);

CKINVDCx5p33_ASAP7_75t_R g3580 ( 
.A(n_2847),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2412),
.Y(n_3581)
);

CKINVDCx5p33_ASAP7_75t_R g3582 ( 
.A(n_1117),
.Y(n_3582)
);

CKINVDCx20_ASAP7_75t_R g3583 ( 
.A(n_1792),
.Y(n_3583)
);

CKINVDCx5p33_ASAP7_75t_R g3584 ( 
.A(n_306),
.Y(n_3584)
);

CKINVDCx20_ASAP7_75t_R g3585 ( 
.A(n_849),
.Y(n_3585)
);

BUFx10_ASAP7_75t_L g3586 ( 
.A(n_139),
.Y(n_3586)
);

CKINVDCx5p33_ASAP7_75t_R g3587 ( 
.A(n_2136),
.Y(n_3587)
);

CKINVDCx5p33_ASAP7_75t_R g3588 ( 
.A(n_93),
.Y(n_3588)
);

CKINVDCx5p33_ASAP7_75t_R g3589 ( 
.A(n_251),
.Y(n_3589)
);

CKINVDCx5p33_ASAP7_75t_R g3590 ( 
.A(n_1604),
.Y(n_3590)
);

CKINVDCx5p33_ASAP7_75t_R g3591 ( 
.A(n_1205),
.Y(n_3591)
);

CKINVDCx5p33_ASAP7_75t_R g3592 ( 
.A(n_977),
.Y(n_3592)
);

CKINVDCx5p33_ASAP7_75t_R g3593 ( 
.A(n_100),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_2824),
.Y(n_3594)
);

CKINVDCx5p33_ASAP7_75t_R g3595 ( 
.A(n_1883),
.Y(n_3595)
);

CKINVDCx5p33_ASAP7_75t_R g3596 ( 
.A(n_923),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_2229),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2164),
.Y(n_3598)
);

CKINVDCx20_ASAP7_75t_R g3599 ( 
.A(n_1852),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_21),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2181),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_1818),
.Y(n_3602)
);

BUFx10_ASAP7_75t_L g3603 ( 
.A(n_1355),
.Y(n_3603)
);

CKINVDCx5p33_ASAP7_75t_R g3604 ( 
.A(n_946),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_2207),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_1090),
.Y(n_3606)
);

CKINVDCx5p33_ASAP7_75t_R g3607 ( 
.A(n_1307),
.Y(n_3607)
);

CKINVDCx5p33_ASAP7_75t_R g3608 ( 
.A(n_2570),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_2832),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_490),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_412),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_791),
.Y(n_3612)
);

CKINVDCx5p33_ASAP7_75t_R g3613 ( 
.A(n_2242),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_856),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_1819),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_2039),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_2852),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_2012),
.Y(n_3618)
);

CKINVDCx5p33_ASAP7_75t_R g3619 ( 
.A(n_1667),
.Y(n_3619)
);

CKINVDCx5p33_ASAP7_75t_R g3620 ( 
.A(n_2846),
.Y(n_3620)
);

CKINVDCx5p33_ASAP7_75t_R g3621 ( 
.A(n_2737),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_267),
.Y(n_3622)
);

CKINVDCx5p33_ASAP7_75t_R g3623 ( 
.A(n_2671),
.Y(n_3623)
);

CKINVDCx20_ASAP7_75t_R g3624 ( 
.A(n_1655),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_2364),
.Y(n_3625)
);

CKINVDCx20_ASAP7_75t_R g3626 ( 
.A(n_2407),
.Y(n_3626)
);

CKINVDCx5p33_ASAP7_75t_R g3627 ( 
.A(n_313),
.Y(n_3627)
);

CKINVDCx20_ASAP7_75t_R g3628 ( 
.A(n_2713),
.Y(n_3628)
);

CKINVDCx5p33_ASAP7_75t_R g3629 ( 
.A(n_2537),
.Y(n_3629)
);

BUFx3_ASAP7_75t_L g3630 ( 
.A(n_2388),
.Y(n_3630)
);

CKINVDCx5p33_ASAP7_75t_R g3631 ( 
.A(n_1087),
.Y(n_3631)
);

CKINVDCx5p33_ASAP7_75t_R g3632 ( 
.A(n_71),
.Y(n_3632)
);

CKINVDCx20_ASAP7_75t_R g3633 ( 
.A(n_1753),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_1161),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_424),
.Y(n_3635)
);

CKINVDCx20_ASAP7_75t_R g3636 ( 
.A(n_913),
.Y(n_3636)
);

INVx2_ASAP7_75t_SL g3637 ( 
.A(n_1546),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_413),
.Y(n_3638)
);

CKINVDCx5p33_ASAP7_75t_R g3639 ( 
.A(n_1601),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_2845),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_2808),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_2683),
.Y(n_3642)
);

CKINVDCx5p33_ASAP7_75t_R g3643 ( 
.A(n_259),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_2900),
.Y(n_3644)
);

CKINVDCx5p33_ASAP7_75t_R g3645 ( 
.A(n_275),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_2761),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_1619),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2624),
.Y(n_3648)
);

BUFx10_ASAP7_75t_L g3649 ( 
.A(n_130),
.Y(n_3649)
);

CKINVDCx20_ASAP7_75t_R g3650 ( 
.A(n_44),
.Y(n_3650)
);

CKINVDCx20_ASAP7_75t_R g3651 ( 
.A(n_197),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_764),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_2209),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_644),
.Y(n_3654)
);

CKINVDCx5p33_ASAP7_75t_R g3655 ( 
.A(n_2458),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_1441),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_885),
.Y(n_3657)
);

CKINVDCx5p33_ASAP7_75t_R g3658 ( 
.A(n_1872),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_1872),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_1236),
.Y(n_3660)
);

BUFx10_ASAP7_75t_L g3661 ( 
.A(n_1369),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_2727),
.Y(n_3662)
);

BUFx10_ASAP7_75t_L g3663 ( 
.A(n_2384),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_2064),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_1041),
.Y(n_3665)
);

CKINVDCx20_ASAP7_75t_R g3666 ( 
.A(n_874),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_2409),
.Y(n_3667)
);

CKINVDCx20_ASAP7_75t_R g3668 ( 
.A(n_353),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_1146),
.Y(n_3669)
);

CKINVDCx20_ASAP7_75t_R g3670 ( 
.A(n_1600),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_2235),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_621),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_1722),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2777),
.Y(n_3674)
);

CKINVDCx5p33_ASAP7_75t_R g3675 ( 
.A(n_488),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_19),
.Y(n_3676)
);

CKINVDCx5p33_ASAP7_75t_R g3677 ( 
.A(n_2710),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_2689),
.Y(n_3678)
);

CKINVDCx5p33_ASAP7_75t_R g3679 ( 
.A(n_2169),
.Y(n_3679)
);

BUFx6f_ASAP7_75t_L g3680 ( 
.A(n_2836),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_338),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_454),
.Y(n_3682)
);

CKINVDCx20_ASAP7_75t_R g3683 ( 
.A(n_402),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_2218),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_310),
.Y(n_3685)
);

CKINVDCx5p33_ASAP7_75t_R g3686 ( 
.A(n_2726),
.Y(n_3686)
);

CKINVDCx5p33_ASAP7_75t_R g3687 ( 
.A(n_2531),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_2816),
.Y(n_3688)
);

BUFx6f_ASAP7_75t_L g3689 ( 
.A(n_2494),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_2754),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_1975),
.Y(n_3691)
);

INVx2_ASAP7_75t_SL g3692 ( 
.A(n_2161),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_801),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_1670),
.Y(n_3694)
);

CKINVDCx20_ASAP7_75t_R g3695 ( 
.A(n_924),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_2694),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_1222),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_2060),
.Y(n_3698)
);

INVx1_ASAP7_75t_SL g3699 ( 
.A(n_1484),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_570),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_2148),
.Y(n_3701)
);

INVx2_ASAP7_75t_SL g3702 ( 
.A(n_2503),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_806),
.Y(n_3703)
);

CKINVDCx5p33_ASAP7_75t_R g3704 ( 
.A(n_2813),
.Y(n_3704)
);

INVx1_ASAP7_75t_SL g3705 ( 
.A(n_1188),
.Y(n_3705)
);

CKINVDCx5p33_ASAP7_75t_R g3706 ( 
.A(n_800),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_2301),
.Y(n_3707)
);

CKINVDCx5p33_ASAP7_75t_R g3708 ( 
.A(n_1487),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_307),
.Y(n_3709)
);

CKINVDCx5p33_ASAP7_75t_R g3710 ( 
.A(n_233),
.Y(n_3710)
);

CKINVDCx5p33_ASAP7_75t_R g3711 ( 
.A(n_770),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_2893),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_319),
.Y(n_3713)
);

CKINVDCx5p33_ASAP7_75t_R g3714 ( 
.A(n_961),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_1976),
.Y(n_3715)
);

CKINVDCx16_ASAP7_75t_R g3716 ( 
.A(n_2542),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_2669),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_2316),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_1326),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_1668),
.Y(n_3720)
);

CKINVDCx5p33_ASAP7_75t_R g3721 ( 
.A(n_517),
.Y(n_3721)
);

CKINVDCx5p33_ASAP7_75t_R g3722 ( 
.A(n_1775),
.Y(n_3722)
);

CKINVDCx5p33_ASAP7_75t_R g3723 ( 
.A(n_995),
.Y(n_3723)
);

CKINVDCx5p33_ASAP7_75t_R g3724 ( 
.A(n_1077),
.Y(n_3724)
);

CKINVDCx5p33_ASAP7_75t_R g3725 ( 
.A(n_2089),
.Y(n_3725)
);

CKINVDCx5p33_ASAP7_75t_R g3726 ( 
.A(n_2542),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_2872),
.Y(n_3727)
);

CKINVDCx20_ASAP7_75t_R g3728 ( 
.A(n_2719),
.Y(n_3728)
);

INVxp67_ASAP7_75t_SL g3729 ( 
.A(n_680),
.Y(n_3729)
);

CKINVDCx5p33_ASAP7_75t_R g3730 ( 
.A(n_856),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_1308),
.Y(n_3731)
);

CKINVDCx5p33_ASAP7_75t_R g3732 ( 
.A(n_138),
.Y(n_3732)
);

CKINVDCx5p33_ASAP7_75t_R g3733 ( 
.A(n_1221),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_1023),
.Y(n_3734)
);

CKINVDCx5p33_ASAP7_75t_R g3735 ( 
.A(n_1866),
.Y(n_3735)
);

CKINVDCx5p33_ASAP7_75t_R g3736 ( 
.A(n_2731),
.Y(n_3736)
);

CKINVDCx5p33_ASAP7_75t_R g3737 ( 
.A(n_2035),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_2858),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_1640),
.Y(n_3739)
);

CKINVDCx5p33_ASAP7_75t_R g3740 ( 
.A(n_2511),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_547),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_646),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_2741),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_644),
.Y(n_3744)
);

CKINVDCx5p33_ASAP7_75t_R g3745 ( 
.A(n_559),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_958),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_1869),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_1096),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_1475),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_2372),
.Y(n_3750)
);

BUFx10_ASAP7_75t_L g3751 ( 
.A(n_274),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_1753),
.Y(n_3752)
);

INVx1_ASAP7_75t_SL g3753 ( 
.A(n_2685),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_2430),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_2148),
.Y(n_3755)
);

CKINVDCx5p33_ASAP7_75t_R g3756 ( 
.A(n_2341),
.Y(n_3756)
);

CKINVDCx5p33_ASAP7_75t_R g3757 ( 
.A(n_2008),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_2696),
.Y(n_3758)
);

CKINVDCx5p33_ASAP7_75t_R g3759 ( 
.A(n_703),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_1448),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_2828),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_2747),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_2632),
.Y(n_3763)
);

CKINVDCx20_ASAP7_75t_R g3764 ( 
.A(n_2416),
.Y(n_3764)
);

CKINVDCx5p33_ASAP7_75t_R g3765 ( 
.A(n_2172),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_736),
.Y(n_3766)
);

CKINVDCx5p33_ASAP7_75t_R g3767 ( 
.A(n_1842),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_1537),
.Y(n_3768)
);

CKINVDCx5p33_ASAP7_75t_R g3769 ( 
.A(n_2442),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_273),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_2817),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_2087),
.Y(n_3772)
);

CKINVDCx5p33_ASAP7_75t_R g3773 ( 
.A(n_1938),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_1664),
.Y(n_3774)
);

CKINVDCx5p33_ASAP7_75t_R g3775 ( 
.A(n_2668),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_1648),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_40),
.Y(n_3777)
);

CKINVDCx20_ASAP7_75t_R g3778 ( 
.A(n_286),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_2877),
.Y(n_3779)
);

CKINVDCx5p33_ASAP7_75t_R g3780 ( 
.A(n_2390),
.Y(n_3780)
);

BUFx2_ASAP7_75t_L g3781 ( 
.A(n_341),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_317),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_265),
.Y(n_3783)
);

CKINVDCx5p33_ASAP7_75t_R g3784 ( 
.A(n_2528),
.Y(n_3784)
);

INVx2_ASAP7_75t_SL g3785 ( 
.A(n_1319),
.Y(n_3785)
);

INVx2_ASAP7_75t_SL g3786 ( 
.A(n_2417),
.Y(n_3786)
);

CKINVDCx5p33_ASAP7_75t_R g3787 ( 
.A(n_2805),
.Y(n_3787)
);

CKINVDCx5p33_ASAP7_75t_R g3788 ( 
.A(n_2264),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_2315),
.Y(n_3789)
);

CKINVDCx20_ASAP7_75t_R g3790 ( 
.A(n_2224),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_1919),
.Y(n_3791)
);

INVx1_ASAP7_75t_SL g3792 ( 
.A(n_989),
.Y(n_3792)
);

CKINVDCx20_ASAP7_75t_R g3793 ( 
.A(n_1406),
.Y(n_3793)
);

BUFx3_ASAP7_75t_L g3794 ( 
.A(n_107),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_1138),
.Y(n_3795)
);

CKINVDCx5p33_ASAP7_75t_R g3796 ( 
.A(n_2359),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_499),
.Y(n_3797)
);

HB1xp67_ASAP7_75t_L g3798 ( 
.A(n_2270),
.Y(n_3798)
);

CKINVDCx5p33_ASAP7_75t_R g3799 ( 
.A(n_2834),
.Y(n_3799)
);

INVx1_ASAP7_75t_SL g3800 ( 
.A(n_1890),
.Y(n_3800)
);

CKINVDCx5p33_ASAP7_75t_R g3801 ( 
.A(n_100),
.Y(n_3801)
);

INVx1_ASAP7_75t_SL g3802 ( 
.A(n_331),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_2151),
.Y(n_3803)
);

CKINVDCx5p33_ASAP7_75t_R g3804 ( 
.A(n_2608),
.Y(n_3804)
);

CKINVDCx5p33_ASAP7_75t_R g3805 ( 
.A(n_652),
.Y(n_3805)
);

CKINVDCx5p33_ASAP7_75t_R g3806 ( 
.A(n_2629),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_908),
.Y(n_3807)
);

CKINVDCx5p33_ASAP7_75t_R g3808 ( 
.A(n_2480),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_130),
.Y(n_3809)
);

CKINVDCx5p33_ASAP7_75t_R g3810 ( 
.A(n_2819),
.Y(n_3810)
);

CKINVDCx5p33_ASAP7_75t_R g3811 ( 
.A(n_1538),
.Y(n_3811)
);

CKINVDCx16_ASAP7_75t_R g3812 ( 
.A(n_1098),
.Y(n_3812)
);

CKINVDCx20_ASAP7_75t_R g3813 ( 
.A(n_2711),
.Y(n_3813)
);

CKINVDCx20_ASAP7_75t_R g3814 ( 
.A(n_2029),
.Y(n_3814)
);

CKINVDCx5p33_ASAP7_75t_R g3815 ( 
.A(n_1517),
.Y(n_3815)
);

CKINVDCx5p33_ASAP7_75t_R g3816 ( 
.A(n_1562),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_2774),
.Y(n_3817)
);

CKINVDCx5p33_ASAP7_75t_R g3818 ( 
.A(n_362),
.Y(n_3818)
);

CKINVDCx5p33_ASAP7_75t_R g3819 ( 
.A(n_439),
.Y(n_3819)
);

CKINVDCx5p33_ASAP7_75t_R g3820 ( 
.A(n_2275),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_2429),
.Y(n_3821)
);

CKINVDCx5p33_ASAP7_75t_R g3822 ( 
.A(n_10),
.Y(n_3822)
);

CKINVDCx5p33_ASAP7_75t_R g3823 ( 
.A(n_2695),
.Y(n_3823)
);

CKINVDCx5p33_ASAP7_75t_R g3824 ( 
.A(n_1008),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_959),
.Y(n_3825)
);

CKINVDCx5p33_ASAP7_75t_R g3826 ( 
.A(n_2857),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_697),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_1050),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_166),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_2716),
.Y(n_3830)
);

CKINVDCx16_ASAP7_75t_R g3831 ( 
.A(n_1198),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_2103),
.Y(n_3832)
);

CKINVDCx5p33_ASAP7_75t_R g3833 ( 
.A(n_2765),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_2818),
.Y(n_3834)
);

CKINVDCx5p33_ASAP7_75t_R g3835 ( 
.A(n_2639),
.Y(n_3835)
);

CKINVDCx5p33_ASAP7_75t_R g3836 ( 
.A(n_484),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_2538),
.Y(n_3837)
);

CKINVDCx5p33_ASAP7_75t_R g3838 ( 
.A(n_1509),
.Y(n_3838)
);

CKINVDCx5p33_ASAP7_75t_R g3839 ( 
.A(n_1238),
.Y(n_3839)
);

BUFx6f_ASAP7_75t_L g3840 ( 
.A(n_2786),
.Y(n_3840)
);

INVx1_ASAP7_75t_SL g3841 ( 
.A(n_132),
.Y(n_3841)
);

CKINVDCx5p33_ASAP7_75t_R g3842 ( 
.A(n_1352),
.Y(n_3842)
);

CKINVDCx5p33_ASAP7_75t_R g3843 ( 
.A(n_1483),
.Y(n_3843)
);

CKINVDCx5p33_ASAP7_75t_R g3844 ( 
.A(n_819),
.Y(n_3844)
);

BUFx6f_ASAP7_75t_L g3845 ( 
.A(n_92),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_2900),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_2053),
.Y(n_3847)
);

CKINVDCx5p33_ASAP7_75t_R g3848 ( 
.A(n_1750),
.Y(n_3848)
);

CKINVDCx5p33_ASAP7_75t_R g3849 ( 
.A(n_1013),
.Y(n_3849)
);

CKINVDCx5p33_ASAP7_75t_R g3850 ( 
.A(n_1783),
.Y(n_3850)
);

CKINVDCx5p33_ASAP7_75t_R g3851 ( 
.A(n_2298),
.Y(n_3851)
);

CKINVDCx5p33_ASAP7_75t_R g3852 ( 
.A(n_1162),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_2097),
.Y(n_3853)
);

CKINVDCx5p33_ASAP7_75t_R g3854 ( 
.A(n_1311),
.Y(n_3854)
);

CKINVDCx16_ASAP7_75t_R g3855 ( 
.A(n_1133),
.Y(n_3855)
);

CKINVDCx5p33_ASAP7_75t_R g3856 ( 
.A(n_368),
.Y(n_3856)
);

CKINVDCx20_ASAP7_75t_R g3857 ( 
.A(n_1737),
.Y(n_3857)
);

CKINVDCx20_ASAP7_75t_R g3858 ( 
.A(n_143),
.Y(n_3858)
);

CKINVDCx5p33_ASAP7_75t_R g3859 ( 
.A(n_1228),
.Y(n_3859)
);

BUFx6f_ASAP7_75t_L g3860 ( 
.A(n_1955),
.Y(n_3860)
);

BUFx2_ASAP7_75t_SL g3861 ( 
.A(n_278),
.Y(n_3861)
);

CKINVDCx5p33_ASAP7_75t_R g3862 ( 
.A(n_109),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_2007),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_1629),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_1904),
.Y(n_3865)
);

CKINVDCx5p33_ASAP7_75t_R g3866 ( 
.A(n_1842),
.Y(n_3866)
);

CKINVDCx5p33_ASAP7_75t_R g3867 ( 
.A(n_2848),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_624),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_2705),
.Y(n_3869)
);

CKINVDCx5p33_ASAP7_75t_R g3870 ( 
.A(n_1517),
.Y(n_3870)
);

CKINVDCx5p33_ASAP7_75t_R g3871 ( 
.A(n_2733),
.Y(n_3871)
);

CKINVDCx5p33_ASAP7_75t_R g3872 ( 
.A(n_133),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_2045),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_1823),
.Y(n_3874)
);

CKINVDCx5p33_ASAP7_75t_R g3875 ( 
.A(n_1327),
.Y(n_3875)
);

CKINVDCx5p33_ASAP7_75t_R g3876 ( 
.A(n_901),
.Y(n_3876)
);

CKINVDCx16_ASAP7_75t_R g3877 ( 
.A(n_2740),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_2850),
.Y(n_3878)
);

CKINVDCx5p33_ASAP7_75t_R g3879 ( 
.A(n_2793),
.Y(n_3879)
);

CKINVDCx20_ASAP7_75t_R g3880 ( 
.A(n_2541),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_2352),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_37),
.Y(n_3882)
);

CKINVDCx5p33_ASAP7_75t_R g3883 ( 
.A(n_2155),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_1214),
.Y(n_3884)
);

BUFx6f_ASAP7_75t_L g3885 ( 
.A(n_286),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_1728),
.Y(n_3886)
);

CKINVDCx5p33_ASAP7_75t_R g3887 ( 
.A(n_1311),
.Y(n_3887)
);

CKINVDCx5p33_ASAP7_75t_R g3888 ( 
.A(n_2046),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_896),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_527),
.Y(n_3890)
);

CKINVDCx5p33_ASAP7_75t_R g3891 ( 
.A(n_2677),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_2732),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_1288),
.Y(n_3893)
);

CKINVDCx20_ASAP7_75t_R g3894 ( 
.A(n_410),
.Y(n_3894)
);

CKINVDCx5p33_ASAP7_75t_R g3895 ( 
.A(n_1157),
.Y(n_3895)
);

CKINVDCx5p33_ASAP7_75t_R g3896 ( 
.A(n_1097),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_723),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_2844),
.Y(n_3898)
);

CKINVDCx5p33_ASAP7_75t_R g3899 ( 
.A(n_181),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_1684),
.Y(n_3900)
);

CKINVDCx5p33_ASAP7_75t_R g3901 ( 
.A(n_227),
.Y(n_3901)
);

BUFx10_ASAP7_75t_L g3902 ( 
.A(n_829),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_2434),
.Y(n_3903)
);

CKINVDCx5p33_ASAP7_75t_R g3904 ( 
.A(n_2830),
.Y(n_3904)
);

CKINVDCx5p33_ASAP7_75t_R g3905 ( 
.A(n_2801),
.Y(n_3905)
);

CKINVDCx5p33_ASAP7_75t_R g3906 ( 
.A(n_19),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_295),
.Y(n_3907)
);

CKINVDCx5p33_ASAP7_75t_R g3908 ( 
.A(n_1784),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_2562),
.Y(n_3909)
);

CKINVDCx20_ASAP7_75t_R g3910 ( 
.A(n_2698),
.Y(n_3910)
);

CKINVDCx5p33_ASAP7_75t_R g3911 ( 
.A(n_1803),
.Y(n_3911)
);

BUFx6f_ASAP7_75t_L g3912 ( 
.A(n_850),
.Y(n_3912)
);

INVx1_ASAP7_75t_SL g3913 ( 
.A(n_1069),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_1869),
.Y(n_3914)
);

CKINVDCx5p33_ASAP7_75t_R g3915 ( 
.A(n_1905),
.Y(n_3915)
);

CKINVDCx5p33_ASAP7_75t_R g3916 ( 
.A(n_864),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_1334),
.Y(n_3917)
);

CKINVDCx20_ASAP7_75t_R g3918 ( 
.A(n_1068),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_247),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_193),
.Y(n_3920)
);

CKINVDCx16_ASAP7_75t_R g3921 ( 
.A(n_2799),
.Y(n_3921)
);

BUFx8_ASAP7_75t_SL g3922 ( 
.A(n_1889),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_2809),
.Y(n_3923)
);

CKINVDCx5p33_ASAP7_75t_R g3924 ( 
.A(n_1356),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_2781),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_2232),
.Y(n_3926)
);

BUFx3_ASAP7_75t_L g3927 ( 
.A(n_2724),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_528),
.Y(n_3928)
);

CKINVDCx5p33_ASAP7_75t_R g3929 ( 
.A(n_2810),
.Y(n_3929)
);

CKINVDCx5p33_ASAP7_75t_R g3930 ( 
.A(n_2717),
.Y(n_3930)
);

CKINVDCx20_ASAP7_75t_R g3931 ( 
.A(n_1008),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_222),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_2646),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_2038),
.Y(n_3934)
);

CKINVDCx5p33_ASAP7_75t_R g3935 ( 
.A(n_355),
.Y(n_3935)
);

CKINVDCx5p33_ASAP7_75t_R g3936 ( 
.A(n_1239),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_1089),
.Y(n_3937)
);

CKINVDCx5p33_ASAP7_75t_R g3938 ( 
.A(n_1471),
.Y(n_3938)
);

BUFx6f_ASAP7_75t_L g3939 ( 
.A(n_1032),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_2859),
.Y(n_3940)
);

BUFx6f_ASAP7_75t_L g3941 ( 
.A(n_975),
.Y(n_3941)
);

CKINVDCx5p33_ASAP7_75t_R g3942 ( 
.A(n_2047),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_931),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_2750),
.Y(n_3944)
);

CKINVDCx5p33_ASAP7_75t_R g3945 ( 
.A(n_2440),
.Y(n_3945)
);

CKINVDCx5p33_ASAP7_75t_R g3946 ( 
.A(n_71),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_1981),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_1420),
.Y(n_3948)
);

CKINVDCx5p33_ASAP7_75t_R g3949 ( 
.A(n_429),
.Y(n_3949)
);

CKINVDCx5p33_ASAP7_75t_R g3950 ( 
.A(n_2124),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_1299),
.Y(n_3951)
);

CKINVDCx5p33_ASAP7_75t_R g3952 ( 
.A(n_1965),
.Y(n_3952)
);

CKINVDCx5p33_ASAP7_75t_R g3953 ( 
.A(n_1949),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_2829),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_2665),
.Y(n_3955)
);

CKINVDCx20_ASAP7_75t_R g3956 ( 
.A(n_1292),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_130),
.Y(n_3957)
);

INVx1_ASAP7_75t_SL g3958 ( 
.A(n_1338),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_1374),
.Y(n_3959)
);

CKINVDCx5p33_ASAP7_75t_R g3960 ( 
.A(n_1588),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_2563),
.Y(n_3961)
);

CKINVDCx5p33_ASAP7_75t_R g3962 ( 
.A(n_2623),
.Y(n_3962)
);

CKINVDCx5p33_ASAP7_75t_R g3963 ( 
.A(n_1801),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_976),
.Y(n_3964)
);

BUFx2_ASAP7_75t_L g3965 ( 
.A(n_2790),
.Y(n_3965)
);

INVx1_ASAP7_75t_SL g3966 ( 
.A(n_1402),
.Y(n_3966)
);

CKINVDCx5p33_ASAP7_75t_R g3967 ( 
.A(n_973),
.Y(n_3967)
);

CKINVDCx5p33_ASAP7_75t_R g3968 ( 
.A(n_1254),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_836),
.Y(n_3969)
);

CKINVDCx5p33_ASAP7_75t_R g3970 ( 
.A(n_869),
.Y(n_3970)
);

CKINVDCx5p33_ASAP7_75t_R g3971 ( 
.A(n_1562),
.Y(n_3971)
);

CKINVDCx5p33_ASAP7_75t_R g3972 ( 
.A(n_329),
.Y(n_3972)
);

CKINVDCx20_ASAP7_75t_R g3973 ( 
.A(n_1739),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_256),
.Y(n_3974)
);

BUFx8_ASAP7_75t_SL g3975 ( 
.A(n_2187),
.Y(n_3975)
);

CKINVDCx5p33_ASAP7_75t_R g3976 ( 
.A(n_2745),
.Y(n_3976)
);

CKINVDCx5p33_ASAP7_75t_R g3977 ( 
.A(n_1887),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_605),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_41),
.Y(n_3979)
);

CKINVDCx20_ASAP7_75t_R g3980 ( 
.A(n_931),
.Y(n_3980)
);

CKINVDCx5p33_ASAP7_75t_R g3981 ( 
.A(n_60),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_2194),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_257),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_2501),
.Y(n_3984)
);

CKINVDCx20_ASAP7_75t_R g3985 ( 
.A(n_2868),
.Y(n_3985)
);

BUFx10_ASAP7_75t_L g3986 ( 
.A(n_2775),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_2739),
.Y(n_3987)
);

CKINVDCx20_ASAP7_75t_R g3988 ( 
.A(n_879),
.Y(n_3988)
);

CKINVDCx5p33_ASAP7_75t_R g3989 ( 
.A(n_1974),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_393),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_2131),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_613),
.Y(n_3992)
);

BUFx2_ASAP7_75t_L g3993 ( 
.A(n_2315),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_2878),
.Y(n_3994)
);

CKINVDCx5p33_ASAP7_75t_R g3995 ( 
.A(n_2868),
.Y(n_3995)
);

BUFx3_ASAP7_75t_L g3996 ( 
.A(n_1919),
.Y(n_3996)
);

HB1xp67_ASAP7_75t_L g3997 ( 
.A(n_952),
.Y(n_3997)
);

CKINVDCx5p33_ASAP7_75t_R g3998 ( 
.A(n_881),
.Y(n_3998)
);

BUFx6f_ASAP7_75t_L g3999 ( 
.A(n_194),
.Y(n_3999)
);

BUFx8_ASAP7_75t_SL g4000 ( 
.A(n_445),
.Y(n_4000)
);

CKINVDCx5p33_ASAP7_75t_R g4001 ( 
.A(n_185),
.Y(n_4001)
);

CKINVDCx5p33_ASAP7_75t_R g4002 ( 
.A(n_1899),
.Y(n_4002)
);

CKINVDCx5p33_ASAP7_75t_R g4003 ( 
.A(n_1286),
.Y(n_4003)
);

CKINVDCx5p33_ASAP7_75t_R g4004 ( 
.A(n_89),
.Y(n_4004)
);

CKINVDCx20_ASAP7_75t_R g4005 ( 
.A(n_1162),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_1141),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_2714),
.Y(n_4007)
);

CKINVDCx5p33_ASAP7_75t_R g4008 ( 
.A(n_980),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_269),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_302),
.Y(n_4010)
);

INVx1_ASAP7_75t_SL g4011 ( 
.A(n_1844),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_2910),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_2116),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_2040),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_2719),
.Y(n_4015)
);

CKINVDCx5p33_ASAP7_75t_R g4016 ( 
.A(n_804),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_2359),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_1515),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_2842),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_1053),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_1336),
.Y(n_4021)
);

CKINVDCx5p33_ASAP7_75t_R g4022 ( 
.A(n_1351),
.Y(n_4022)
);

CKINVDCx5p33_ASAP7_75t_R g4023 ( 
.A(n_2706),
.Y(n_4023)
);

INVx2_ASAP7_75t_L g4024 ( 
.A(n_550),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_2714),
.Y(n_4025)
);

BUFx6f_ASAP7_75t_L g4026 ( 
.A(n_2556),
.Y(n_4026)
);

CKINVDCx5p33_ASAP7_75t_R g4027 ( 
.A(n_247),
.Y(n_4027)
);

CKINVDCx5p33_ASAP7_75t_R g4028 ( 
.A(n_2089),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_1779),
.Y(n_4029)
);

CKINVDCx5p33_ASAP7_75t_R g4030 ( 
.A(n_128),
.Y(n_4030)
);

CKINVDCx5p33_ASAP7_75t_R g4031 ( 
.A(n_2839),
.Y(n_4031)
);

CKINVDCx5p33_ASAP7_75t_R g4032 ( 
.A(n_463),
.Y(n_4032)
);

CKINVDCx5p33_ASAP7_75t_R g4033 ( 
.A(n_2650),
.Y(n_4033)
);

CKINVDCx5p33_ASAP7_75t_R g4034 ( 
.A(n_778),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_907),
.Y(n_4035)
);

CKINVDCx5p33_ASAP7_75t_R g4036 ( 
.A(n_1320),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_2595),
.Y(n_4037)
);

HB1xp67_ASAP7_75t_L g4038 ( 
.A(n_1224),
.Y(n_4038)
);

CKINVDCx5p33_ASAP7_75t_R g4039 ( 
.A(n_667),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_786),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_2085),
.Y(n_4041)
);

BUFx6f_ASAP7_75t_L g4042 ( 
.A(n_2043),
.Y(n_4042)
);

INVx1_ASAP7_75t_SL g4043 ( 
.A(n_1478),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_2139),
.Y(n_4044)
);

CKINVDCx5p33_ASAP7_75t_R g4045 ( 
.A(n_561),
.Y(n_4045)
);

CKINVDCx20_ASAP7_75t_R g4046 ( 
.A(n_305),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_1453),
.Y(n_4047)
);

CKINVDCx5p33_ASAP7_75t_R g4048 ( 
.A(n_2545),
.Y(n_4048)
);

INVx2_ASAP7_75t_SL g4049 ( 
.A(n_769),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_441),
.Y(n_4050)
);

INVx2_ASAP7_75t_SL g4051 ( 
.A(n_1028),
.Y(n_4051)
);

CKINVDCx5p33_ASAP7_75t_R g4052 ( 
.A(n_2789),
.Y(n_4052)
);

INVxp67_ASAP7_75t_SL g4053 ( 
.A(n_171),
.Y(n_4053)
);

BUFx3_ASAP7_75t_L g4054 ( 
.A(n_2837),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_1548),
.Y(n_4055)
);

CKINVDCx5p33_ASAP7_75t_R g4056 ( 
.A(n_2835),
.Y(n_4056)
);

BUFx2_ASAP7_75t_L g4057 ( 
.A(n_686),
.Y(n_4057)
);

CKINVDCx5p33_ASAP7_75t_R g4058 ( 
.A(n_717),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_1230),
.Y(n_4059)
);

CKINVDCx5p33_ASAP7_75t_R g4060 ( 
.A(n_2172),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_2691),
.Y(n_4061)
);

CKINVDCx5p33_ASAP7_75t_R g4062 ( 
.A(n_2472),
.Y(n_4062)
);

CKINVDCx5p33_ASAP7_75t_R g4063 ( 
.A(n_2721),
.Y(n_4063)
);

CKINVDCx5p33_ASAP7_75t_R g4064 ( 
.A(n_259),
.Y(n_4064)
);

CKINVDCx20_ASAP7_75t_R g4065 ( 
.A(n_1767),
.Y(n_4065)
);

BUFx3_ASAP7_75t_L g4066 ( 
.A(n_1124),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_1403),
.Y(n_4067)
);

CKINVDCx20_ASAP7_75t_R g4068 ( 
.A(n_511),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_1472),
.Y(n_4069)
);

CKINVDCx20_ASAP7_75t_R g4070 ( 
.A(n_1421),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_2749),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_553),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_224),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_60),
.Y(n_4074)
);

CKINVDCx14_ASAP7_75t_R g4075 ( 
.A(n_933),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_595),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_732),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_711),
.Y(n_4078)
);

BUFx2_ASAP7_75t_L g4079 ( 
.A(n_895),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_1742),
.Y(n_4080)
);

CKINVDCx5p33_ASAP7_75t_R g4081 ( 
.A(n_761),
.Y(n_4081)
);

BUFx6f_ASAP7_75t_L g4082 ( 
.A(n_365),
.Y(n_4082)
);

CKINVDCx5p33_ASAP7_75t_R g4083 ( 
.A(n_1220),
.Y(n_4083)
);

BUFx6f_ASAP7_75t_L g4084 ( 
.A(n_1448),
.Y(n_4084)
);

CKINVDCx5p33_ASAP7_75t_R g4085 ( 
.A(n_2140),
.Y(n_4085)
);

CKINVDCx5p33_ASAP7_75t_R g4086 ( 
.A(n_2688),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_2757),
.Y(n_4087)
);

CKINVDCx20_ASAP7_75t_R g4088 ( 
.A(n_2449),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_126),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_2199),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_2811),
.Y(n_4091)
);

INVxp67_ASAP7_75t_L g4092 ( 
.A(n_339),
.Y(n_4092)
);

CKINVDCx5p33_ASAP7_75t_R g4093 ( 
.A(n_1760),
.Y(n_4093)
);

CKINVDCx5p33_ASAP7_75t_R g4094 ( 
.A(n_519),
.Y(n_4094)
);

BUFx6f_ASAP7_75t_L g4095 ( 
.A(n_131),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_2815),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_414),
.Y(n_4097)
);

CKINVDCx5p33_ASAP7_75t_R g4098 ( 
.A(n_338),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_1553),
.Y(n_4099)
);

CKINVDCx5p33_ASAP7_75t_R g4100 ( 
.A(n_2763),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_1199),
.Y(n_4101)
);

CKINVDCx5p33_ASAP7_75t_R g4102 ( 
.A(n_2046),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_62),
.Y(n_4103)
);

CKINVDCx5p33_ASAP7_75t_R g4104 ( 
.A(n_1870),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_1762),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_1644),
.Y(n_4106)
);

CKINVDCx5p33_ASAP7_75t_R g4107 ( 
.A(n_2559),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_2769),
.Y(n_4108)
);

INVx3_ASAP7_75t_L g4109 ( 
.A(n_2458),
.Y(n_4109)
);

CKINVDCx5p33_ASAP7_75t_R g4110 ( 
.A(n_2209),
.Y(n_4110)
);

BUFx2_ASAP7_75t_L g4111 ( 
.A(n_1483),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_2636),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_2427),
.Y(n_4113)
);

CKINVDCx5p33_ASAP7_75t_R g4114 ( 
.A(n_766),
.Y(n_4114)
);

INVx1_ASAP7_75t_SL g4115 ( 
.A(n_957),
.Y(n_4115)
);

CKINVDCx20_ASAP7_75t_R g4116 ( 
.A(n_2405),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_880),
.Y(n_4117)
);

CKINVDCx5p33_ASAP7_75t_R g4118 ( 
.A(n_2331),
.Y(n_4118)
);

HB1xp67_ASAP7_75t_L g4119 ( 
.A(n_1498),
.Y(n_4119)
);

BUFx10_ASAP7_75t_L g4120 ( 
.A(n_1903),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_2523),
.Y(n_4121)
);

CKINVDCx5p33_ASAP7_75t_R g4122 ( 
.A(n_2778),
.Y(n_4122)
);

CKINVDCx14_ASAP7_75t_R g4123 ( 
.A(n_2590),
.Y(n_4123)
);

INVxp67_ASAP7_75t_SL g4124 ( 
.A(n_1120),
.Y(n_4124)
);

CKINVDCx5p33_ASAP7_75t_R g4125 ( 
.A(n_1211),
.Y(n_4125)
);

CKINVDCx5p33_ASAP7_75t_R g4126 ( 
.A(n_2693),
.Y(n_4126)
);

CKINVDCx5p33_ASAP7_75t_R g4127 ( 
.A(n_2412),
.Y(n_4127)
);

CKINVDCx5p33_ASAP7_75t_R g4128 ( 
.A(n_1154),
.Y(n_4128)
);

CKINVDCx5p33_ASAP7_75t_R g4129 ( 
.A(n_483),
.Y(n_4129)
);

CKINVDCx20_ASAP7_75t_R g4130 ( 
.A(n_2507),
.Y(n_4130)
);

INVx1_ASAP7_75t_SL g4131 ( 
.A(n_2335),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_1993),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_2679),
.Y(n_4133)
);

INVx2_ASAP7_75t_SL g4134 ( 
.A(n_2051),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_2826),
.Y(n_4135)
);

CKINVDCx5p33_ASAP7_75t_R g4136 ( 
.A(n_391),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_2301),
.Y(n_4137)
);

CKINVDCx20_ASAP7_75t_R g4138 ( 
.A(n_21),
.Y(n_4138)
);

INVx2_ASAP7_75t_SL g4139 ( 
.A(n_2617),
.Y(n_4139)
);

CKINVDCx5p33_ASAP7_75t_R g4140 ( 
.A(n_2429),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_595),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_1177),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_1832),
.Y(n_4143)
);

CKINVDCx20_ASAP7_75t_R g4144 ( 
.A(n_1074),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_2259),
.Y(n_4145)
);

CKINVDCx5p33_ASAP7_75t_R g4146 ( 
.A(n_1270),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_698),
.Y(n_4147)
);

CKINVDCx5p33_ASAP7_75t_R g4148 ( 
.A(n_1509),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_458),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_1800),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_1274),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_1252),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_1914),
.Y(n_4153)
);

CKINVDCx20_ASAP7_75t_R g4154 ( 
.A(n_1323),
.Y(n_4154)
);

CKINVDCx5p33_ASAP7_75t_R g4155 ( 
.A(n_1455),
.Y(n_4155)
);

CKINVDCx14_ASAP7_75t_R g4156 ( 
.A(n_2796),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_1861),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_900),
.Y(n_4158)
);

BUFx10_ASAP7_75t_L g4159 ( 
.A(n_109),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_2132),
.Y(n_4160)
);

CKINVDCx5p33_ASAP7_75t_R g4161 ( 
.A(n_957),
.Y(n_4161)
);

CKINVDCx5p33_ASAP7_75t_R g4162 ( 
.A(n_2678),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_2700),
.Y(n_4163)
);

INVx1_ASAP7_75t_SL g4164 ( 
.A(n_29),
.Y(n_4164)
);

BUFx8_ASAP7_75t_SL g4165 ( 
.A(n_2322),
.Y(n_4165)
);

CKINVDCx20_ASAP7_75t_R g4166 ( 
.A(n_2634),
.Y(n_4166)
);

CKINVDCx20_ASAP7_75t_R g4167 ( 
.A(n_2033),
.Y(n_4167)
);

CKINVDCx5p33_ASAP7_75t_R g4168 ( 
.A(n_1179),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_1663),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_2800),
.Y(n_4170)
);

CKINVDCx5p33_ASAP7_75t_R g4171 ( 
.A(n_2109),
.Y(n_4171)
);

CKINVDCx5p33_ASAP7_75t_R g4172 ( 
.A(n_464),
.Y(n_4172)
);

CKINVDCx5p33_ASAP7_75t_R g4173 ( 
.A(n_880),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_467),
.Y(n_4174)
);

CKINVDCx20_ASAP7_75t_R g4175 ( 
.A(n_2366),
.Y(n_4175)
);

CKINVDCx5p33_ASAP7_75t_R g4176 ( 
.A(n_506),
.Y(n_4176)
);

CKINVDCx5p33_ASAP7_75t_R g4177 ( 
.A(n_2239),
.Y(n_4177)
);

CKINVDCx5p33_ASAP7_75t_R g4178 ( 
.A(n_469),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_603),
.Y(n_4179)
);

INVx1_ASAP7_75t_SL g4180 ( 
.A(n_493),
.Y(n_4180)
);

CKINVDCx5p33_ASAP7_75t_R g4181 ( 
.A(n_2840),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_2309),
.Y(n_4182)
);

CKINVDCx20_ASAP7_75t_R g4183 ( 
.A(n_860),
.Y(n_4183)
);

CKINVDCx5p33_ASAP7_75t_R g4184 ( 
.A(n_468),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_74),
.Y(n_4185)
);

CKINVDCx20_ASAP7_75t_R g4186 ( 
.A(n_2608),
.Y(n_4186)
);

BUFx6f_ASAP7_75t_L g4187 ( 
.A(n_2814),
.Y(n_4187)
);

CKINVDCx5p33_ASAP7_75t_R g4188 ( 
.A(n_1196),
.Y(n_4188)
);

CKINVDCx20_ASAP7_75t_R g4189 ( 
.A(n_2099),
.Y(n_4189)
);

CKINVDCx5p33_ASAP7_75t_R g4190 ( 
.A(n_199),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_739),
.Y(n_4191)
);

CKINVDCx5p33_ASAP7_75t_R g4192 ( 
.A(n_982),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_670),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_609),
.Y(n_4194)
);

CKINVDCx5p33_ASAP7_75t_R g4195 ( 
.A(n_843),
.Y(n_4195)
);

CKINVDCx5p33_ASAP7_75t_R g4196 ( 
.A(n_2126),
.Y(n_4196)
);

CKINVDCx5p33_ASAP7_75t_R g4197 ( 
.A(n_1295),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_784),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_1742),
.Y(n_4199)
);

INVx2_ASAP7_75t_SL g4200 ( 
.A(n_2280),
.Y(n_4200)
);

BUFx3_ASAP7_75t_L g4201 ( 
.A(n_2433),
.Y(n_4201)
);

CKINVDCx5p33_ASAP7_75t_R g4202 ( 
.A(n_2751),
.Y(n_4202)
);

CKINVDCx5p33_ASAP7_75t_R g4203 ( 
.A(n_770),
.Y(n_4203)
);

CKINVDCx5p33_ASAP7_75t_R g4204 ( 
.A(n_294),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_1903),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_1576),
.Y(n_4206)
);

CKINVDCx5p33_ASAP7_75t_R g4207 ( 
.A(n_2681),
.Y(n_4207)
);

CKINVDCx5p33_ASAP7_75t_R g4208 ( 
.A(n_1997),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_1111),
.Y(n_4209)
);

CKINVDCx5p33_ASAP7_75t_R g4210 ( 
.A(n_1840),
.Y(n_4210)
);

CKINVDCx5p33_ASAP7_75t_R g4211 ( 
.A(n_2853),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_1831),
.Y(n_4212)
);

CKINVDCx5p33_ASAP7_75t_R g4213 ( 
.A(n_784),
.Y(n_4213)
);

CKINVDCx5p33_ASAP7_75t_R g4214 ( 
.A(n_631),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_916),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_2214),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_794),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_1070),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_548),
.Y(n_4219)
);

CKINVDCx5p33_ASAP7_75t_R g4220 ( 
.A(n_2709),
.Y(n_4220)
);

CKINVDCx5p33_ASAP7_75t_R g4221 ( 
.A(n_1412),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_2621),
.Y(n_4222)
);

CKINVDCx5p33_ASAP7_75t_R g4223 ( 
.A(n_88),
.Y(n_4223)
);

CKINVDCx5p33_ASAP7_75t_R g4224 ( 
.A(n_147),
.Y(n_4224)
);

CKINVDCx20_ASAP7_75t_R g4225 ( 
.A(n_1135),
.Y(n_4225)
);

CKINVDCx5p33_ASAP7_75t_R g4226 ( 
.A(n_2501),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_1345),
.Y(n_4227)
);

BUFx8_ASAP7_75t_SL g4228 ( 
.A(n_273),
.Y(n_4228)
);

CKINVDCx20_ASAP7_75t_R g4229 ( 
.A(n_2722),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_235),
.Y(n_4230)
);

CKINVDCx20_ASAP7_75t_R g4231 ( 
.A(n_1895),
.Y(n_4231)
);

BUFx6f_ASAP7_75t_L g4232 ( 
.A(n_2563),
.Y(n_4232)
);

INVxp67_ASAP7_75t_L g4233 ( 
.A(n_1522),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_2865),
.Y(n_4234)
);

CKINVDCx5p33_ASAP7_75t_R g4235 ( 
.A(n_701),
.Y(n_4235)
);

INVxp67_ASAP7_75t_L g4236 ( 
.A(n_292),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_801),
.Y(n_4237)
);

BUFx3_ASAP7_75t_L g4238 ( 
.A(n_176),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_2242),
.Y(n_4239)
);

CKINVDCx5p33_ASAP7_75t_R g4240 ( 
.A(n_1687),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_1821),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_857),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_1291),
.Y(n_4243)
);

CKINVDCx20_ASAP7_75t_R g4244 ( 
.A(n_2063),
.Y(n_4244)
);

CKINVDCx5p33_ASAP7_75t_R g4245 ( 
.A(n_2385),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_1915),
.Y(n_4246)
);

CKINVDCx20_ASAP7_75t_R g4247 ( 
.A(n_80),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_2762),
.Y(n_4248)
);

CKINVDCx20_ASAP7_75t_R g4249 ( 
.A(n_1135),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_283),
.Y(n_4250)
);

CKINVDCx5p33_ASAP7_75t_R g4251 ( 
.A(n_2305),
.Y(n_4251)
);

CKINVDCx20_ASAP7_75t_R g4252 ( 
.A(n_2870),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_624),
.Y(n_4253)
);

CKINVDCx5p33_ASAP7_75t_R g4254 ( 
.A(n_1885),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_89),
.Y(n_4255)
);

CKINVDCx5p33_ASAP7_75t_R g4256 ( 
.A(n_1991),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_2691),
.Y(n_4257)
);

CKINVDCx5p33_ASAP7_75t_R g4258 ( 
.A(n_2701),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_1988),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_1029),
.Y(n_4260)
);

INVx1_ASAP7_75t_SL g4261 ( 
.A(n_1389),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_1053),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_2035),
.Y(n_4263)
);

CKINVDCx5p33_ASAP7_75t_R g4264 ( 
.A(n_502),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_749),
.Y(n_4265)
);

CKINVDCx5p33_ASAP7_75t_R g4266 ( 
.A(n_689),
.Y(n_4266)
);

CKINVDCx5p33_ASAP7_75t_R g4267 ( 
.A(n_1705),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_890),
.Y(n_4268)
);

CKINVDCx5p33_ASAP7_75t_R g4269 ( 
.A(n_2752),
.Y(n_4269)
);

CKINVDCx5p33_ASAP7_75t_R g4270 ( 
.A(n_496),
.Y(n_4270)
);

CKINVDCx5p33_ASAP7_75t_R g4271 ( 
.A(n_484),
.Y(n_4271)
);

CKINVDCx5p33_ASAP7_75t_R g4272 ( 
.A(n_2707),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_982),
.Y(n_4273)
);

CKINVDCx5p33_ASAP7_75t_R g4274 ( 
.A(n_2838),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_274),
.Y(n_4275)
);

CKINVDCx5p33_ASAP7_75t_R g4276 ( 
.A(n_1347),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_115),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_2824),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_1976),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_2874),
.Y(n_4280)
);

CKINVDCx5p33_ASAP7_75t_R g4281 ( 
.A(n_466),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_423),
.Y(n_4282)
);

HB1xp67_ASAP7_75t_L g4283 ( 
.A(n_2837),
.Y(n_4283)
);

BUFx10_ASAP7_75t_L g4284 ( 
.A(n_1082),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_2137),
.Y(n_4285)
);

CKINVDCx5p33_ASAP7_75t_R g4286 ( 
.A(n_1650),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_55),
.Y(n_4287)
);

CKINVDCx5p33_ASAP7_75t_R g4288 ( 
.A(n_1623),
.Y(n_4288)
);

CKINVDCx5p33_ASAP7_75t_R g4289 ( 
.A(n_2486),
.Y(n_4289)
);

BUFx5_ASAP7_75t_L g4290 ( 
.A(n_2143),
.Y(n_4290)
);

CKINVDCx5p33_ASAP7_75t_R g4291 ( 
.A(n_780),
.Y(n_4291)
);

CKINVDCx5p33_ASAP7_75t_R g4292 ( 
.A(n_2556),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_1862),
.Y(n_4293)
);

INVx1_ASAP7_75t_SL g4294 ( 
.A(n_2055),
.Y(n_4294)
);

CKINVDCx20_ASAP7_75t_R g4295 ( 
.A(n_1986),
.Y(n_4295)
);

BUFx10_ASAP7_75t_L g4296 ( 
.A(n_2653),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_2686),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_715),
.Y(n_4298)
);

BUFx10_ASAP7_75t_L g4299 ( 
.A(n_2684),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_1969),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_1834),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_2286),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_2169),
.Y(n_4303)
);

CKINVDCx5p33_ASAP7_75t_R g4304 ( 
.A(n_2626),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_578),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_1834),
.Y(n_4306)
);

CKINVDCx5p33_ASAP7_75t_R g4307 ( 
.A(n_651),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_2720),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_2566),
.Y(n_4309)
);

CKINVDCx5p33_ASAP7_75t_R g4310 ( 
.A(n_4228),
.Y(n_4310)
);

INVxp67_ASAP7_75t_L g4311 ( 
.A(n_3453),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3110),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3110),
.Y(n_4313)
);

CKINVDCx14_ASAP7_75t_R g4314 ( 
.A(n_3300),
.Y(n_4314)
);

BUFx3_ASAP7_75t_L g4315 ( 
.A(n_3266),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3110),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3110),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3110),
.Y(n_4318)
);

INVxp67_ASAP7_75t_SL g4319 ( 
.A(n_3060),
.Y(n_4319)
);

CKINVDCx5p33_ASAP7_75t_R g4320 ( 
.A(n_3262),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3523),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_3523),
.Y(n_4322)
);

BUFx3_ASAP7_75t_L g4323 ( 
.A(n_3794),
.Y(n_4323)
);

CKINVDCx20_ASAP7_75t_R g4324 ( 
.A(n_3357),
.Y(n_4324)
);

CKINVDCx5p33_ASAP7_75t_R g4325 ( 
.A(n_3265),
.Y(n_4325)
);

INVxp33_ASAP7_75t_L g4326 ( 
.A(n_3020),
.Y(n_4326)
);

CKINVDCx5p33_ASAP7_75t_R g4327 ( 
.A(n_3379),
.Y(n_4327)
);

CKINVDCx20_ASAP7_75t_R g4328 ( 
.A(n_3426),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3523),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3523),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_3523),
.Y(n_4331)
);

INVx2_ASAP7_75t_SL g4332 ( 
.A(n_3586),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_3922),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4290),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4290),
.Y(n_4335)
);

CKINVDCx5p33_ASAP7_75t_R g4336 ( 
.A(n_3975),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4290),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4290),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4290),
.Y(n_4339)
);

CKINVDCx20_ASAP7_75t_R g4340 ( 
.A(n_4075),
.Y(n_4340)
);

CKINVDCx5p33_ASAP7_75t_R g4341 ( 
.A(n_4000),
.Y(n_4341)
);

BUFx3_ASAP7_75t_L g4342 ( 
.A(n_4238),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_3033),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_4165),
.Y(n_4344)
);

CKINVDCx5p33_ASAP7_75t_R g4345 ( 
.A(n_3188),
.Y(n_4345)
);

CKINVDCx5p33_ASAP7_75t_R g4346 ( 
.A(n_3219),
.Y(n_4346)
);

CKINVDCx16_ASAP7_75t_R g4347 ( 
.A(n_2953),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_3160),
.Y(n_4348)
);

CKINVDCx16_ASAP7_75t_R g4349 ( 
.A(n_2958),
.Y(n_4349)
);

BUFx3_ASAP7_75t_L g4350 ( 
.A(n_2998),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_3192),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3196),
.Y(n_4352)
);

CKINVDCx14_ASAP7_75t_R g4353 ( 
.A(n_4123),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3227),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3247),
.Y(n_4355)
);

INVx3_ASAP7_75t_L g4356 ( 
.A(n_3011),
.Y(n_4356)
);

INVxp33_ASAP7_75t_L g4357 ( 
.A(n_3907),
.Y(n_4357)
);

INVxp33_ASAP7_75t_SL g4358 ( 
.A(n_3057),
.Y(n_4358)
);

CKINVDCx5p33_ASAP7_75t_R g4359 ( 
.A(n_4156),
.Y(n_4359)
);

BUFx6f_ASAP7_75t_L g4360 ( 
.A(n_3018),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3331),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3333),
.Y(n_4362)
);

CKINVDCx5p33_ASAP7_75t_R g4363 ( 
.A(n_2987),
.Y(n_4363)
);

CKINVDCx14_ASAP7_75t_R g4364 ( 
.A(n_3781),
.Y(n_4364)
);

INVxp33_ASAP7_75t_SL g4365 ( 
.A(n_3070),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_3355),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_3377),
.Y(n_4367)
);

BUFx5_ASAP7_75t_L g4368 ( 
.A(n_2922),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3431),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3443),
.Y(n_4370)
);

CKINVDCx16_ASAP7_75t_R g4371 ( 
.A(n_3104),
.Y(n_4371)
);

INVxp33_ASAP7_75t_SL g4372 ( 
.A(n_3162),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3455),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_3521),
.Y(n_4374)
);

INVx1_ASAP7_75t_SL g4375 ( 
.A(n_3107),
.Y(n_4375)
);

HB1xp67_ASAP7_75t_L g4376 ( 
.A(n_3482),
.Y(n_4376)
);

CKINVDCx14_ASAP7_75t_R g4377 ( 
.A(n_3151),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_3528),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3534),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3536),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3539),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_3572),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_3513),
.Y(n_4383)
);

CKINVDCx16_ASAP7_75t_R g4384 ( 
.A(n_3716),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_3600),
.Y(n_4385)
);

BUFx3_ASAP7_75t_L g4386 ( 
.A(n_3049),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_3611),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3676),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_3685),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_3060),
.B(n_4109),
.Y(n_4390)
);

INVxp67_ASAP7_75t_L g4391 ( 
.A(n_3309),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_3709),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3713),
.Y(n_4393)
);

CKINVDCx16_ASAP7_75t_R g4394 ( 
.A(n_3812),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_3770),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_3809),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_3829),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3882),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_3919),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_3920),
.Y(n_4400)
);

INVxp67_ASAP7_75t_L g4401 ( 
.A(n_3342),
.Y(n_4401)
);

CKINVDCx5p33_ASAP7_75t_R g4402 ( 
.A(n_3831),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3957),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3974),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_3983),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_3855),
.Y(n_4406)
);

CKINVDCx20_ASAP7_75t_R g4407 ( 
.A(n_3877),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4009),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_3921),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4010),
.Y(n_4410)
);

CKINVDCx14_ASAP7_75t_R g4411 ( 
.A(n_3567),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_2947),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4074),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4089),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_2974),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4103),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4185),
.Y(n_4417)
);

CKINVDCx16_ASAP7_75t_R g4418 ( 
.A(n_3586),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4250),
.Y(n_4419)
);

INVx1_ASAP7_75t_SL g4420 ( 
.A(n_3965),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4255),
.Y(n_4421)
);

CKINVDCx5p33_ASAP7_75t_R g4422 ( 
.A(n_2978),
.Y(n_4422)
);

INVx2_ASAP7_75t_SL g4423 ( 
.A(n_3649),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4275),
.Y(n_4424)
);

CKINVDCx5p33_ASAP7_75t_R g4425 ( 
.A(n_3007),
.Y(n_4425)
);

INVxp67_ASAP7_75t_L g4426 ( 
.A(n_3993),
.Y(n_4426)
);

CKINVDCx5p33_ASAP7_75t_R g4427 ( 
.A(n_3032),
.Y(n_4427)
);

CKINVDCx20_ASAP7_75t_R g4428 ( 
.A(n_2928),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4277),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4287),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_3018),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3018),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3083),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_3083),
.Y(n_4434)
);

CKINVDCx20_ASAP7_75t_R g4435 ( 
.A(n_2934),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_3083),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3420),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_3420),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_2939),
.Y(n_4439)
);

BUFx2_ASAP7_75t_SL g4440 ( 
.A(n_3649),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3420),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_3042),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_3044),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3845),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3845),
.Y(n_4445)
);

INVxp67_ASAP7_75t_SL g4446 ( 
.A(n_4109),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3845),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4057),
.B(n_0),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_3014),
.Y(n_4449)
);

CKINVDCx5p33_ASAP7_75t_R g4450 ( 
.A(n_3084),
.Y(n_4450)
);

CKINVDCx5p33_ASAP7_75t_R g4451 ( 
.A(n_3121),
.Y(n_4451)
);

HB1xp67_ASAP7_75t_L g4452 ( 
.A(n_3239),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_3123),
.Y(n_4453)
);

INVxp67_ASAP7_75t_L g4454 ( 
.A(n_4079),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_3136),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_3157),
.Y(n_4456)
);

CKINVDCx20_ASAP7_75t_R g4457 ( 
.A(n_2943),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_3885),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_3885),
.Y(n_4459)
);

INVxp67_ASAP7_75t_L g4460 ( 
.A(n_4111),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_3885),
.Y(n_4461)
);

BUFx2_ASAP7_75t_L g4462 ( 
.A(n_3167),
.Y(n_4462)
);

BUFx3_ASAP7_75t_L g4463 ( 
.A(n_3050),
.Y(n_4463)
);

INVx1_ASAP7_75t_SL g4464 ( 
.A(n_4046),
.Y(n_4464)
);

CKINVDCx5p33_ASAP7_75t_R g4465 ( 
.A(n_3179),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_3999),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_3999),
.Y(n_4467)
);

BUFx3_ASAP7_75t_L g4468 ( 
.A(n_3126),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_3999),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_3206),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4082),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4082),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4082),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4095),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4095),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4095),
.Y(n_4476)
);

CKINVDCx5p33_ASAP7_75t_R g4477 ( 
.A(n_3207),
.Y(n_4477)
);

CKINVDCx5p33_ASAP7_75t_R g4478 ( 
.A(n_3208),
.Y(n_4478)
);

CKINVDCx16_ASAP7_75t_R g4479 ( 
.A(n_3751),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_3228),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_3783),
.Y(n_4481)
);

INVxp67_ASAP7_75t_SL g4482 ( 
.A(n_3350),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3990),
.Y(n_4483)
);

CKINVDCx5p33_ASAP7_75t_R g4484 ( 
.A(n_3253),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4230),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_2954),
.Y(n_4486)
);

HB1xp67_ASAP7_75t_L g4487 ( 
.A(n_3380),
.Y(n_4487)
);

HB1xp67_ASAP7_75t_L g4488 ( 
.A(n_3798),
.Y(n_4488)
);

CKINVDCx5p33_ASAP7_75t_R g4489 ( 
.A(n_3254),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_2954),
.Y(n_4490)
);

INVxp33_ASAP7_75t_SL g4491 ( 
.A(n_3997),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_3310),
.Y(n_4492)
);

INVxp67_ASAP7_75t_SL g4493 ( 
.A(n_3821),
.Y(n_4493)
);

INVxp67_ASAP7_75t_SL g4494 ( 
.A(n_4038),
.Y(n_4494)
);

CKINVDCx20_ASAP7_75t_R g4495 ( 
.A(n_2950),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_2954),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_3318),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_3074),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3074),
.Y(n_4499)
);

INVx2_ASAP7_75t_SL g4500 ( 
.A(n_3751),
.Y(n_4500)
);

BUFx3_ASAP7_75t_L g4501 ( 
.A(n_3177),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_3074),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_3319),
.Y(n_4503)
);

CKINVDCx5p33_ASAP7_75t_R g4504 ( 
.A(n_3330),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_3140),
.Y(n_4505)
);

NOR2xp67_ASAP7_75t_L g4506 ( 
.A(n_3230),
.B(n_0),
.Y(n_4506)
);

CKINVDCx5p33_ASAP7_75t_R g4507 ( 
.A(n_3332),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_3140),
.Y(n_4508)
);

CKINVDCx5p33_ASAP7_75t_R g4509 ( 
.A(n_3336),
.Y(n_4509)
);

CKINVDCx5p33_ASAP7_75t_R g4510 ( 
.A(n_3346),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_3140),
.Y(n_4511)
);

CKINVDCx14_ASAP7_75t_R g4512 ( 
.A(n_4159),
.Y(n_4512)
);

BUFx6f_ASAP7_75t_L g4513 ( 
.A(n_3166),
.Y(n_4513)
);

CKINVDCx16_ASAP7_75t_R g4514 ( 
.A(n_4159),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_3166),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_3166),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_3244),
.Y(n_4517)
);

INVxp67_ASAP7_75t_L g4518 ( 
.A(n_4119),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_3244),
.Y(n_4519)
);

CKINVDCx20_ASAP7_75t_R g4520 ( 
.A(n_2972),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3244),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_3468),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_3468),
.Y(n_4523)
);

INVx3_ASAP7_75t_L g4524 ( 
.A(n_3213),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3468),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3540),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_3540),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_3540),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_3365),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3551),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_3399),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_3551),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_3551),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_3618),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3618),
.Y(n_4535)
);

CKINVDCx20_ASAP7_75t_R g4536 ( 
.A(n_3005),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3618),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_3680),
.Y(n_4538)
);

INVx2_ASAP7_75t_SL g4539 ( 
.A(n_2938),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_3680),
.Y(n_4540)
);

CKINVDCx5p33_ASAP7_75t_R g4541 ( 
.A(n_3409),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_3680),
.Y(n_4542)
);

BUFx3_ASAP7_75t_L g4543 ( 
.A(n_3218),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3689),
.Y(n_4544)
);

CKINVDCx16_ASAP7_75t_R g4545 ( 
.A(n_2938),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_3689),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_3412),
.Y(n_4547)
);

INVxp67_ASAP7_75t_L g4548 ( 
.A(n_4283),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_3689),
.Y(n_4549)
);

INVx1_ASAP7_75t_SL g4550 ( 
.A(n_3209),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_3840),
.Y(n_4551)
);

BUFx3_ASAP7_75t_L g4552 ( 
.A(n_3225),
.Y(n_4552)
);

CKINVDCx20_ASAP7_75t_R g4553 ( 
.A(n_3021),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_3840),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_3840),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_3860),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_3860),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_3860),
.Y(n_4558)
);

CKINVDCx5p33_ASAP7_75t_R g4559 ( 
.A(n_3435),
.Y(n_4559)
);

INVxp33_ASAP7_75t_L g4560 ( 
.A(n_2923),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3912),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_3912),
.Y(n_4562)
);

CKINVDCx5p33_ASAP7_75t_R g4563 ( 
.A(n_3445),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_3912),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_3939),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3939),
.Y(n_4566)
);

CKINVDCx5p33_ASAP7_75t_R g4567 ( 
.A(n_3446),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_3939),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_3941),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_3941),
.Y(n_4570)
);

INVxp67_ASAP7_75t_SL g4571 ( 
.A(n_3941),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4026),
.Y(n_4572)
);

CKINVDCx20_ASAP7_75t_R g4573 ( 
.A(n_3027),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4026),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4026),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4042),
.Y(n_4576)
);

INVxp67_ASAP7_75t_L g4577 ( 
.A(n_3015),
.Y(n_4577)
);

BUFx6f_ASAP7_75t_L g4578 ( 
.A(n_4042),
.Y(n_4578)
);

CKINVDCx5p33_ASAP7_75t_R g4579 ( 
.A(n_3472),
.Y(n_4579)
);

CKINVDCx16_ASAP7_75t_R g4580 ( 
.A(n_3015),
.Y(n_4580)
);

CKINVDCx5p33_ASAP7_75t_R g4581 ( 
.A(n_3487),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4042),
.Y(n_4582)
);

CKINVDCx20_ASAP7_75t_R g4583 ( 
.A(n_3075),
.Y(n_4583)
);

BUFx6f_ASAP7_75t_L g4584 ( 
.A(n_4084),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4084),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4084),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4187),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4187),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4187),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4232),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4232),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4232),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4273),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4273),
.Y(n_4594)
);

CKINVDCx14_ASAP7_75t_R g4595 ( 
.A(n_3072),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4273),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_3231),
.Y(n_4597)
);

CKINVDCx5p33_ASAP7_75t_R g4598 ( 
.A(n_3488),
.Y(n_4598)
);

INVx2_ASAP7_75t_SL g4599 ( 
.A(n_3072),
.Y(n_4599)
);

INVx1_ASAP7_75t_SL g4600 ( 
.A(n_3668),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_3237),
.Y(n_4601)
);

CKINVDCx16_ASAP7_75t_R g4602 ( 
.A(n_3086),
.Y(n_4602)
);

BUFx3_ASAP7_75t_L g4603 ( 
.A(n_3250),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_3282),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_3316),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_3504),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_3415),
.Y(n_4607)
);

CKINVDCx16_ASAP7_75t_R g4608 ( 
.A(n_3086),
.Y(n_4608)
);

INVx2_ASAP7_75t_L g4609 ( 
.A(n_3444),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_3459),
.Y(n_4610)
);

CKINVDCx5p33_ASAP7_75t_R g4611 ( 
.A(n_3522),
.Y(n_4611)
);

CKINVDCx5p33_ASAP7_75t_R g4612 ( 
.A(n_3560),
.Y(n_4612)
);

CKINVDCx5p33_ASAP7_75t_R g4613 ( 
.A(n_3563),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_3467),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_3470),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_3479),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_3480),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_3485),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_3543),
.Y(n_4619)
);

BUFx6f_ASAP7_75t_L g4620 ( 
.A(n_3554),
.Y(n_4620)
);

CKINVDCx16_ASAP7_75t_R g4621 ( 
.A(n_3178),
.Y(n_4621)
);

BUFx6f_ASAP7_75t_L g4622 ( 
.A(n_3630),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_3671),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_3927),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_3996),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_3584),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4054),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_3588),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4066),
.Y(n_4629)
);

INVxp67_ASAP7_75t_SL g4630 ( 
.A(n_4201),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4300),
.Y(n_4631)
);

BUFx6f_ASAP7_75t_L g4632 ( 
.A(n_2970),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4301),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4305),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_2926),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4306),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4308),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4309),
.Y(n_4638)
);

BUFx2_ASAP7_75t_L g4639 ( 
.A(n_3589),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_2929),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_2930),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_2931),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_2935),
.Y(n_4643)
);

CKINVDCx20_ASAP7_75t_R g4644 ( 
.A(n_3109),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_3593),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_2937),
.Y(n_4646)
);

INVxp33_ASAP7_75t_L g4647 ( 
.A(n_2948),
.Y(n_4647)
);

OR2x2_ASAP7_75t_L g4648 ( 
.A(n_3802),
.B(n_0),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_2949),
.Y(n_4649)
);

INVxp67_ASAP7_75t_L g4650 ( 
.A(n_3178),
.Y(n_4650)
);

BUFx3_ASAP7_75t_L g4651 ( 
.A(n_3220),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_2956),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_2959),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_3622),
.Y(n_4654)
);

BUFx3_ASAP7_75t_L g4655 ( 
.A(n_3220),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_2968),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_2975),
.Y(n_4657)
);

CKINVDCx5p33_ASAP7_75t_R g4658 ( 
.A(n_3627),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_3632),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_2976),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_3293),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_2977),
.Y(n_4662)
);

BUFx5_ASAP7_75t_L g4663 ( 
.A(n_2980),
.Y(n_4663)
);

BUFx3_ASAP7_75t_L g4664 ( 
.A(n_3293),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_2982),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_3643),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_2985),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_3645),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_2986),
.Y(n_4669)
);

CKINVDCx5p33_ASAP7_75t_R g4670 ( 
.A(n_3681),
.Y(n_4670)
);

CKINVDCx5p33_ASAP7_75t_R g4671 ( 
.A(n_3710),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_2988),
.Y(n_4672)
);

CKINVDCx5p33_ASAP7_75t_R g4673 ( 
.A(n_3732),
.Y(n_4673)
);

BUFx6f_ASAP7_75t_L g4674 ( 
.A(n_3038),
.Y(n_4674)
);

BUFx3_ASAP7_75t_L g4675 ( 
.A(n_3308),
.Y(n_4675)
);

CKINVDCx16_ASAP7_75t_R g4676 ( 
.A(n_3308),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_2990),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_3777),
.Y(n_4678)
);

BUFx2_ASAP7_75t_L g4679 ( 
.A(n_3782),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_2991),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_3000),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_3001),
.Y(n_4682)
);

CKINVDCx20_ASAP7_75t_R g4683 ( 
.A(n_3116),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_3003),
.Y(n_4684)
);

CKINVDCx5p33_ASAP7_75t_R g4685 ( 
.A(n_3801),
.Y(n_4685)
);

CKINVDCx20_ASAP7_75t_R g4686 ( 
.A(n_3119),
.Y(n_4686)
);

CKINVDCx5p33_ASAP7_75t_R g4687 ( 
.A(n_3818),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_3006),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_3008),
.Y(n_4689)
);

CKINVDCx5p33_ASAP7_75t_R g4690 ( 
.A(n_3822),
.Y(n_4690)
);

INVxp67_ASAP7_75t_SL g4691 ( 
.A(n_4092),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_3029),
.Y(n_4692)
);

BUFx3_ASAP7_75t_L g4693 ( 
.A(n_3428),
.Y(n_4693)
);

INVxp67_ASAP7_75t_L g4694 ( 
.A(n_3428),
.Y(n_4694)
);

BUFx6f_ASAP7_75t_L g4695 ( 
.A(n_3082),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_3856),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_3035),
.Y(n_4697)
);

CKINVDCx5p33_ASAP7_75t_R g4698 ( 
.A(n_3862),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_3039),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_3045),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_3046),
.Y(n_4701)
);

NOR2xp67_ASAP7_75t_L g4702 ( 
.A(n_3305),
.B(n_1),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_3054),
.Y(n_4703)
);

CKINVDCx20_ASAP7_75t_R g4704 ( 
.A(n_3129),
.Y(n_4704)
);

INVxp33_ASAP7_75t_L g4705 ( 
.A(n_3055),
.Y(n_4705)
);

CKINVDCx16_ASAP7_75t_R g4706 ( 
.A(n_4299),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_3058),
.Y(n_4707)
);

INVxp67_ASAP7_75t_L g4708 ( 
.A(n_3489),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_3063),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_3090),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_3093),
.Y(n_4711)
);

CKINVDCx20_ASAP7_75t_R g4712 ( 
.A(n_3145),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_3094),
.Y(n_4713)
);

BUFx3_ASAP7_75t_L g4714 ( 
.A(n_3489),
.Y(n_4714)
);

CKINVDCx5p33_ASAP7_75t_R g4715 ( 
.A(n_3872),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_3097),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_3573),
.B(n_1),
.Y(n_4717)
);

INVxp33_ASAP7_75t_L g4718 ( 
.A(n_3098),
.Y(n_4718)
);

CKINVDCx20_ASAP7_75t_R g4719 ( 
.A(n_3171),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_3106),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_3124),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_3125),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_3133),
.Y(n_4723)
);

INVxp67_ASAP7_75t_SL g4724 ( 
.A(n_4236),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_3137),
.Y(n_4725)
);

BUFx2_ASAP7_75t_L g4726 ( 
.A(n_3899),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_3901),
.Y(n_4727)
);

BUFx3_ASAP7_75t_L g4728 ( 
.A(n_3509),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_3142),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_3143),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_3147),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_3148),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_3906),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_3150),
.Y(n_4734)
);

CKINVDCx5p33_ASAP7_75t_R g4735 ( 
.A(n_4320),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4319),
.B(n_3023),
.Y(n_4736)
);

CKINVDCx20_ASAP7_75t_R g4737 ( 
.A(n_4428),
.Y(n_4737)
);

CKINVDCx5p33_ASAP7_75t_R g4738 ( 
.A(n_4325),
.Y(n_4738)
);

CKINVDCx5p33_ASAP7_75t_R g4739 ( 
.A(n_4327),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4571),
.Y(n_4740)
);

INVxp67_ASAP7_75t_SL g4741 ( 
.A(n_4390),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4360),
.Y(n_4742)
);

CKINVDCx20_ASAP7_75t_R g4743 ( 
.A(n_4435),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_4333),
.Y(n_4744)
);

BUFx6f_ASAP7_75t_L g4745 ( 
.A(n_4360),
.Y(n_4745)
);

INVxp67_ASAP7_75t_SL g4746 ( 
.A(n_4356),
.Y(n_4746)
);

CKINVDCx5p33_ASAP7_75t_R g4747 ( 
.A(n_4336),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4513),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4446),
.B(n_3127),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4486),
.Y(n_4750)
);

CKINVDCx5p33_ASAP7_75t_R g4751 ( 
.A(n_4341),
.Y(n_4751)
);

INVx3_ASAP7_75t_L g4752 ( 
.A(n_4513),
.Y(n_4752)
);

INVxp33_ASAP7_75t_L g4753 ( 
.A(n_4376),
.Y(n_4753)
);

CKINVDCx20_ASAP7_75t_R g4754 ( 
.A(n_4457),
.Y(n_4754)
);

CKINVDCx16_ASAP7_75t_R g4755 ( 
.A(n_4324),
.Y(n_4755)
);

CKINVDCx20_ASAP7_75t_R g4756 ( 
.A(n_4495),
.Y(n_4756)
);

HB1xp67_ASAP7_75t_L g4757 ( 
.A(n_4363),
.Y(n_4757)
);

CKINVDCx5p33_ASAP7_75t_R g4758 ( 
.A(n_4344),
.Y(n_4758)
);

HB1xp67_ASAP7_75t_L g4759 ( 
.A(n_4383),
.Y(n_4759)
);

NOR2xp33_ASAP7_75t_L g4760 ( 
.A(n_4359),
.B(n_3932),
.Y(n_4760)
);

INVxp67_ASAP7_75t_SL g4761 ( 
.A(n_4524),
.Y(n_4761)
);

CKINVDCx20_ASAP7_75t_R g4762 ( 
.A(n_4520),
.Y(n_4762)
);

CKINVDCx5p33_ASAP7_75t_R g4763 ( 
.A(n_4412),
.Y(n_4763)
);

CKINVDCx5p33_ASAP7_75t_R g4764 ( 
.A(n_4415),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4578),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4578),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4584),
.Y(n_4767)
);

BUFx3_ASAP7_75t_L g4768 ( 
.A(n_4315),
.Y(n_4768)
);

HB1xp67_ASAP7_75t_L g4769 ( 
.A(n_4402),
.Y(n_4769)
);

INVxp67_ASAP7_75t_SL g4770 ( 
.A(n_4350),
.Y(n_4770)
);

CKINVDCx5p33_ASAP7_75t_R g4771 ( 
.A(n_4422),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4584),
.Y(n_4772)
);

CKINVDCx5p33_ASAP7_75t_R g4773 ( 
.A(n_4425),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_4427),
.Y(n_4774)
);

CKINVDCx16_ASAP7_75t_R g4775 ( 
.A(n_4328),
.Y(n_4775)
);

CKINVDCx20_ASAP7_75t_R g4776 ( 
.A(n_4536),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4431),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4432),
.Y(n_4778)
);

CKINVDCx5p33_ASAP7_75t_R g4779 ( 
.A(n_4442),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4433),
.Y(n_4780)
);

CKINVDCx20_ASAP7_75t_R g4781 ( 
.A(n_4553),
.Y(n_4781)
);

CKINVDCx5p33_ASAP7_75t_R g4782 ( 
.A(n_4443),
.Y(n_4782)
);

HB1xp67_ASAP7_75t_L g4783 ( 
.A(n_4406),
.Y(n_4783)
);

BUFx6f_ASAP7_75t_L g4784 ( 
.A(n_4620),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4434),
.Y(n_4785)
);

INVxp33_ASAP7_75t_SL g4786 ( 
.A(n_4310),
.Y(n_4786)
);

CKINVDCx5p33_ASAP7_75t_R g4787 ( 
.A(n_4450),
.Y(n_4787)
);

CKINVDCx5p33_ASAP7_75t_R g4788 ( 
.A(n_4451),
.Y(n_4788)
);

CKINVDCx5p33_ASAP7_75t_R g4789 ( 
.A(n_4453),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4436),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4437),
.Y(n_4791)
);

CKINVDCx5p33_ASAP7_75t_R g4792 ( 
.A(n_4455),
.Y(n_4792)
);

CKINVDCx20_ASAP7_75t_R g4793 ( 
.A(n_4573),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4438),
.Y(n_4794)
);

CKINVDCx20_ASAP7_75t_R g4795 ( 
.A(n_4583),
.Y(n_4795)
);

CKINVDCx20_ASAP7_75t_R g4796 ( 
.A(n_4644),
.Y(n_4796)
);

CKINVDCx5p33_ASAP7_75t_R g4797 ( 
.A(n_4456),
.Y(n_4797)
);

CKINVDCx5p33_ASAP7_75t_R g4798 ( 
.A(n_4465),
.Y(n_4798)
);

HB1xp67_ASAP7_75t_L g4799 ( 
.A(n_4409),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4441),
.Y(n_4800)
);

INVxp67_ASAP7_75t_SL g4801 ( 
.A(n_4386),
.Y(n_4801)
);

INVxp33_ASAP7_75t_L g4802 ( 
.A(n_4452),
.Y(n_4802)
);

INVxp33_ASAP7_75t_SL g4803 ( 
.A(n_4345),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4444),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4445),
.Y(n_4805)
);

CKINVDCx20_ASAP7_75t_R g4806 ( 
.A(n_4683),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4447),
.Y(n_4807)
);

CKINVDCx5p33_ASAP7_75t_R g4808 ( 
.A(n_4470),
.Y(n_4808)
);

INVxp67_ASAP7_75t_L g4809 ( 
.A(n_4440),
.Y(n_4809)
);

CKINVDCx20_ASAP7_75t_R g4810 ( 
.A(n_4686),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4458),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4459),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4461),
.Y(n_4813)
);

NOR2xp33_ASAP7_75t_L g4814 ( 
.A(n_4358),
.B(n_3935),
.Y(n_4814)
);

CKINVDCx20_ASAP7_75t_R g4815 ( 
.A(n_4704),
.Y(n_4815)
);

INVxp67_ASAP7_75t_SL g4816 ( 
.A(n_4463),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4466),
.Y(n_4817)
);

CKINVDCx20_ASAP7_75t_R g4818 ( 
.A(n_4712),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4365),
.B(n_3946),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4467),
.Y(n_4820)
);

INVxp67_ASAP7_75t_SL g4821 ( 
.A(n_4468),
.Y(n_4821)
);

INVx2_ASAP7_75t_L g4822 ( 
.A(n_4511),
.Y(n_4822)
);

INVxp67_ASAP7_75t_SL g4823 ( 
.A(n_4501),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4523),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4469),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4471),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_4477),
.Y(n_4827)
);

CKINVDCx5p33_ASAP7_75t_R g4828 ( 
.A(n_4478),
.Y(n_4828)
);

CKINVDCx14_ASAP7_75t_R g4829 ( 
.A(n_4314),
.Y(n_4829)
);

INVxp67_ASAP7_75t_L g4830 ( 
.A(n_4462),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4472),
.Y(n_4831)
);

CKINVDCx20_ASAP7_75t_R g4832 ( 
.A(n_4719),
.Y(n_4832)
);

CKINVDCx20_ASAP7_75t_R g4833 ( 
.A(n_4340),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4473),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4474),
.Y(n_4835)
);

CKINVDCx5p33_ASAP7_75t_R g4836 ( 
.A(n_4480),
.Y(n_4836)
);

INVxp67_ASAP7_75t_SL g4837 ( 
.A(n_4543),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4475),
.Y(n_4838)
);

CKINVDCx20_ASAP7_75t_R g4839 ( 
.A(n_4407),
.Y(n_4839)
);

CKINVDCx5p33_ASAP7_75t_R g4840 ( 
.A(n_4484),
.Y(n_4840)
);

CKINVDCx20_ASAP7_75t_R g4841 ( 
.A(n_4347),
.Y(n_4841)
);

INVxp67_ASAP7_75t_SL g4842 ( 
.A(n_4552),
.Y(n_4842)
);

INVx2_ASAP7_75t_L g4843 ( 
.A(n_4556),
.Y(n_4843)
);

INVxp67_ASAP7_75t_SL g4844 ( 
.A(n_4603),
.Y(n_4844)
);

OR2x2_ASAP7_75t_L g4845 ( 
.A(n_4375),
.B(n_3841),
.Y(n_4845)
);

CKINVDCx5p33_ASAP7_75t_R g4846 ( 
.A(n_4489),
.Y(n_4846)
);

CKINVDCx16_ASAP7_75t_R g4847 ( 
.A(n_4349),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4476),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4353),
.B(n_4053),
.Y(n_4849)
);

CKINVDCx20_ASAP7_75t_R g4850 ( 
.A(n_4371),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4490),
.Y(n_4851)
);

BUFx2_ASAP7_75t_L g4852 ( 
.A(n_4346),
.Y(n_4852)
);

INVx1_ASAP7_75t_SL g4853 ( 
.A(n_4464),
.Y(n_4853)
);

CKINVDCx20_ASAP7_75t_R g4854 ( 
.A(n_4384),
.Y(n_4854)
);

INVxp67_ASAP7_75t_SL g4855 ( 
.A(n_4620),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4496),
.Y(n_4856)
);

INVxp67_ASAP7_75t_SL g4857 ( 
.A(n_4622),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4498),
.Y(n_4858)
);

CKINVDCx20_ASAP7_75t_R g4859 ( 
.A(n_4394),
.Y(n_4859)
);

CKINVDCx5p33_ASAP7_75t_R g4860 ( 
.A(n_4492),
.Y(n_4860)
);

CKINVDCx20_ASAP7_75t_R g4861 ( 
.A(n_4512),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4499),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4502),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_4497),
.Y(n_4864)
);

CKINVDCx20_ASAP7_75t_R g4865 ( 
.A(n_4595),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4505),
.Y(n_4866)
);

NOR2xp33_ASAP7_75t_L g4867 ( 
.A(n_4372),
.B(n_3972),
.Y(n_4867)
);

BUFx6f_ASAP7_75t_L g4868 ( 
.A(n_4622),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4508),
.Y(n_4869)
);

CKINVDCx5p33_ASAP7_75t_R g4870 ( 
.A(n_4503),
.Y(n_4870)
);

CKINVDCx20_ASAP7_75t_R g4871 ( 
.A(n_4364),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4515),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4516),
.Y(n_4873)
);

CKINVDCx20_ASAP7_75t_R g4874 ( 
.A(n_4377),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4517),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4519),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4521),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4630),
.B(n_3729),
.Y(n_4878)
);

INVxp67_ASAP7_75t_L g4879 ( 
.A(n_4628),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4522),
.Y(n_4880)
);

CKINVDCx5p33_ASAP7_75t_R g4881 ( 
.A(n_4504),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4525),
.Y(n_4882)
);

CKINVDCx20_ASAP7_75t_R g4883 ( 
.A(n_4411),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4526),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4527),
.Y(n_4885)
);

CKINVDCx20_ASAP7_75t_R g4886 ( 
.A(n_4550),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4691),
.B(n_3246),
.Y(n_4887)
);

CKINVDCx20_ASAP7_75t_R g4888 ( 
.A(n_4600),
.Y(n_4888)
);

INVxp67_ASAP7_75t_SL g4889 ( 
.A(n_4661),
.Y(n_4889)
);

CKINVDCx16_ASAP7_75t_R g4890 ( 
.A(n_4418),
.Y(n_4890)
);

HB1xp67_ASAP7_75t_L g4891 ( 
.A(n_4507),
.Y(n_4891)
);

CKINVDCx5p33_ASAP7_75t_R g4892 ( 
.A(n_4509),
.Y(n_4892)
);

CKINVDCx20_ASAP7_75t_R g4893 ( 
.A(n_4510),
.Y(n_4893)
);

CKINVDCx20_ASAP7_75t_R g4894 ( 
.A(n_4529),
.Y(n_4894)
);

CKINVDCx20_ASAP7_75t_R g4895 ( 
.A(n_4531),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_4491),
.B(n_4541),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_4547),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4528),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4530),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4532),
.Y(n_4900)
);

CKINVDCx20_ASAP7_75t_R g4901 ( 
.A(n_4559),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4533),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4534),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4535),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4537),
.Y(n_4905)
);

CKINVDCx5p33_ASAP7_75t_R g4906 ( 
.A(n_4563),
.Y(n_4906)
);

CKINVDCx5p33_ASAP7_75t_R g4907 ( 
.A(n_4567),
.Y(n_4907)
);

CKINVDCx20_ASAP7_75t_R g4908 ( 
.A(n_4579),
.Y(n_4908)
);

INVxp67_ASAP7_75t_L g4909 ( 
.A(n_4639),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4538),
.Y(n_4910)
);

CKINVDCx5p33_ASAP7_75t_R g4911 ( 
.A(n_4581),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4540),
.Y(n_4912)
);

HB1xp67_ASAP7_75t_L g4913 ( 
.A(n_4598),
.Y(n_4913)
);

CKINVDCx5p33_ASAP7_75t_R g4914 ( 
.A(n_4606),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4542),
.Y(n_4915)
);

CKINVDCx20_ASAP7_75t_R g4916 ( 
.A(n_4611),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4544),
.Y(n_4917)
);

AND2x4_ASAP7_75t_L g4918 ( 
.A(n_4482),
.B(n_3091),
.Y(n_4918)
);

CKINVDCx20_ASAP7_75t_R g4919 ( 
.A(n_4612),
.Y(n_4919)
);

HB1xp67_ASAP7_75t_L g4920 ( 
.A(n_4613),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4546),
.Y(n_4921)
);

CKINVDCx5p33_ASAP7_75t_R g4922 ( 
.A(n_4626),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_4645),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4549),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4551),
.Y(n_4925)
);

CKINVDCx5p33_ASAP7_75t_R g4926 ( 
.A(n_4654),
.Y(n_4926)
);

CKINVDCx20_ASAP7_75t_R g4927 ( 
.A(n_4658),
.Y(n_4927)
);

CKINVDCx20_ASAP7_75t_R g4928 ( 
.A(n_4659),
.Y(n_4928)
);

INVxp67_ASAP7_75t_L g4929 ( 
.A(n_4679),
.Y(n_4929)
);

CKINVDCx16_ASAP7_75t_R g4930 ( 
.A(n_4479),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4554),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4555),
.Y(n_4932)
);

CKINVDCx20_ASAP7_75t_R g4933 ( 
.A(n_4666),
.Y(n_4933)
);

CKINVDCx20_ASAP7_75t_R g4934 ( 
.A(n_4668),
.Y(n_4934)
);

CKINVDCx20_ASAP7_75t_R g4935 ( 
.A(n_4670),
.Y(n_4935)
);

HB1xp67_ASAP7_75t_L g4936 ( 
.A(n_4671),
.Y(n_4936)
);

CKINVDCx20_ASAP7_75t_R g4937 ( 
.A(n_4673),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4557),
.Y(n_4938)
);

CKINVDCx5p33_ASAP7_75t_R g4939 ( 
.A(n_4678),
.Y(n_4939)
);

INVxp67_ASAP7_75t_L g4940 ( 
.A(n_4726),
.Y(n_4940)
);

INVxp33_ASAP7_75t_SL g4941 ( 
.A(n_4685),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4558),
.Y(n_4942)
);

INVxp67_ASAP7_75t_L g4943 ( 
.A(n_4651),
.Y(n_4943)
);

CKINVDCx20_ASAP7_75t_R g4944 ( 
.A(n_4687),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4690),
.B(n_4696),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_4698),
.Y(n_4946)
);

CKINVDCx14_ASAP7_75t_R g4947 ( 
.A(n_4715),
.Y(n_4947)
);

CKINVDCx5p33_ASAP7_75t_R g4948 ( 
.A(n_4727),
.Y(n_4948)
);

CKINVDCx20_ASAP7_75t_R g4949 ( 
.A(n_4733),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4561),
.Y(n_4950)
);

NOR2xp67_ASAP7_75t_L g4951 ( 
.A(n_4577),
.B(n_3389),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4562),
.Y(n_4952)
);

CKINVDCx5p33_ASAP7_75t_R g4953 ( 
.A(n_4545),
.Y(n_4953)
);

NOR2xp67_ASAP7_75t_L g4954 ( 
.A(n_4650),
.B(n_4233),
.Y(n_4954)
);

INVx2_ASAP7_75t_L g4955 ( 
.A(n_4564),
.Y(n_4955)
);

INVxp67_ASAP7_75t_SL g4956 ( 
.A(n_4323),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4565),
.Y(n_4957)
);

NOR2xp33_ASAP7_75t_L g4958 ( 
.A(n_4518),
.B(n_3979),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_4580),
.Y(n_4959)
);

CKINVDCx20_ASAP7_75t_R g4960 ( 
.A(n_4514),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4566),
.Y(n_4961)
);

CKINVDCx20_ASAP7_75t_R g4962 ( 
.A(n_4602),
.Y(n_4962)
);

HB1xp67_ASAP7_75t_L g4963 ( 
.A(n_4655),
.Y(n_4963)
);

CKINVDCx5p33_ASAP7_75t_R g4964 ( 
.A(n_4608),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_4621),
.Y(n_4965)
);

BUFx6f_ASAP7_75t_SL g4966 ( 
.A(n_4664),
.Y(n_4966)
);

CKINVDCx5p33_ASAP7_75t_R g4967 ( 
.A(n_4676),
.Y(n_4967)
);

CKINVDCx5p33_ASAP7_75t_R g4968 ( 
.A(n_4706),
.Y(n_4968)
);

INVxp67_ASAP7_75t_L g4969 ( 
.A(n_4675),
.Y(n_4969)
);

CKINVDCx16_ASAP7_75t_R g4970 ( 
.A(n_4693),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4568),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_4420),
.Y(n_4972)
);

HB1xp67_ASAP7_75t_L g4973 ( 
.A(n_4714),
.Y(n_4973)
);

CKINVDCx5p33_ASAP7_75t_R g4974 ( 
.A(n_4728),
.Y(n_4974)
);

CKINVDCx5p33_ASAP7_75t_R g4975 ( 
.A(n_4342),
.Y(n_4975)
);

CKINVDCx20_ASAP7_75t_R g4976 ( 
.A(n_4487),
.Y(n_4976)
);

INVx3_ASAP7_75t_L g4977 ( 
.A(n_4632),
.Y(n_4977)
);

CKINVDCx20_ASAP7_75t_R g4978 ( 
.A(n_4488),
.Y(n_4978)
);

HB1xp67_ASAP7_75t_L g4979 ( 
.A(n_4694),
.Y(n_4979)
);

CKINVDCx5p33_ASAP7_75t_R g4980 ( 
.A(n_4539),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_4599),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4569),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4570),
.Y(n_4983)
);

NOR2xp33_ASAP7_75t_L g4984 ( 
.A(n_4548),
.B(n_3981),
.Y(n_4984)
);

CKINVDCx20_ASAP7_75t_R g4985 ( 
.A(n_4391),
.Y(n_4985)
);

CKINVDCx5p33_ASAP7_75t_R g4986 ( 
.A(n_4332),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4724),
.B(n_3349),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4572),
.Y(n_4988)
);

CKINVDCx5p33_ASAP7_75t_R g4989 ( 
.A(n_4423),
.Y(n_4989)
);

CKINVDCx20_ASAP7_75t_R g4990 ( 
.A(n_4401),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_4500),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4574),
.Y(n_4992)
);

CKINVDCx5p33_ASAP7_75t_R g4993 ( 
.A(n_4426),
.Y(n_4993)
);

CKINVDCx5p33_ASAP7_75t_R g4994 ( 
.A(n_4454),
.Y(n_4994)
);

NOR2xp33_ASAP7_75t_L g4995 ( 
.A(n_4460),
.B(n_4001),
.Y(n_4995)
);

NOR2xp33_ASAP7_75t_L g4996 ( 
.A(n_4493),
.B(n_4004),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4575),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4576),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4582),
.Y(n_4999)
);

CKINVDCx5p33_ASAP7_75t_R g5000 ( 
.A(n_4311),
.Y(n_5000)
);

BUFx3_ASAP7_75t_L g5001 ( 
.A(n_4605),
.Y(n_5001)
);

INVxp67_ASAP7_75t_SL g5002 ( 
.A(n_4609),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4585),
.Y(n_5003)
);

CKINVDCx20_ASAP7_75t_R g5004 ( 
.A(n_4708),
.Y(n_5004)
);

INVx3_ASAP7_75t_L g5005 ( 
.A(n_4632),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4586),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4587),
.Y(n_5007)
);

CKINVDCx5p33_ASAP7_75t_R g5008 ( 
.A(n_4494),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_4610),
.Y(n_5009)
);

CKINVDCx20_ASAP7_75t_R g5010 ( 
.A(n_4448),
.Y(n_5010)
);

INVxp67_ASAP7_75t_SL g5011 ( 
.A(n_4618),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4588),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4589),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4590),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4591),
.Y(n_5015)
);

NOR2xp67_ASAP7_75t_L g5016 ( 
.A(n_4312),
.B(n_3458),
.Y(n_5016)
);

CKINVDCx5p33_ASAP7_75t_R g5017 ( 
.A(n_4597),
.Y(n_5017)
);

INVxp67_ASAP7_75t_SL g5018 ( 
.A(n_4601),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4592),
.Y(n_5019)
);

CKINVDCx20_ASAP7_75t_R g5020 ( 
.A(n_4604),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4593),
.Y(n_5021)
);

CKINVDCx20_ASAP7_75t_R g5022 ( 
.A(n_4607),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4594),
.Y(n_5023)
);

BUFx6f_ASAP7_75t_L g5024 ( 
.A(n_4674),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4614),
.B(n_4615),
.Y(n_5025)
);

CKINVDCx5p33_ASAP7_75t_R g5026 ( 
.A(n_4616),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4596),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_L g5028 ( 
.A(n_4326),
.B(n_4027),
.Y(n_5028)
);

CKINVDCx5p33_ASAP7_75t_R g5029 ( 
.A(n_4617),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4313),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4316),
.Y(n_5031)
);

CKINVDCx20_ASAP7_75t_R g5032 ( 
.A(n_4619),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4317),
.Y(n_5033)
);

INVxp67_ASAP7_75t_L g5034 ( 
.A(n_4623),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4318),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4321),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4322),
.Y(n_5037)
);

CKINVDCx20_ASAP7_75t_R g5038 ( 
.A(n_4624),
.Y(n_5038)
);

CKINVDCx5p33_ASAP7_75t_R g5039 ( 
.A(n_4625),
.Y(n_5039)
);

CKINVDCx5p33_ASAP7_75t_R g5040 ( 
.A(n_4627),
.Y(n_5040)
);

INVxp67_ASAP7_75t_SL g5041 ( 
.A(n_4629),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4329),
.Y(n_5042)
);

INVxp67_ASAP7_75t_L g5043 ( 
.A(n_4648),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4330),
.Y(n_5044)
);

CKINVDCx20_ASAP7_75t_R g5045 ( 
.A(n_4368),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4331),
.Y(n_5046)
);

CKINVDCx5p33_ASAP7_75t_R g5047 ( 
.A(n_4368),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_4368),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4357),
.B(n_4124),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4334),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4335),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4337),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4338),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4339),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_4368),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4631),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4633),
.Y(n_5057)
);

HB1xp67_ASAP7_75t_L g5058 ( 
.A(n_4674),
.Y(n_5058)
);

INVxp67_ASAP7_75t_SL g5059 ( 
.A(n_4695),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_4663),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4634),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_4397),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4663),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4636),
.Y(n_5064)
);

OR2x2_ASAP7_75t_L g5065 ( 
.A(n_4560),
.B(n_4164),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4637),
.Y(n_5066)
);

CKINVDCx5p33_ASAP7_75t_R g5067 ( 
.A(n_4663),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4638),
.Y(n_5068)
);

CKINVDCx5p33_ASAP7_75t_R g5069 ( 
.A(n_4663),
.Y(n_5069)
);

CKINVDCx5p33_ASAP7_75t_R g5070 ( 
.A(n_4695),
.Y(n_5070)
);

INVx2_ASAP7_75t_L g5071 ( 
.A(n_4439),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4640),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4641),
.Y(n_5073)
);

CKINVDCx20_ASAP7_75t_R g5074 ( 
.A(n_4642),
.Y(n_5074)
);

CKINVDCx5p33_ASAP7_75t_R g5075 ( 
.A(n_4635),
.Y(n_5075)
);

CKINVDCx20_ASAP7_75t_R g5076 ( 
.A(n_4643),
.Y(n_5076)
);

CKINVDCx5p33_ASAP7_75t_R g5077 ( 
.A(n_4667),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4646),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4649),
.Y(n_5079)
);

INVxp67_ASAP7_75t_SL g5080 ( 
.A(n_4506),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_4709),
.Y(n_5081)
);

INVxp67_ASAP7_75t_L g5082 ( 
.A(n_4717),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_4730),
.Y(n_5083)
);

CKINVDCx20_ASAP7_75t_R g5084 ( 
.A(n_4652),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4653),
.Y(n_5085)
);

BUFx3_ASAP7_75t_L g5086 ( 
.A(n_4656),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4657),
.Y(n_5087)
);

CKINVDCx5p33_ASAP7_75t_R g5088 ( 
.A(n_4660),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4662),
.Y(n_5089)
);

BUFx3_ASAP7_75t_L g5090 ( 
.A(n_4665),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4669),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4672),
.Y(n_5092)
);

INVxp33_ASAP7_75t_L g5093 ( 
.A(n_4647),
.Y(n_5093)
);

CKINVDCx20_ASAP7_75t_R g5094 ( 
.A(n_4677),
.Y(n_5094)
);

INVxp67_ASAP7_75t_SL g5095 ( 
.A(n_4702),
.Y(n_5095)
);

NOR2xp67_ASAP7_75t_L g5096 ( 
.A(n_4483),
.B(n_3499),
.Y(n_5096)
);

CKINVDCx5p33_ASAP7_75t_R g5097 ( 
.A(n_4680),
.Y(n_5097)
);

BUFx6f_ASAP7_75t_L g5098 ( 
.A(n_4449),
.Y(n_5098)
);

INVxp67_ASAP7_75t_L g5099 ( 
.A(n_4343),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_4681),
.Y(n_5100)
);

NOR2xp33_ASAP7_75t_L g5101 ( 
.A(n_4705),
.B(n_4030),
.Y(n_5101)
);

CKINVDCx20_ASAP7_75t_R g5102 ( 
.A(n_4682),
.Y(n_5102)
);

INVxp67_ASAP7_75t_SL g5103 ( 
.A(n_4684),
.Y(n_5103)
);

CKINVDCx5p33_ASAP7_75t_R g5104 ( 
.A(n_4688),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4689),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4692),
.Y(n_5106)
);

NOR2xp67_ASAP7_75t_L g5107 ( 
.A(n_4485),
.B(n_3535),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4697),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4348),
.Y(n_5109)
);

CKINVDCx5p33_ASAP7_75t_R g5110 ( 
.A(n_4699),
.Y(n_5110)
);

CKINVDCx20_ASAP7_75t_R g5111 ( 
.A(n_4700),
.Y(n_5111)
);

CKINVDCx5p33_ASAP7_75t_R g5112 ( 
.A(n_4701),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4703),
.Y(n_5113)
);

CKINVDCx5p33_ASAP7_75t_R g5114 ( 
.A(n_4707),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4710),
.Y(n_5115)
);

CKINVDCx20_ASAP7_75t_R g5116 ( 
.A(n_4711),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4713),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_4481),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4716),
.Y(n_5119)
);

CKINVDCx20_ASAP7_75t_R g5120 ( 
.A(n_4720),
.Y(n_5120)
);

CKINVDCx5p33_ASAP7_75t_R g5121 ( 
.A(n_4721),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4722),
.Y(n_5122)
);

CKINVDCx20_ASAP7_75t_R g5123 ( 
.A(n_4723),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4725),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_4729),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4731),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_4732),
.Y(n_5127)
);

CKINVDCx20_ASAP7_75t_R g5128 ( 
.A(n_4734),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_4351),
.B(n_3637),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_4352),
.Y(n_5130)
);

INVxp67_ASAP7_75t_SL g5131 ( 
.A(n_4718),
.Y(n_5131)
);

CKINVDCx20_ASAP7_75t_R g5132 ( 
.A(n_4354),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4355),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_4361),
.B(n_3692),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4362),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_4366),
.B(n_4367),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_4369),
.Y(n_5137)
);

INVxp67_ASAP7_75t_L g5138 ( 
.A(n_4370),
.Y(n_5138)
);

BUFx2_ASAP7_75t_L g5139 ( 
.A(n_4373),
.Y(n_5139)
);

CKINVDCx20_ASAP7_75t_R g5140 ( 
.A(n_4374),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4378),
.Y(n_5141)
);

BUFx10_ASAP7_75t_L g5142 ( 
.A(n_4379),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4380),
.Y(n_5143)
);

BUFx2_ASAP7_75t_L g5144 ( 
.A(n_4381),
.Y(n_5144)
);

CKINVDCx5p33_ASAP7_75t_R g5145 ( 
.A(n_4382),
.Y(n_5145)
);

CKINVDCx5p33_ASAP7_75t_R g5146 ( 
.A(n_4430),
.Y(n_5146)
);

CKINVDCx5p33_ASAP7_75t_R g5147 ( 
.A(n_4385),
.Y(n_5147)
);

CKINVDCx5p33_ASAP7_75t_R g5148 ( 
.A(n_4429),
.Y(n_5148)
);

CKINVDCx20_ASAP7_75t_R g5149 ( 
.A(n_4387),
.Y(n_5149)
);

CKINVDCx20_ASAP7_75t_R g5150 ( 
.A(n_4388),
.Y(n_5150)
);

INVxp67_ASAP7_75t_L g5151 ( 
.A(n_4389),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_4424),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4392),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4393),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4395),
.Y(n_5155)
);

INVxp67_ASAP7_75t_L g5156 ( 
.A(n_4396),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4398),
.Y(n_5157)
);

CKINVDCx20_ASAP7_75t_R g5158 ( 
.A(n_4399),
.Y(n_5158)
);

CKINVDCx16_ASAP7_75t_R g5159 ( 
.A(n_4400),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_4421),
.Y(n_5160)
);

BUFx6f_ASAP7_75t_L g5161 ( 
.A(n_4403),
.Y(n_5161)
);

INVxp67_ASAP7_75t_SL g5162 ( 
.A(n_4404),
.Y(n_5162)
);

CKINVDCx5p33_ASAP7_75t_R g5163 ( 
.A(n_4405),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4408),
.Y(n_5164)
);

CKINVDCx20_ASAP7_75t_R g5165 ( 
.A(n_4410),
.Y(n_5165)
);

BUFx6f_ASAP7_75t_SL g5166 ( 
.A(n_4413),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_4414),
.Y(n_5167)
);

NOR2xp33_ASAP7_75t_L g5168 ( 
.A(n_4416),
.B(n_4064),
.Y(n_5168)
);

CKINVDCx5p33_ASAP7_75t_R g5169 ( 
.A(n_4417),
.Y(n_5169)
);

CKINVDCx5p33_ASAP7_75t_R g5170 ( 
.A(n_4419),
.Y(n_5170)
);

CKINVDCx5p33_ASAP7_75t_R g5171 ( 
.A(n_4320),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4571),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_4320),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4571),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4571),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4571),
.Y(n_5176)
);

NOR2xp33_ASAP7_75t_L g5177 ( 
.A(n_4359),
.B(n_4073),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_4571),
.Y(n_5178)
);

CKINVDCx20_ASAP7_75t_R g5179 ( 
.A(n_4428),
.Y(n_5179)
);

CKINVDCx5p33_ASAP7_75t_R g5180 ( 
.A(n_4320),
.Y(n_5180)
);

INVxp67_ASAP7_75t_L g5181 ( 
.A(n_4440),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4571),
.Y(n_5182)
);

CKINVDCx5p33_ASAP7_75t_R g5183 ( 
.A(n_4320),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_4319),
.B(n_3702),
.Y(n_5184)
);

CKINVDCx5p33_ASAP7_75t_R g5185 ( 
.A(n_4320),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4571),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_4571),
.Y(n_5187)
);

CKINVDCx5p33_ASAP7_75t_R g5188 ( 
.A(n_4320),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4571),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4571),
.Y(n_5190)
);

HB1xp67_ASAP7_75t_L g5191 ( 
.A(n_4363),
.Y(n_5191)
);

CKINVDCx5p33_ASAP7_75t_R g5192 ( 
.A(n_4320),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_4571),
.Y(n_5193)
);

CKINVDCx5p33_ASAP7_75t_R g5194 ( 
.A(n_4320),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_4571),
.Y(n_5195)
);

BUFx2_ASAP7_75t_SL g5196 ( 
.A(n_4324),
.Y(n_5196)
);

CKINVDCx20_ASAP7_75t_R g5197 ( 
.A(n_4428),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_4571),
.Y(n_5198)
);

CKINVDCx5p33_ASAP7_75t_R g5199 ( 
.A(n_4320),
.Y(n_5199)
);

INVxp33_ASAP7_75t_SL g5200 ( 
.A(n_4310),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_4320),
.Y(n_5201)
);

CKINVDCx20_ASAP7_75t_R g5202 ( 
.A(n_4428),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4571),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4571),
.Y(n_5204)
);

CKINVDCx20_ASAP7_75t_R g5205 ( 
.A(n_4428),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4571),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4571),
.Y(n_5207)
);

NOR2xp67_ASAP7_75t_L g5208 ( 
.A(n_4412),
.B(n_3785),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4571),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_4571),
.Y(n_5210)
);

CKINVDCx20_ASAP7_75t_R g5211 ( 
.A(n_4428),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_4320),
.Y(n_5212)
);

CKINVDCx5p33_ASAP7_75t_R g5213 ( 
.A(n_4320),
.Y(n_5213)
);

CKINVDCx5p33_ASAP7_75t_R g5214 ( 
.A(n_4320),
.Y(n_5214)
);

CKINVDCx20_ASAP7_75t_R g5215 ( 
.A(n_4428),
.Y(n_5215)
);

CKINVDCx20_ASAP7_75t_R g5216 ( 
.A(n_4428),
.Y(n_5216)
);

CKINVDCx5p33_ASAP7_75t_R g5217 ( 
.A(n_4320),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_4571),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_4571),
.Y(n_5219)
);

NOR2xp33_ASAP7_75t_L g5220 ( 
.A(n_4359),
.B(n_4098),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_4571),
.Y(n_5221)
);

CKINVDCx5p33_ASAP7_75t_R g5222 ( 
.A(n_4320),
.Y(n_5222)
);

NOR2xp33_ASAP7_75t_R g5223 ( 
.A(n_4314),
.B(n_2921),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_4571),
.Y(n_5224)
);

CKINVDCx20_ASAP7_75t_R g5225 ( 
.A(n_4428),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4571),
.Y(n_5226)
);

CKINVDCx20_ASAP7_75t_R g5227 ( 
.A(n_4428),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_4571),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4571),
.Y(n_5229)
);

CKINVDCx20_ASAP7_75t_R g5230 ( 
.A(n_4428),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4571),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_4320),
.Y(n_5232)
);

INVxp67_ASAP7_75t_SL g5233 ( 
.A(n_4571),
.Y(n_5233)
);

CKINVDCx5p33_ASAP7_75t_R g5234 ( 
.A(n_4320),
.Y(n_5234)
);

INVxp67_ASAP7_75t_SL g5235 ( 
.A(n_4571),
.Y(n_5235)
);

NOR2xp33_ASAP7_75t_L g5236 ( 
.A(n_5093),
.B(n_4136),
.Y(n_5236)
);

NAND2xp5_ASAP7_75t_L g5237 ( 
.A(n_5047),
.B(n_3786),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_SL g5238 ( 
.A(n_4972),
.B(n_4190),
.Y(n_5238)
);

NOR2xp33_ASAP7_75t_L g5239 ( 
.A(n_4741),
.B(n_5131),
.Y(n_5239)
);

BUFx6f_ASAP7_75t_L g5240 ( 
.A(n_4784),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_5048),
.B(n_3991),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5098),
.Y(n_5242)
);

AND2x4_ASAP7_75t_L g5243 ( 
.A(n_4768),
.B(n_4049),
.Y(n_5243)
);

BUFx6f_ASAP7_75t_L g5244 ( 
.A(n_4784),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5058),
.Y(n_5245)
);

CKINVDCx5p33_ASAP7_75t_R g5246 ( 
.A(n_4763),
.Y(n_5246)
);

INVxp67_ASAP7_75t_L g5247 ( 
.A(n_5065),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_5098),
.Y(n_5248)
);

NAND2xp5_ASAP7_75t_L g5249 ( 
.A(n_5055),
.B(n_4051),
.Y(n_5249)
);

INVx3_ASAP7_75t_L g5250 ( 
.A(n_4784),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5060),
.B(n_4134),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_5098),
.Y(n_5252)
);

BUFx6f_ASAP7_75t_L g5253 ( 
.A(n_4868),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5001),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5159),
.B(n_3509),
.Y(n_5255)
);

BUFx3_ASAP7_75t_L g5256 ( 
.A(n_5070),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_4764),
.Y(n_5257)
);

CKINVDCx11_ASAP7_75t_R g5258 ( 
.A(n_4861),
.Y(n_5258)
);

OAI22xp5_ASAP7_75t_SL g5259 ( 
.A1(n_5010),
.A2(n_3243),
.B1(n_3462),
.B2(n_3051),
.Y(n_5259)
);

BUFx6f_ASAP7_75t_L g5260 ( 
.A(n_4868),
.Y(n_5260)
);

INVx3_ASAP7_75t_L g5261 ( 
.A(n_4868),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5136),
.Y(n_5262)
);

BUFx6f_ASAP7_75t_L g5263 ( 
.A(n_5024),
.Y(n_5263)
);

NOR2x1_ASAP7_75t_L g5264 ( 
.A(n_5045),
.B(n_3030),
.Y(n_5264)
);

XOR2xp5_ASAP7_75t_L g5265 ( 
.A(n_4737),
.B(n_3176),
.Y(n_5265)
);

AND2x4_ASAP7_75t_L g5266 ( 
.A(n_4746),
.B(n_4139),
.Y(n_5266)
);

BUFx12f_ASAP7_75t_L g5267 ( 
.A(n_4953),
.Y(n_5267)
);

BUFx6f_ASAP7_75t_L g5268 ( 
.A(n_5024),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5056),
.Y(n_5269)
);

INVx3_ASAP7_75t_L g5270 ( 
.A(n_5024),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_5071),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5057),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_5061),
.Y(n_5273)
);

CKINVDCx5p33_ASAP7_75t_R g5274 ( 
.A(n_4771),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_5064),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5066),
.Y(n_5276)
);

BUFx6f_ASAP7_75t_L g5277 ( 
.A(n_4745),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_5068),
.Y(n_5278)
);

OAI22xp5_ASAP7_75t_L g5279 ( 
.A1(n_5082),
.A2(n_4223),
.B1(n_4224),
.B2(n_4204),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_5118),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5072),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4750),
.Y(n_5282)
);

OAI21x1_ASAP7_75t_L g5283 ( 
.A1(n_4736),
.A2(n_3146),
.B(n_3120),
.Y(n_5283)
);

BUFx3_ASAP7_75t_L g5284 ( 
.A(n_4975),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_4822),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5073),
.Y(n_5286)
);

INVx3_ASAP7_75t_L g5287 ( 
.A(n_4745),
.Y(n_5287)
);

CKINVDCx5p33_ASAP7_75t_R g5288 ( 
.A(n_4773),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_5063),
.B(n_4200),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5078),
.Y(n_5290)
);

INVx2_ASAP7_75t_L g5291 ( 
.A(n_4824),
.Y(n_5291)
);

AND2x4_ASAP7_75t_L g5292 ( 
.A(n_4761),
.B(n_3154),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5079),
.Y(n_5293)
);

OR2x2_ASAP7_75t_L g5294 ( 
.A(n_4845),
.B(n_3861),
.Y(n_5294)
);

AOI22xp5_ASAP7_75t_L g5295 ( 
.A1(n_4814),
.A2(n_2951),
.B1(n_2965),
.B2(n_2933),
.Y(n_5295)
);

INVx2_ASAP7_75t_L g5296 ( 
.A(n_4843),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5085),
.Y(n_5297)
);

OA21x2_ASAP7_75t_L g5298 ( 
.A1(n_5067),
.A2(n_3174),
.B(n_3155),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_5062),
.Y(n_5299)
);

INVx3_ASAP7_75t_L g5300 ( 
.A(n_4745),
.Y(n_5300)
);

INVx2_ASAP7_75t_L g5301 ( 
.A(n_4884),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5087),
.Y(n_5302)
);

AND2x4_ASAP7_75t_L g5303 ( 
.A(n_4956),
.B(n_3181),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_5089),
.Y(n_5304)
);

INVx2_ASAP7_75t_L g5305 ( 
.A(n_4932),
.Y(n_5305)
);

BUFx6f_ASAP7_75t_L g5306 ( 
.A(n_5161),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_4952),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_5049),
.B(n_3519),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5091),
.Y(n_5309)
);

BUFx3_ASAP7_75t_L g5310 ( 
.A(n_5086),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_5092),
.Y(n_5311)
);

INVx3_ASAP7_75t_L g5312 ( 
.A(n_4977),
.Y(n_5312)
);

AND2x2_ASAP7_75t_L g5313 ( 
.A(n_5101),
.B(n_3519),
.Y(n_5313)
);

HB1xp67_ASAP7_75t_L g5314 ( 
.A(n_4853),
.Y(n_5314)
);

BUFx6f_ASAP7_75t_L g5315 ( 
.A(n_5161),
.Y(n_5315)
);

BUFx6f_ASAP7_75t_L g5316 ( 
.A(n_5161),
.Y(n_5316)
);

BUFx6f_ASAP7_75t_L g5317 ( 
.A(n_4977),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_4955),
.Y(n_5318)
);

BUFx2_ASAP7_75t_L g5319 ( 
.A(n_4886),
.Y(n_5319)
);

NAND2xp5_ASAP7_75t_L g5320 ( 
.A(n_5069),
.B(n_3156),
.Y(n_5320)
);

AND2x2_ASAP7_75t_L g5321 ( 
.A(n_5043),
.B(n_3525),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5008),
.B(n_3525),
.Y(n_5322)
);

AND2x4_ASAP7_75t_L g5323 ( 
.A(n_4770),
.B(n_4801),
.Y(n_5323)
);

AND2x6_ASAP7_75t_L g5324 ( 
.A(n_4945),
.B(n_2983),
.Y(n_5324)
);

BUFx8_ASAP7_75t_L g5325 ( 
.A(n_4966),
.Y(n_5325)
);

AND2x2_ASAP7_75t_L g5326 ( 
.A(n_5028),
.B(n_3526),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_4749),
.A2(n_3185),
.B(n_3175),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5105),
.Y(n_5328)
);

CKINVDCx5p33_ASAP7_75t_R g5329 ( 
.A(n_4774),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5106),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5108),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5113),
.Y(n_5332)
);

AND2x6_ASAP7_75t_L g5333 ( 
.A(n_4849),
.B(n_4760),
.Y(n_5333)
);

AND2x2_ASAP7_75t_L g5334 ( 
.A(n_5080),
.B(n_3526),
.Y(n_5334)
);

INVx2_ASAP7_75t_L g5335 ( 
.A(n_4777),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_5233),
.B(n_3197),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5115),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_4778),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5117),
.Y(n_5339)
);

AND2x2_ASAP7_75t_L g5340 ( 
.A(n_5095),
.B(n_3547),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_5119),
.Y(n_5341)
);

OR2x2_ASAP7_75t_L g5342 ( 
.A(n_5184),
.B(n_2989),
.Y(n_5342)
);

BUFx6f_ASAP7_75t_L g5343 ( 
.A(n_5005),
.Y(n_5343)
);

BUFx2_ASAP7_75t_L g5344 ( 
.A(n_4888),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5122),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_L g5346 ( 
.A(n_5235),
.B(n_3205),
.Y(n_5346)
);

BUFx6f_ASAP7_75t_L g5347 ( 
.A(n_5005),
.Y(n_5347)
);

INVx3_ASAP7_75t_L g5348 ( 
.A(n_4752),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_5124),
.Y(n_5349)
);

INVx2_ASAP7_75t_L g5350 ( 
.A(n_4780),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_4785),
.Y(n_5351)
);

BUFx6f_ASAP7_75t_L g5352 ( 
.A(n_4752),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_SL g5353 ( 
.A1(n_4985),
.A2(n_3650),
.B1(n_3651),
.B2(n_3494),
.Y(n_5353)
);

INVx2_ASAP7_75t_L g5354 ( 
.A(n_4790),
.Y(n_5354)
);

NOR2xp33_ASAP7_75t_SL g5355 ( 
.A(n_4941),
.B(n_3683),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5030),
.B(n_3216),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5126),
.Y(n_5357)
);

AND2x2_ASAP7_75t_L g5358 ( 
.A(n_4819),
.B(n_3547),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5031),
.B(n_3245),
.Y(n_5359)
);

HB1xp67_ASAP7_75t_L g5360 ( 
.A(n_5000),
.Y(n_5360)
);

BUFx6f_ASAP7_75t_L g5361 ( 
.A(n_5090),
.Y(n_5361)
);

INVx6_ASAP7_75t_L g5362 ( 
.A(n_5142),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_L g5363 ( 
.A(n_5033),
.B(n_3258),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5127),
.Y(n_5364)
);

BUFx8_ASAP7_75t_SL g5365 ( 
.A(n_4865),
.Y(n_5365)
);

AND2x4_ASAP7_75t_L g5366 ( 
.A(n_4816),
.B(n_3182),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_5035),
.B(n_3264),
.Y(n_5367)
);

AND2x6_ASAP7_75t_L g5368 ( 
.A(n_5177),
.B(n_3019),
.Y(n_5368)
);

HB1xp67_ASAP7_75t_L g5369 ( 
.A(n_4993),
.Y(n_5369)
);

INVxp67_ASAP7_75t_L g5370 ( 
.A(n_4979),
.Y(n_5370)
);

OAI22xp5_ASAP7_75t_SL g5371 ( 
.A1(n_4990),
.A2(n_3858),
.B1(n_3894),
.B2(n_3778),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5036),
.B(n_3274),
.Y(n_5372)
);

BUFx6f_ASAP7_75t_L g5373 ( 
.A(n_5155),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5130),
.Y(n_5374)
);

INVx2_ASAP7_75t_L g5375 ( 
.A(n_4791),
.Y(n_5375)
);

OAI21x1_ASAP7_75t_L g5376 ( 
.A1(n_5037),
.A2(n_3405),
.B(n_3359),
.Y(n_5376)
);

INVx5_ASAP7_75t_L g5377 ( 
.A(n_4847),
.Y(n_5377)
);

BUFx3_ASAP7_75t_L g5378 ( 
.A(n_5139),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5133),
.Y(n_5379)
);

BUFx6f_ASAP7_75t_L g5380 ( 
.A(n_4748),
.Y(n_5380)
);

CKINVDCx20_ASAP7_75t_R g5381 ( 
.A(n_4743),
.Y(n_5381)
);

INVx3_ASAP7_75t_L g5382 ( 
.A(n_5142),
.Y(n_5382)
);

AND2x4_ASAP7_75t_L g5383 ( 
.A(n_4821),
.B(n_3183),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5135),
.Y(n_5384)
);

AND2x4_ASAP7_75t_L g5385 ( 
.A(n_4823),
.B(n_3186),
.Y(n_5385)
);

BUFx6f_ASAP7_75t_L g5386 ( 
.A(n_4765),
.Y(n_5386)
);

NAND2xp5_ASAP7_75t_SL g5387 ( 
.A(n_5208),
.B(n_2924),
.Y(n_5387)
);

HB1xp67_ASAP7_75t_L g5388 ( 
.A(n_4994),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_4794),
.Y(n_5389)
);

AND2x2_ASAP7_75t_SL g5390 ( 
.A(n_4852),
.B(n_3406),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_SL g5391 ( 
.A(n_4980),
.B(n_2925),
.Y(n_5391)
);

CKINVDCx5p33_ASAP7_75t_R g5392 ( 
.A(n_4779),
.Y(n_5392)
);

NAND2xp5_ASAP7_75t_L g5393 ( 
.A(n_5042),
.B(n_3424),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4800),
.Y(n_5394)
);

AND2x4_ASAP7_75t_L g5395 ( 
.A(n_4837),
.B(n_3189),
.Y(n_5395)
);

OAI22xp5_ASAP7_75t_L g5396 ( 
.A1(n_4867),
.A2(n_2932),
.B1(n_2936),
.B2(n_2927),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_5137),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_4804),
.Y(n_5398)
);

INVx3_ASAP7_75t_L g5399 ( 
.A(n_4766),
.Y(n_5399)
);

BUFx6f_ASAP7_75t_L g5400 ( 
.A(n_4767),
.Y(n_5400)
);

AOI22x1_ASAP7_75t_L g5401 ( 
.A1(n_4878),
.A2(n_2941),
.B1(n_2942),
.B2(n_2940),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5141),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_4782),
.Y(n_5403)
);

AND2x4_ASAP7_75t_L g5404 ( 
.A(n_4842),
.B(n_3195),
.Y(n_5404)
);

AND2x2_ASAP7_75t_L g5405 ( 
.A(n_4947),
.B(n_3603),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_L g5406 ( 
.A(n_5044),
.B(n_3457),
.Y(n_5406)
);

OAI22xp5_ASAP7_75t_L g5407 ( 
.A1(n_4830),
.A2(n_4909),
.B1(n_4929),
.B2(n_4879),
.Y(n_5407)
);

AND2x2_ASAP7_75t_L g5408 ( 
.A(n_4802),
.B(n_3603),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5143),
.Y(n_5409)
);

AND2x4_ASAP7_75t_L g5410 ( 
.A(n_4844),
.B(n_3214),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5153),
.Y(n_5411)
);

AND2x2_ASAP7_75t_L g5412 ( 
.A(n_4809),
.B(n_3661),
.Y(n_5412)
);

AND2x6_ASAP7_75t_L g5413 ( 
.A(n_5220),
.B(n_3048),
.Y(n_5413)
);

INVx1_ASAP7_75t_SL g5414 ( 
.A(n_4976),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5154),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5157),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5164),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5167),
.Y(n_5418)
);

BUFx2_ASAP7_75t_L g5419 ( 
.A(n_4978),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_4805),
.Y(n_5420)
);

BUFx6f_ASAP7_75t_L g5421 ( 
.A(n_4772),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5002),
.Y(n_5422)
);

OAI22xp5_ASAP7_75t_L g5423 ( 
.A1(n_4940),
.A2(n_2945),
.B1(n_2946),
.B2(n_2944),
.Y(n_5423)
);

AOI22xp5_ASAP7_75t_L g5424 ( 
.A1(n_4996),
.A2(n_3080),
.B1(n_3089),
.B2(n_3052),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5011),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_4807),
.Y(n_5426)
);

BUFx3_ASAP7_75t_L g5427 ( 
.A(n_5144),
.Y(n_5427)
);

OR2x6_ASAP7_75t_L g5428 ( 
.A(n_5196),
.B(n_3102),
.Y(n_5428)
);

INVx4_ASAP7_75t_L g5429 ( 
.A(n_5017),
.Y(n_5429)
);

BUFx6f_ASAP7_75t_L g5430 ( 
.A(n_4742),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5046),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_4811),
.Y(n_5432)
);

INVx2_ASAP7_75t_L g5433 ( 
.A(n_4812),
.Y(n_5433)
);

OA21x2_ASAP7_75t_L g5434 ( 
.A1(n_5050),
.A2(n_3224),
.B(n_3221),
.Y(n_5434)
);

AND2x4_ASAP7_75t_L g5435 ( 
.A(n_4889),
.B(n_3233),
.Y(n_5435)
);

INVx3_ASAP7_75t_L g5436 ( 
.A(n_5051),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_4896),
.A2(n_3108),
.B1(n_3161),
.B2(n_3096),
.Y(n_5437)
);

BUFx3_ASAP7_75t_L g5438 ( 
.A(n_4740),
.Y(n_5438)
);

OAI22xp5_ASAP7_75t_SL g5439 ( 
.A1(n_4841),
.A2(n_4247),
.B1(n_4138),
.B2(n_3202),
.Y(n_5439)
);

AOI22xp5_ASAP7_75t_L g5440 ( 
.A1(n_5020),
.A2(n_3353),
.B1(n_3407),
.B2(n_3200),
.Y(n_5440)
);

BUFx6f_ASAP7_75t_L g5441 ( 
.A(n_4813),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_L g5442 ( 
.A(n_5052),
.B(n_5053),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5054),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5059),
.Y(n_5444)
);

BUFx8_ASAP7_75t_L g5445 ( 
.A(n_4966),
.Y(n_5445)
);

BUFx6f_ASAP7_75t_L g5446 ( 
.A(n_4817),
.Y(n_5446)
);

BUFx6f_ASAP7_75t_L g5447 ( 
.A(n_4820),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5109),
.Y(n_5448)
);

BUFx6f_ASAP7_75t_L g5449 ( 
.A(n_4825),
.Y(n_5449)
);

BUFx6f_ASAP7_75t_L g5450 ( 
.A(n_4826),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_4831),
.Y(n_5451)
);

INVx3_ASAP7_75t_L g5452 ( 
.A(n_5172),
.Y(n_5452)
);

OAI22xp5_ASAP7_75t_L g5453 ( 
.A1(n_4995),
.A2(n_2955),
.B1(n_2957),
.B2(n_2952),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_4834),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_4835),
.Y(n_5455)
);

BUFx6f_ASAP7_75t_L g5456 ( 
.A(n_4838),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_4848),
.Y(n_5457)
);

AND2x4_ASAP7_75t_L g5458 ( 
.A(n_4855),
.B(n_3234),
.Y(n_5458)
);

INVx3_ASAP7_75t_L g5459 ( 
.A(n_5174),
.Y(n_5459)
);

INVx3_ASAP7_75t_L g5460 ( 
.A(n_5175),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5176),
.Y(n_5461)
);

NAND2xp5_ASAP7_75t_L g5462 ( 
.A(n_5178),
.B(n_3498),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_5182),
.B(n_3503),
.Y(n_5463)
);

BUFx6f_ASAP7_75t_L g5464 ( 
.A(n_4851),
.Y(n_5464)
);

OAI21x1_ASAP7_75t_L g5465 ( 
.A1(n_5186),
.A2(n_3594),
.B(n_3577),
.Y(n_5465)
);

INVx3_ASAP7_75t_L g5466 ( 
.A(n_5187),
.Y(n_5466)
);

OAI22xp5_ASAP7_75t_SL g5467 ( 
.A1(n_4850),
.A2(n_3215),
.B1(n_3242),
.B2(n_3204),
.Y(n_5467)
);

OAI22xp5_ASAP7_75t_SL g5468 ( 
.A1(n_4854),
.A2(n_3249),
.B1(n_3279),
.B2(n_3248),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5181),
.B(n_3661),
.Y(n_5469)
);

BUFx6f_ASAP7_75t_L g5470 ( 
.A(n_4856),
.Y(n_5470)
);

NAND2xp5_ASAP7_75t_L g5471 ( 
.A(n_5189),
.B(n_3612),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5190),
.Y(n_5472)
);

INVx2_ASAP7_75t_L g5473 ( 
.A(n_4858),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5193),
.Y(n_5474)
);

INVx4_ASAP7_75t_L g5475 ( 
.A(n_5026),
.Y(n_5475)
);

AND2x2_ASAP7_75t_L g5476 ( 
.A(n_4958),
.B(n_3663),
.Y(n_5476)
);

AND2x4_ASAP7_75t_L g5477 ( 
.A(n_4857),
.B(n_3238),
.Y(n_5477)
);

CKINVDCx5p33_ASAP7_75t_R g5478 ( 
.A(n_4787),
.Y(n_5478)
);

AND2x4_ASAP7_75t_L g5479 ( 
.A(n_5162),
.B(n_3241),
.Y(n_5479)
);

INVx2_ASAP7_75t_L g5480 ( 
.A(n_4862),
.Y(n_5480)
);

BUFx3_ASAP7_75t_L g5481 ( 
.A(n_5195),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5198),
.B(n_3615),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5203),
.A2(n_3690),
.B(n_3644),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5204),
.B(n_3731),
.Y(n_5484)
);

NOR2xp33_ASAP7_75t_L g5485 ( 
.A(n_5206),
.B(n_2960),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_4863),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5207),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5209),
.Y(n_5488)
);

HB1xp67_ASAP7_75t_L g5489 ( 
.A(n_4963),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5210),
.Y(n_5490)
);

OAI22xp5_ASAP7_75t_SL g5491 ( 
.A1(n_4859),
.A2(n_3322),
.B1(n_3323),
.B2(n_3320),
.Y(n_5491)
);

BUFx3_ASAP7_75t_L g5492 ( 
.A(n_5218),
.Y(n_5492)
);

BUFx12f_ASAP7_75t_L g5493 ( 
.A(n_4959),
.Y(n_5493)
);

AND2x6_ASAP7_75t_L g5494 ( 
.A(n_4918),
.B(n_3408),
.Y(n_5494)
);

INVx4_ASAP7_75t_L g5495 ( 
.A(n_5029),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5219),
.Y(n_5496)
);

BUFx2_ASAP7_75t_L g5497 ( 
.A(n_4871),
.Y(n_5497)
);

BUFx6f_ASAP7_75t_L g5498 ( 
.A(n_4866),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5221),
.Y(n_5499)
);

AND2x4_ASAP7_75t_L g5500 ( 
.A(n_5103),
.B(n_3255),
.Y(n_5500)
);

BUFx3_ASAP7_75t_L g5501 ( 
.A(n_5224),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_5226),
.B(n_3746),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5228),
.Y(n_5503)
);

AND2x2_ASAP7_75t_SL g5504 ( 
.A(n_4755),
.B(n_3755),
.Y(n_5504)
);

OAI21x1_ASAP7_75t_L g5505 ( 
.A1(n_5229),
.A2(n_3830),
.B(n_3817),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_4984),
.B(n_3663),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_5231),
.B(n_3865),
.Y(n_5507)
);

INVx4_ASAP7_75t_L g5508 ( 
.A(n_5039),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_SL g5509 ( 
.A(n_4981),
.B(n_2961),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_4869),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_4872),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_4873),
.Y(n_5512)
);

NOR2xp33_ASAP7_75t_L g5513 ( 
.A(n_5040),
.B(n_2962),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_R g5514 ( 
.A(n_4829),
.B(n_3361),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_4875),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_4876),
.Y(n_5516)
);

BUFx6f_ASAP7_75t_L g5517 ( 
.A(n_4877),
.Y(n_5517)
);

INVx3_ASAP7_75t_L g5518 ( 
.A(n_5009),
.Y(n_5518)
);

INVx3_ASAP7_75t_L g5519 ( 
.A(n_4880),
.Y(n_5519)
);

NOR2xp33_ASAP7_75t_L g5520 ( 
.A(n_4753),
.B(n_4788),
.Y(n_5520)
);

AND2x4_ASAP7_75t_L g5521 ( 
.A(n_5018),
.B(n_3261),
.Y(n_5521)
);

OAI22xp5_ASAP7_75t_SL g5522 ( 
.A1(n_4839),
.A2(n_3451),
.B1(n_3474),
.B2(n_3402),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_L g5523 ( 
.A(n_5041),
.B(n_3873),
.Y(n_5523)
);

BUFx2_ASAP7_75t_L g5524 ( 
.A(n_4874),
.Y(n_5524)
);

HB1xp67_ASAP7_75t_L g5525 ( 
.A(n_4973),
.Y(n_5525)
);

CKINVDCx5p33_ASAP7_75t_R g5526 ( 
.A(n_4789),
.Y(n_5526)
);

AND2x6_ASAP7_75t_L g5527 ( 
.A(n_4918),
.B(n_3441),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5088),
.B(n_3874),
.Y(n_5528)
);

INVx3_ASAP7_75t_L g5529 ( 
.A(n_4882),
.Y(n_5529)
);

INVx3_ASAP7_75t_L g5530 ( 
.A(n_4885),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_4898),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_4899),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_4900),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_4902),
.Y(n_5534)
);

INVx2_ASAP7_75t_L g5535 ( 
.A(n_4903),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_4904),
.Y(n_5536)
);

INVx2_ASAP7_75t_L g5537 ( 
.A(n_4905),
.Y(n_5537)
);

INVx2_ASAP7_75t_SL g5538 ( 
.A(n_4974),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_4910),
.Y(n_5539)
);

INVx4_ASAP7_75t_L g5540 ( 
.A(n_5075),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_4912),
.Y(n_5541)
);

AND2x2_ASAP7_75t_L g5542 ( 
.A(n_5145),
.B(n_3902),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_4915),
.Y(n_5543)
);

BUFx2_ASAP7_75t_L g5544 ( 
.A(n_4883),
.Y(n_5544)
);

NOR2x1_ASAP7_75t_L g5545 ( 
.A(n_5025),
.B(n_3263),
.Y(n_5545)
);

CKINVDCx6p67_ASAP7_75t_R g5546 ( 
.A(n_4890),
.Y(n_5546)
);

OAI22x1_ASAP7_75t_L g5547 ( 
.A1(n_4986),
.A2(n_3699),
.B1(n_3705),
.B2(n_3486),
.Y(n_5547)
);

AND2x2_ASAP7_75t_L g5548 ( 
.A(n_5146),
.B(n_3902),
.Y(n_5548)
);

BUFx6f_ASAP7_75t_L g5549 ( 
.A(n_4917),
.Y(n_5549)
);

BUFx3_ASAP7_75t_L g5550 ( 
.A(n_4893),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_4921),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_4924),
.Y(n_5552)
);

BUFx2_ASAP7_75t_L g5553 ( 
.A(n_5223),
.Y(n_5553)
);

BUFx6f_ASAP7_75t_L g5554 ( 
.A(n_4925),
.Y(n_5554)
);

INVx3_ASAP7_75t_L g5555 ( 
.A(n_4931),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_4938),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4942),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_4950),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_4957),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4961),
.Y(n_5560)
);

HB1xp67_ASAP7_75t_L g5561 ( 
.A(n_4951),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_4971),
.Y(n_5562)
);

BUFx2_ASAP7_75t_L g5563 ( 
.A(n_5004),
.Y(n_5563)
);

INVx2_ASAP7_75t_SL g5564 ( 
.A(n_4989),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_5097),
.B(n_3926),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_SL g5566 ( 
.A(n_4991),
.B(n_2963),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_4982),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_4983),
.Y(n_5568)
);

INVx2_ASAP7_75t_L g5569 ( 
.A(n_4988),
.Y(n_5569)
);

INVx3_ASAP7_75t_L g5570 ( 
.A(n_4992),
.Y(n_5570)
);

INVx3_ASAP7_75t_L g5571 ( 
.A(n_4997),
.Y(n_5571)
);

AND2x2_ASAP7_75t_L g5572 ( 
.A(n_5147),
.B(n_5148),
.Y(n_5572)
);

AOI22xp5_ASAP7_75t_L g5573 ( 
.A1(n_5022),
.A2(n_3792),
.B1(n_3800),
.B2(n_3753),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_5100),
.B(n_3940),
.Y(n_5574)
);

INVx2_ASAP7_75t_L g5575 ( 
.A(n_4998),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_4999),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_5003),
.Y(n_5577)
);

OA21x2_ASAP7_75t_L g5578 ( 
.A1(n_4887),
.A2(n_3270),
.B(n_3268),
.Y(n_5578)
);

INVx3_ASAP7_75t_L g5579 ( 
.A(n_5006),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5007),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_L g5581 ( 
.A(n_5104),
.B(n_3948),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5012),
.Y(n_5582)
);

OAI21x1_ASAP7_75t_L g5583 ( 
.A1(n_4987),
.A2(n_4012),
.B(n_3969),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_5013),
.Y(n_5584)
);

OAI21x1_ASAP7_75t_L g5585 ( 
.A1(n_5129),
.A2(n_4019),
.B(n_4018),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5110),
.B(n_4020),
.Y(n_5586)
);

INVx5_ASAP7_75t_L g5587 ( 
.A(n_4970),
.Y(n_5587)
);

AND2x2_ASAP7_75t_L g5588 ( 
.A(n_5152),
.B(n_3986),
.Y(n_5588)
);

INVx3_ASAP7_75t_L g5589 ( 
.A(n_5014),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5015),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5019),
.Y(n_5591)
);

INVx5_ASAP7_75t_L g5592 ( 
.A(n_4930),
.Y(n_5592)
);

BUFx6f_ASAP7_75t_L g5593 ( 
.A(n_5021),
.Y(n_5593)
);

INVx1_ASAP7_75t_SL g5594 ( 
.A(n_4754),
.Y(n_5594)
);

OAI22xp5_ASAP7_75t_L g5595 ( 
.A1(n_5160),
.A2(n_2966),
.B1(n_2967),
.B2(n_2964),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5023),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5027),
.Y(n_5597)
);

INVx2_ASAP7_75t_L g5598 ( 
.A(n_5077),
.Y(n_5598)
);

BUFx6f_ASAP7_75t_L g5599 ( 
.A(n_5134),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5081),
.Y(n_5600)
);

OAI22xp5_ASAP7_75t_L g5601 ( 
.A1(n_5163),
.A2(n_2971),
.B1(n_2973),
.B2(n_2969),
.Y(n_5601)
);

BUFx6f_ASAP7_75t_L g5602 ( 
.A(n_5083),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5099),
.Y(n_5603)
);

CKINVDCx5p33_ASAP7_75t_R g5604 ( 
.A(n_4792),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_5169),
.B(n_3986),
.Y(n_5605)
);

CKINVDCx5p33_ASAP7_75t_R g5606 ( 
.A(n_4797),
.Y(n_5606)
);

AOI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_5032),
.A2(n_3958),
.B1(n_3966),
.B2(n_3913),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_L g5608 ( 
.A(n_5112),
.B(n_5114),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5138),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_5151),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_5156),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5034),
.Y(n_5612)
);

NAND2xp33_ASAP7_75t_L g5613 ( 
.A(n_5121),
.B(n_2979),
.Y(n_5613)
);

AND2x2_ASAP7_75t_SL g5614 ( 
.A(n_4775),
.B(n_4024),
.Y(n_5614)
);

AOI22xp5_ASAP7_75t_L g5615 ( 
.A1(n_5038),
.A2(n_4011),
.B1(n_4043),
.B2(n_4007),
.Y(n_5615)
);

CKINVDCx5p33_ASAP7_75t_R g5616 ( 
.A(n_4798),
.Y(n_5616)
);

OA21x2_ASAP7_75t_L g5617 ( 
.A1(n_5016),
.A2(n_3277),
.B(n_3273),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_5125),
.B(n_4055),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_5170),
.Y(n_5619)
);

OAI22xp5_ASAP7_75t_L g5620 ( 
.A1(n_5074),
.A2(n_2984),
.B1(n_2992),
.B2(n_2981),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5076),
.Y(n_5621)
);

AND2x4_ASAP7_75t_L g5622 ( 
.A(n_4943),
.B(n_3280),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5168),
.B(n_4067),
.Y(n_5623)
);

AOI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_5084),
.A2(n_4131),
.B1(n_4180),
.B2(n_4115),
.Y(n_5624)
);

INVx2_ASAP7_75t_L g5625 ( 
.A(n_5166),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5166),
.Y(n_5626)
);

NOR2x1_ASAP7_75t_L g5627 ( 
.A(n_4954),
.B(n_3281),
.Y(n_5627)
);

AND2x2_ASAP7_75t_L g5628 ( 
.A(n_4891),
.B(n_4120),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5094),
.Y(n_5629)
);

HB1xp67_ASAP7_75t_L g5630 ( 
.A(n_4969),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_5102),
.Y(n_5631)
);

BUFx3_ASAP7_75t_L g5632 ( 
.A(n_4894),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5111),
.Y(n_5633)
);

AND2x4_ASAP7_75t_L g5634 ( 
.A(n_5132),
.B(n_3284),
.Y(n_5634)
);

BUFx6f_ASAP7_75t_L g5635 ( 
.A(n_4808),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5116),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5140),
.B(n_3286),
.Y(n_5637)
);

AND2x6_ASAP7_75t_L g5638 ( 
.A(n_4803),
.B(n_4261),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_5096),
.B(n_4071),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5107),
.B(n_4097),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_5120),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_4827),
.B(n_4108),
.Y(n_5642)
);

OAI22xp5_ASAP7_75t_L g5643 ( 
.A1(n_5123),
.A2(n_2994),
.B1(n_2995),
.B2(n_2993),
.Y(n_5643)
);

AND2x6_ASAP7_75t_L g5644 ( 
.A(n_4786),
.B(n_4294),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5128),
.Y(n_5645)
);

HB1xp67_ASAP7_75t_L g5646 ( 
.A(n_5149),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5150),
.Y(n_5647)
);

HB1xp67_ASAP7_75t_L g5648 ( 
.A(n_5158),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_5165),
.Y(n_5649)
);

BUFx6f_ASAP7_75t_L g5650 ( 
.A(n_4828),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_4913),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_4920),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_4936),
.Y(n_5653)
);

NAND2xp5_ASAP7_75t_L g5654 ( 
.A(n_4836),
.B(n_4113),
.Y(n_5654)
);

OAI21x1_ASAP7_75t_L g5655 ( 
.A1(n_4757),
.A2(n_4206),
.B(n_4145),
.Y(n_5655)
);

AND2x4_ASAP7_75t_L g5656 ( 
.A(n_4759),
.B(n_3290),
.Y(n_5656)
);

AND2x2_ASAP7_75t_L g5657 ( 
.A(n_4840),
.B(n_4120),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_4846),
.B(n_4860),
.Y(n_5658)
);

BUFx6f_ASAP7_75t_L g5659 ( 
.A(n_4864),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_4769),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_4870),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_4783),
.Y(n_5662)
);

AND2x2_ASAP7_75t_L g5663 ( 
.A(n_4881),
.B(n_4284),
.Y(n_5663)
);

INVx3_ASAP7_75t_L g5664 ( 
.A(n_4892),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_4799),
.Y(n_5665)
);

OA21x2_ASAP7_75t_L g5666 ( 
.A1(n_4897),
.A2(n_3298),
.B(n_3295),
.Y(n_5666)
);

AND2x2_ASAP7_75t_L g5667 ( 
.A(n_4906),
.B(n_4284),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_4907),
.B(n_4296),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_5191),
.B(n_3302),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_4911),
.Y(n_5670)
);

AOI22xp5_ASAP7_75t_L g5671 ( 
.A1(n_4914),
.A2(n_2997),
.B1(n_2999),
.B2(n_2996),
.Y(n_5671)
);

BUFx6f_ASAP7_75t_L g5672 ( 
.A(n_4922),
.Y(n_5672)
);

BUFx6f_ASAP7_75t_L g5673 ( 
.A(n_4923),
.Y(n_5673)
);

INVx2_ASAP7_75t_L g5674 ( 
.A(n_4926),
.Y(n_5674)
);

BUFx6f_ASAP7_75t_L g5675 ( 
.A(n_4939),
.Y(n_5675)
);

AND2x4_ASAP7_75t_L g5676 ( 
.A(n_4946),
.B(n_3307),
.Y(n_5676)
);

INVx3_ASAP7_75t_L g5677 ( 
.A(n_4948),
.Y(n_5677)
);

BUFx12f_ASAP7_75t_L g5678 ( 
.A(n_4964),
.Y(n_5678)
);

INVx2_ASAP7_75t_L g5679 ( 
.A(n_4895),
.Y(n_5679)
);

INVx4_ASAP7_75t_L g5680 ( 
.A(n_4735),
.Y(n_5680)
);

AND2x4_ASAP7_75t_L g5681 ( 
.A(n_4901),
.B(n_3311),
.Y(n_5681)
);

OA21x2_ASAP7_75t_L g5682 ( 
.A1(n_4738),
.A2(n_3314),
.B(n_3312),
.Y(n_5682)
);

BUFx6f_ASAP7_75t_L g5683 ( 
.A(n_4965),
.Y(n_5683)
);

BUFx6f_ASAP7_75t_L g5684 ( 
.A(n_4967),
.Y(n_5684)
);

INVx3_ASAP7_75t_L g5685 ( 
.A(n_4968),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_4739),
.Y(n_5686)
);

INVx2_ASAP7_75t_L g5687 ( 
.A(n_4908),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_4744),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_4916),
.Y(n_5689)
);

INVx3_ASAP7_75t_L g5690 ( 
.A(n_4747),
.Y(n_5690)
);

NAND2xp5_ASAP7_75t_L g5691 ( 
.A(n_4751),
.B(n_4293),
.Y(n_5691)
);

CKINVDCx11_ASAP7_75t_R g5692 ( 
.A(n_4960),
.Y(n_5692)
);

OAI22xp5_ASAP7_75t_L g5693 ( 
.A1(n_4919),
.A2(n_3004),
.B1(n_3009),
.B2(n_3002),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_4758),
.Y(n_5694)
);

HB1xp67_ASAP7_75t_L g5695 ( 
.A(n_4756),
.Y(n_5695)
);

BUFx6f_ASAP7_75t_L g5696 ( 
.A(n_5171),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5173),
.Y(n_5697)
);

INVx2_ASAP7_75t_L g5698 ( 
.A(n_4927),
.Y(n_5698)
);

BUFx2_ASAP7_75t_L g5699 ( 
.A(n_4962),
.Y(n_5699)
);

BUFx6f_ASAP7_75t_L g5700 ( 
.A(n_5180),
.Y(n_5700)
);

INVx2_ASAP7_75t_L g5701 ( 
.A(n_4928),
.Y(n_5701)
);

HB1xp67_ASAP7_75t_L g5702 ( 
.A(n_4762),
.Y(n_5702)
);

HB1xp67_ASAP7_75t_L g5703 ( 
.A(n_4776),
.Y(n_5703)
);

AND2x4_ASAP7_75t_L g5704 ( 
.A(n_4933),
.B(n_3317),
.Y(n_5704)
);

HB1xp67_ASAP7_75t_L g5705 ( 
.A(n_4781),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_4934),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_4935),
.Y(n_5707)
);

INVx2_ASAP7_75t_L g5708 ( 
.A(n_4937),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5183),
.B(n_4303),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_4944),
.Y(n_5710)
);

CKINVDCx16_ASAP7_75t_R g5711 ( 
.A(n_4793),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5185),
.Y(n_5712)
);

BUFx6f_ASAP7_75t_L g5713 ( 
.A(n_5188),
.Y(n_5713)
);

BUFx6f_ASAP7_75t_L g5714 ( 
.A(n_5192),
.Y(n_5714)
);

OAI22xp5_ASAP7_75t_L g5715 ( 
.A1(n_4949),
.A2(n_3013),
.B1(n_3016),
.B2(n_3010),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5194),
.Y(n_5716)
);

HB1xp67_ASAP7_75t_L g5717 ( 
.A(n_4795),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5199),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5201),
.Y(n_5719)
);

INVx5_ASAP7_75t_L g5720 ( 
.A(n_5200),
.Y(n_5720)
);

CKINVDCx5p33_ASAP7_75t_R g5721 ( 
.A(n_5212),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5213),
.Y(n_5722)
);

NAND2xp5_ASAP7_75t_L g5723 ( 
.A(n_5214),
.B(n_3321),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5217),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_L g5725 ( 
.A(n_5222),
.B(n_3324),
.Y(n_5725)
);

INVx1_ASAP7_75t_SL g5726 ( 
.A(n_4796),
.Y(n_5726)
);

BUFx6f_ASAP7_75t_L g5727 ( 
.A(n_5232),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_5234),
.Y(n_5728)
);

BUFx6f_ASAP7_75t_L g5729 ( 
.A(n_4806),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_5230),
.Y(n_5730)
);

BUFx2_ASAP7_75t_L g5731 ( 
.A(n_4833),
.Y(n_5731)
);

NOR2x1_ASAP7_75t_L g5732 ( 
.A(n_4810),
.B(n_3326),
.Y(n_5732)
);

OAI21x1_ASAP7_75t_L g5733 ( 
.A1(n_4815),
.A2(n_3341),
.B(n_3338),
.Y(n_5733)
);

BUFx6f_ASAP7_75t_L g5734 ( 
.A(n_4818),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_4832),
.Y(n_5735)
);

INVx2_ASAP7_75t_L g5736 ( 
.A(n_5179),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5197),
.Y(n_5737)
);

BUFx2_ASAP7_75t_L g5738 ( 
.A(n_5202),
.Y(n_5738)
);

NAND2xp33_ASAP7_75t_L g5739 ( 
.A(n_5205),
.B(n_3017),
.Y(n_5739)
);

HB1xp67_ASAP7_75t_L g5740 ( 
.A(n_5211),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5215),
.Y(n_5741)
);

CKINVDCx11_ASAP7_75t_R g5742 ( 
.A(n_5216),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5225),
.Y(n_5743)
);

CKINVDCx5p33_ASAP7_75t_R g5744 ( 
.A(n_5227),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5058),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5058),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5058),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5058),
.Y(n_5748)
);

AND2x6_ASAP7_75t_L g5749 ( 
.A(n_4945),
.B(n_3345),
.Y(n_5749)
);

BUFx6f_ASAP7_75t_L g5750 ( 
.A(n_4784),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5098),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5058),
.Y(n_5752)
);

BUFx3_ASAP7_75t_L g5753 ( 
.A(n_4768),
.Y(n_5753)
);

OA21x2_ASAP7_75t_L g5754 ( 
.A1(n_5047),
.A2(n_3354),
.B(n_3347),
.Y(n_5754)
);

OAI22xp5_ASAP7_75t_SL g5755 ( 
.A1(n_5010),
.A2(n_3495),
.B1(n_3579),
.B2(n_3478),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5098),
.Y(n_5756)
);

AND2x6_ASAP7_75t_L g5757 ( 
.A(n_4945),
.B(n_3356),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_4768),
.Y(n_5758)
);

OAI22xp5_ASAP7_75t_SL g5759 ( 
.A1(n_5010),
.A2(n_3585),
.B1(n_3599),
.B2(n_3583),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5058),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5058),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5098),
.Y(n_5762)
);

AOI22xp5_ASAP7_75t_L g5763 ( 
.A1(n_5045),
.A2(n_3022),
.B1(n_3025),
.B2(n_3024),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5058),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5098),
.Y(n_5765)
);

OAI22xp5_ASAP7_75t_SL g5766 ( 
.A1(n_5010),
.A2(n_3626),
.B1(n_3628),
.B2(n_3624),
.Y(n_5766)
);

OAI21x1_ASAP7_75t_L g5767 ( 
.A1(n_4736),
.A2(n_3362),
.B(n_3360),
.Y(n_5767)
);

AND2x4_ASAP7_75t_L g5768 ( 
.A(n_4768),
.B(n_3364),
.Y(n_5768)
);

OAI22xp5_ASAP7_75t_L g5769 ( 
.A1(n_5082),
.A2(n_3026),
.B1(n_3031),
.B2(n_3028),
.Y(n_5769)
);

INVx5_ASAP7_75t_L g5770 ( 
.A(n_4847),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5058),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5058),
.Y(n_5772)
);

AND2x4_ASAP7_75t_L g5773 ( 
.A(n_4768),
.B(n_3367),
.Y(n_5773)
);

OAI22xp5_ASAP7_75t_SL g5774 ( 
.A1(n_5010),
.A2(n_3636),
.B1(n_3666),
.B2(n_3633),
.Y(n_5774)
);

INVx2_ASAP7_75t_L g5775 ( 
.A(n_5098),
.Y(n_5775)
);

INVx2_ASAP7_75t_SL g5776 ( 
.A(n_4972),
.Y(n_5776)
);

AND2x2_ASAP7_75t_L g5777 ( 
.A(n_5093),
.B(n_4296),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5058),
.Y(n_5778)
);

CKINVDCx11_ASAP7_75t_R g5779 ( 
.A(n_4861),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5098),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5098),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5098),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5093),
.B(n_4299),
.Y(n_5783)
);

NAND2xp5_ASAP7_75t_L g5784 ( 
.A(n_5047),
.B(n_3371),
.Y(n_5784)
);

BUFx2_ASAP7_75t_L g5785 ( 
.A(n_4972),
.Y(n_5785)
);

BUFx2_ASAP7_75t_L g5786 ( 
.A(n_4972),
.Y(n_5786)
);

AND2x4_ASAP7_75t_L g5787 ( 
.A(n_4768),
.B(n_3375),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5098),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5058),
.Y(n_5789)
);

BUFx3_ASAP7_75t_L g5790 ( 
.A(n_4768),
.Y(n_5790)
);

AND2x4_ASAP7_75t_L g5791 ( 
.A(n_4768),
.B(n_3376),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5098),
.Y(n_5792)
);

AND2x2_ASAP7_75t_L g5793 ( 
.A(n_5093),
.B(n_3034),
.Y(n_5793)
);

AND2x2_ASAP7_75t_L g5794 ( 
.A(n_5093),
.B(n_3036),
.Y(n_5794)
);

NOR2xp33_ASAP7_75t_L g5795 ( 
.A(n_5093),
.B(n_3037),
.Y(n_5795)
);

AND2x2_ASAP7_75t_L g5796 ( 
.A(n_5093),
.B(n_3040),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5098),
.Y(n_5797)
);

NOR2xp33_ASAP7_75t_R g5798 ( 
.A(n_4829),
.B(n_3670),
.Y(n_5798)
);

INVx2_ASAP7_75t_L g5799 ( 
.A(n_5098),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5058),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5098),
.Y(n_5801)
);

INVx3_ASAP7_75t_L g5802 ( 
.A(n_4784),
.Y(n_5802)
);

INVx3_ASAP7_75t_L g5803 ( 
.A(n_4784),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5058),
.Y(n_5804)
);

NAND2xp33_ASAP7_75t_L g5805 ( 
.A(n_5047),
.B(n_3041),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_5058),
.Y(n_5806)
);

AND2x4_ASAP7_75t_L g5807 ( 
.A(n_4768),
.B(n_3378),
.Y(n_5807)
);

AND2x2_ASAP7_75t_L g5808 ( 
.A(n_5093),
.B(n_3043),
.Y(n_5808)
);

BUFx6f_ASAP7_75t_L g5809 ( 
.A(n_4784),
.Y(n_5809)
);

NAND2xp33_ASAP7_75t_L g5810 ( 
.A(n_5047),
.B(n_3047),
.Y(n_5810)
);

INVx2_ASAP7_75t_L g5811 ( 
.A(n_5098),
.Y(n_5811)
);

AND2x4_ASAP7_75t_L g5812 ( 
.A(n_4768),
.B(n_3386),
.Y(n_5812)
);

CKINVDCx5p33_ASAP7_75t_R g5813 ( 
.A(n_4763),
.Y(n_5813)
);

HB1xp67_ASAP7_75t_L g5814 ( 
.A(n_5314),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5777),
.Y(n_5815)
);

CKINVDCx5p33_ASAP7_75t_R g5816 ( 
.A(n_5246),
.Y(n_5816)
);

CKINVDCx5p33_ASAP7_75t_R g5817 ( 
.A(n_5813),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_5257),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_5274),
.Y(n_5819)
);

CKINVDCx5p33_ASAP7_75t_R g5820 ( 
.A(n_5288),
.Y(n_5820)
);

CKINVDCx5p33_ASAP7_75t_R g5821 ( 
.A(n_5329),
.Y(n_5821)
);

CKINVDCx5p33_ASAP7_75t_R g5822 ( 
.A(n_5392),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5269),
.Y(n_5823)
);

CKINVDCx5p33_ASAP7_75t_R g5824 ( 
.A(n_5403),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5776),
.B(n_3695),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_5272),
.Y(n_5826)
);

CKINVDCx20_ASAP7_75t_R g5827 ( 
.A(n_5381),
.Y(n_5827)
);

CKINVDCx20_ASAP7_75t_R g5828 ( 
.A(n_5742),
.Y(n_5828)
);

INVx2_ASAP7_75t_L g5829 ( 
.A(n_5299),
.Y(n_5829)
);

CKINVDCx20_ASAP7_75t_R g5830 ( 
.A(n_5711),
.Y(n_5830)
);

NOR2xp33_ASAP7_75t_R g5831 ( 
.A(n_5478),
.B(n_3701),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5271),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5280),
.Y(n_5833)
);

BUFx6f_ASAP7_75t_L g5834 ( 
.A(n_5263),
.Y(n_5834)
);

BUFx3_ASAP7_75t_L g5835 ( 
.A(n_5753),
.Y(n_5835)
);

BUFx2_ASAP7_75t_L g5836 ( 
.A(n_5319),
.Y(n_5836)
);

CKINVDCx5p33_ASAP7_75t_R g5837 ( 
.A(n_5526),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_5604),
.Y(n_5838)
);

HB1xp67_ASAP7_75t_L g5839 ( 
.A(n_5783),
.Y(n_5839)
);

CKINVDCx20_ASAP7_75t_R g5840 ( 
.A(n_5692),
.Y(n_5840)
);

CKINVDCx5p33_ASAP7_75t_R g5841 ( 
.A(n_5606),
.Y(n_5841)
);

CKINVDCx5p33_ASAP7_75t_R g5842 ( 
.A(n_5616),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5273),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5275),
.Y(n_5844)
);

CKINVDCx5p33_ASAP7_75t_R g5845 ( 
.A(n_5721),
.Y(n_5845)
);

CKINVDCx20_ASAP7_75t_R g5846 ( 
.A(n_5744),
.Y(n_5846)
);

CKINVDCx5p33_ASAP7_75t_R g5847 ( 
.A(n_5365),
.Y(n_5847)
);

CKINVDCx20_ASAP7_75t_R g5848 ( 
.A(n_5258),
.Y(n_5848)
);

CKINVDCx5p33_ASAP7_75t_R g5849 ( 
.A(n_5635),
.Y(n_5849)
);

CKINVDCx5p33_ASAP7_75t_R g5850 ( 
.A(n_5650),
.Y(n_5850)
);

CKINVDCx20_ASAP7_75t_R g5851 ( 
.A(n_5779),
.Y(n_5851)
);

AND2x2_ASAP7_75t_L g5852 ( 
.A(n_5308),
.B(n_3728),
.Y(n_5852)
);

CKINVDCx5p33_ASAP7_75t_R g5853 ( 
.A(n_5659),
.Y(n_5853)
);

AND3x2_ASAP7_75t_L g5854 ( 
.A(n_5785),
.B(n_3395),
.C(n_3387),
.Y(n_5854)
);

INVxp67_ASAP7_75t_L g5855 ( 
.A(n_5795),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5276),
.Y(n_5856)
);

CKINVDCx5p33_ASAP7_75t_R g5857 ( 
.A(n_5672),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_5673),
.Y(n_5858)
);

CKINVDCx5p33_ASAP7_75t_R g5859 ( 
.A(n_5675),
.Y(n_5859)
);

NOR2xp33_ASAP7_75t_R g5860 ( 
.A(n_5685),
.B(n_3764),
.Y(n_5860)
);

CKINVDCx20_ASAP7_75t_R g5861 ( 
.A(n_5546),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_5514),
.Y(n_5862)
);

CKINVDCx5p33_ASAP7_75t_R g5863 ( 
.A(n_5798),
.Y(n_5863)
);

INVx2_ASAP7_75t_L g5864 ( 
.A(n_5282),
.Y(n_5864)
);

CKINVDCx20_ASAP7_75t_R g5865 ( 
.A(n_5786),
.Y(n_5865)
);

BUFx3_ASAP7_75t_L g5866 ( 
.A(n_5758),
.Y(n_5866)
);

HB1xp67_ASAP7_75t_L g5867 ( 
.A(n_5344),
.Y(n_5867)
);

NOR2xp33_ASAP7_75t_R g5868 ( 
.A(n_5690),
.B(n_3790),
.Y(n_5868)
);

AND2x2_ASAP7_75t_L g5869 ( 
.A(n_5247),
.B(n_3793),
.Y(n_5869)
);

CKINVDCx5p33_ASAP7_75t_R g5870 ( 
.A(n_5696),
.Y(n_5870)
);

CKINVDCx5p33_ASAP7_75t_R g5871 ( 
.A(n_5700),
.Y(n_5871)
);

BUFx2_ASAP7_75t_L g5872 ( 
.A(n_5419),
.Y(n_5872)
);

CKINVDCx5p33_ASAP7_75t_R g5873 ( 
.A(n_5713),
.Y(n_5873)
);

CKINVDCx5p33_ASAP7_75t_R g5874 ( 
.A(n_5714),
.Y(n_5874)
);

NOR2xp33_ASAP7_75t_L g5875 ( 
.A(n_5239),
.B(n_3053),
.Y(n_5875)
);

CKINVDCx20_ASAP7_75t_R g5876 ( 
.A(n_5738),
.Y(n_5876)
);

CKINVDCx20_ASAP7_75t_R g5877 ( 
.A(n_5550),
.Y(n_5877)
);

NOR2xp33_ASAP7_75t_R g5878 ( 
.A(n_5664),
.B(n_5677),
.Y(n_5878)
);

BUFx6f_ASAP7_75t_L g5879 ( 
.A(n_5268),
.Y(n_5879)
);

INVx2_ASAP7_75t_L g5880 ( 
.A(n_5285),
.Y(n_5880)
);

CKINVDCx5p33_ASAP7_75t_R g5881 ( 
.A(n_5727),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5278),
.Y(n_5882)
);

NOR2xp33_ASAP7_75t_R g5883 ( 
.A(n_5267),
.B(n_3813),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5281),
.Y(n_5884)
);

CKINVDCx5p33_ASAP7_75t_R g5885 ( 
.A(n_5493),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5286),
.Y(n_5886)
);

CKINVDCx20_ASAP7_75t_R g5887 ( 
.A(n_5632),
.Y(n_5887)
);

CKINVDCx5p33_ASAP7_75t_R g5888 ( 
.A(n_5678),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5291),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_5284),
.Y(n_5890)
);

CKINVDCx5p33_ASAP7_75t_R g5891 ( 
.A(n_5729),
.Y(n_5891)
);

CKINVDCx20_ASAP7_75t_R g5892 ( 
.A(n_5731),
.Y(n_5892)
);

CKINVDCx20_ASAP7_75t_R g5893 ( 
.A(n_5377),
.Y(n_5893)
);

CKINVDCx5p33_ASAP7_75t_R g5894 ( 
.A(n_5734),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5296),
.Y(n_5895)
);

CKINVDCx5p33_ASAP7_75t_R g5896 ( 
.A(n_5680),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5290),
.Y(n_5897)
);

NOR2xp33_ASAP7_75t_L g5898 ( 
.A(n_5642),
.B(n_3056),
.Y(n_5898)
);

CKINVDCx5p33_ASAP7_75t_R g5899 ( 
.A(n_5553),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5293),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5301),
.Y(n_5901)
);

HB1xp67_ASAP7_75t_L g5902 ( 
.A(n_5298),
.Y(n_5902)
);

INVx3_ASAP7_75t_L g5903 ( 
.A(n_5242),
.Y(n_5903)
);

BUFx2_ASAP7_75t_L g5904 ( 
.A(n_5494),
.Y(n_5904)
);

CKINVDCx20_ASAP7_75t_R g5905 ( 
.A(n_5770),
.Y(n_5905)
);

BUFx2_ASAP7_75t_L g5906 ( 
.A(n_5494),
.Y(n_5906)
);

CKINVDCx5p33_ASAP7_75t_R g5907 ( 
.A(n_5256),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5297),
.Y(n_5908)
);

CKINVDCx5p33_ASAP7_75t_R g5909 ( 
.A(n_5658),
.Y(n_5909)
);

CKINVDCx20_ASAP7_75t_R g5910 ( 
.A(n_5695),
.Y(n_5910)
);

INVx3_ASAP7_75t_L g5911 ( 
.A(n_5248),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_5305),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_L g5913 ( 
.A(n_5320),
.B(n_3059),
.Y(n_5913)
);

CKINVDCx20_ASAP7_75t_R g5914 ( 
.A(n_5702),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5302),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5304),
.Y(n_5916)
);

CKINVDCx5p33_ASAP7_75t_R g5917 ( 
.A(n_5594),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5309),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5311),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5328),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5572),
.B(n_3814),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_5726),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5330),
.Y(n_5923)
);

BUFx3_ASAP7_75t_L g5924 ( 
.A(n_5790),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_SL g5925 ( 
.A(n_5599),
.B(n_3061),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5331),
.Y(n_5926)
);

INVx2_ASAP7_75t_SL g5927 ( 
.A(n_5378),
.Y(n_5927)
);

CKINVDCx5p33_ASAP7_75t_R g5928 ( 
.A(n_5720),
.Y(n_5928)
);

CKINVDCx5p33_ASAP7_75t_R g5929 ( 
.A(n_5587),
.Y(n_5929)
);

NOR2xp33_ASAP7_75t_R g5930 ( 
.A(n_5382),
.B(n_3857),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5332),
.Y(n_5931)
);

CKINVDCx5p33_ASAP7_75t_R g5932 ( 
.A(n_5683),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5337),
.Y(n_5933)
);

CKINVDCx5p33_ASAP7_75t_R g5934 ( 
.A(n_5684),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_5592),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5307),
.Y(n_5936)
);

CKINVDCx5p33_ASAP7_75t_R g5937 ( 
.A(n_5602),
.Y(n_5937)
);

CKINVDCx5p33_ASAP7_75t_R g5938 ( 
.A(n_5703),
.Y(n_5938)
);

CKINVDCx5p33_ASAP7_75t_R g5939 ( 
.A(n_5705),
.Y(n_5939)
);

CKINVDCx5p33_ASAP7_75t_R g5940 ( 
.A(n_5717),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5339),
.Y(n_5941)
);

CKINVDCx20_ASAP7_75t_R g5942 ( 
.A(n_5740),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5318),
.Y(n_5943)
);

BUFx2_ASAP7_75t_L g5944 ( 
.A(n_5527),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_5452),
.B(n_3062),
.Y(n_5945)
);

AND2x4_ASAP7_75t_L g5946 ( 
.A(n_5254),
.B(n_5310),
.Y(n_5946)
);

AO21x2_ASAP7_75t_L g5947 ( 
.A1(n_5655),
.A2(n_3397),
.B(n_3396),
.Y(n_5947)
);

CKINVDCx5p33_ASAP7_75t_R g5948 ( 
.A(n_5538),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_5520),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_5661),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5341),
.Y(n_5951)
);

CKINVDCx5p33_ASAP7_75t_R g5952 ( 
.A(n_5674),
.Y(n_5952)
);

CKINVDCx5p33_ASAP7_75t_R g5953 ( 
.A(n_5362),
.Y(n_5953)
);

NAND2xp33_ASAP7_75t_R g5954 ( 
.A(n_5681),
.B(n_3064),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_5699),
.Y(n_5955)
);

OR2x2_ASAP7_75t_L g5956 ( 
.A(n_5294),
.B(n_3065),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5345),
.Y(n_5957)
);

CKINVDCx5p33_ASAP7_75t_R g5958 ( 
.A(n_5716),
.Y(n_5958)
);

BUFx3_ASAP7_75t_L g5959 ( 
.A(n_5361),
.Y(n_5959)
);

BUFx6f_ASAP7_75t_L g5960 ( 
.A(n_5277),
.Y(n_5960)
);

XOR2xp5_ASAP7_75t_L g5961 ( 
.A(n_5265),
.B(n_3880),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5349),
.Y(n_5962)
);

INVxp67_ASAP7_75t_SL g5963 ( 
.A(n_5436),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5358),
.B(n_3910),
.Y(n_5964)
);

HB1xp67_ASAP7_75t_L g5965 ( 
.A(n_5754),
.Y(n_5965)
);

CKINVDCx5p33_ASAP7_75t_R g5966 ( 
.A(n_5718),
.Y(n_5966)
);

CKINVDCx20_ASAP7_75t_R g5967 ( 
.A(n_5497),
.Y(n_5967)
);

CKINVDCx5p33_ASAP7_75t_R g5968 ( 
.A(n_5728),
.Y(n_5968)
);

CKINVDCx5p33_ASAP7_75t_R g5969 ( 
.A(n_5524),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5357),
.Y(n_5970)
);

CKINVDCx5p33_ASAP7_75t_R g5971 ( 
.A(n_5544),
.Y(n_5971)
);

AND3x2_ASAP7_75t_L g5972 ( 
.A(n_5355),
.B(n_3410),
.C(n_3401),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5459),
.B(n_5460),
.Y(n_5973)
);

CKINVDCx5p33_ASAP7_75t_R g5974 ( 
.A(n_5670),
.Y(n_5974)
);

BUFx2_ASAP7_75t_L g5975 ( 
.A(n_5527),
.Y(n_5975)
);

CKINVDCx20_ASAP7_75t_R g5976 ( 
.A(n_5360),
.Y(n_5976)
);

CKINVDCx5p33_ASAP7_75t_R g5977 ( 
.A(n_5369),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5364),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5335),
.Y(n_5979)
);

INVx8_ASAP7_75t_L g5980 ( 
.A(n_5749),
.Y(n_5980)
);

CKINVDCx5p33_ASAP7_75t_R g5981 ( 
.A(n_5388),
.Y(n_5981)
);

CKINVDCx20_ASAP7_75t_R g5982 ( 
.A(n_5563),
.Y(n_5982)
);

BUFx6f_ASAP7_75t_L g5983 ( 
.A(n_5240),
.Y(n_5983)
);

NOR2xp33_ASAP7_75t_R g5984 ( 
.A(n_5805),
.B(n_3918),
.Y(n_5984)
);

CKINVDCx5p33_ASAP7_75t_R g5985 ( 
.A(n_5429),
.Y(n_5985)
);

CKINVDCx5p33_ASAP7_75t_R g5986 ( 
.A(n_5475),
.Y(n_5986)
);

CKINVDCx5p33_ASAP7_75t_R g5987 ( 
.A(n_5495),
.Y(n_5987)
);

CKINVDCx5p33_ASAP7_75t_R g5988 ( 
.A(n_5508),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5374),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5379),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_5686),
.Y(n_5991)
);

CKINVDCx5p33_ASAP7_75t_R g5992 ( 
.A(n_5688),
.Y(n_5992)
);

CKINVDCx5p33_ASAP7_75t_R g5993 ( 
.A(n_5694),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5384),
.Y(n_5994)
);

CKINVDCx20_ASAP7_75t_R g5995 ( 
.A(n_5414),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5397),
.Y(n_5996)
);

CKINVDCx5p33_ASAP7_75t_R g5997 ( 
.A(n_5697),
.Y(n_5997)
);

CKINVDCx5p33_ASAP7_75t_R g5998 ( 
.A(n_5712),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5338),
.Y(n_5999)
);

INVx2_ASAP7_75t_L g6000 ( 
.A(n_5350),
.Y(n_6000)
);

CKINVDCx5p33_ASAP7_75t_R g6001 ( 
.A(n_5719),
.Y(n_6001)
);

CKINVDCx5p33_ASAP7_75t_R g6002 ( 
.A(n_5722),
.Y(n_6002)
);

BUFx6f_ASAP7_75t_L g6003 ( 
.A(n_5244),
.Y(n_6003)
);

HB1xp67_ASAP7_75t_L g6004 ( 
.A(n_5793),
.Y(n_6004)
);

CKINVDCx5p33_ASAP7_75t_R g6005 ( 
.A(n_5724),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5402),
.Y(n_6006)
);

NOR2xp33_ASAP7_75t_R g6007 ( 
.A(n_5810),
.B(n_3931),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5409),
.Y(n_6008)
);

CKINVDCx5p33_ASAP7_75t_R g6009 ( 
.A(n_5540),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5411),
.Y(n_6010)
);

CKINVDCx5p33_ASAP7_75t_R g6011 ( 
.A(n_5518),
.Y(n_6011)
);

CKINVDCx5p33_ASAP7_75t_R g6012 ( 
.A(n_5564),
.Y(n_6012)
);

CKINVDCx5p33_ASAP7_75t_R g6013 ( 
.A(n_5325),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5351),
.Y(n_6014)
);

INVx2_ASAP7_75t_L g6015 ( 
.A(n_5354),
.Y(n_6015)
);

CKINVDCx5p33_ASAP7_75t_R g6016 ( 
.A(n_5445),
.Y(n_6016)
);

INVx2_ASAP7_75t_L g6017 ( 
.A(n_5375),
.Y(n_6017)
);

CKINVDCx20_ASAP7_75t_R g6018 ( 
.A(n_5646),
.Y(n_6018)
);

CKINVDCx5p33_ASAP7_75t_R g6019 ( 
.A(n_5735),
.Y(n_6019)
);

HB1xp67_ASAP7_75t_L g6020 ( 
.A(n_5794),
.Y(n_6020)
);

NOR2xp33_ASAP7_75t_R g6021 ( 
.A(n_5739),
.B(n_3956),
.Y(n_6021)
);

NOR2xp33_ASAP7_75t_R g6022 ( 
.A(n_5613),
.B(n_5730),
.Y(n_6022)
);

CKINVDCx5p33_ASAP7_75t_R g6023 ( 
.A(n_5736),
.Y(n_6023)
);

CKINVDCx5p33_ASAP7_75t_R g6024 ( 
.A(n_5428),
.Y(n_6024)
);

CKINVDCx6p67_ASAP7_75t_R g6025 ( 
.A(n_5644),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_L g6026 ( 
.A(n_5466),
.B(n_3066),
.Y(n_6026)
);

INVx2_ASAP7_75t_L g6027 ( 
.A(n_5389),
.Y(n_6027)
);

CKINVDCx20_ASAP7_75t_R g6028 ( 
.A(n_5648),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5415),
.Y(n_6029)
);

BUFx6f_ASAP7_75t_L g6030 ( 
.A(n_5253),
.Y(n_6030)
);

CKINVDCx5p33_ASAP7_75t_R g6031 ( 
.A(n_5679),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5416),
.Y(n_6032)
);

INVx3_ASAP7_75t_L g6033 ( 
.A(n_5252),
.Y(n_6033)
);

CKINVDCx5p33_ASAP7_75t_R g6034 ( 
.A(n_5687),
.Y(n_6034)
);

NOR2xp67_ASAP7_75t_L g6035 ( 
.A(n_5370),
.B(n_3067),
.Y(n_6035)
);

CKINVDCx20_ASAP7_75t_R g6036 ( 
.A(n_5522),
.Y(n_6036)
);

AND2x2_ASAP7_75t_L g6037 ( 
.A(n_5796),
.B(n_3973),
.Y(n_6037)
);

CKINVDCx5p33_ASAP7_75t_R g6038 ( 
.A(n_5689),
.Y(n_6038)
);

CKINVDCx20_ASAP7_75t_R g6039 ( 
.A(n_5427),
.Y(n_6039)
);

NOR2xp33_ASAP7_75t_R g6040 ( 
.A(n_5737),
.B(n_3980),
.Y(n_6040)
);

CKINVDCx5p33_ASAP7_75t_R g6041 ( 
.A(n_5698),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5417),
.Y(n_6042)
);

AOI22xp5_ASAP7_75t_L g6043 ( 
.A1(n_5333),
.A2(n_3988),
.B1(n_4005),
.B2(n_3985),
.Y(n_6043)
);

HB1xp67_ASAP7_75t_L g6044 ( 
.A(n_5808),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5418),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_5511),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5515),
.Y(n_6047)
);

CKINVDCx5p33_ASAP7_75t_R g6048 ( 
.A(n_5701),
.Y(n_6048)
);

NAND2xp33_ASAP7_75t_R g6049 ( 
.A(n_5704),
.B(n_3068),
.Y(n_6049)
);

NOR2xp33_ASAP7_75t_L g6050 ( 
.A(n_5654),
.B(n_3069),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5531),
.Y(n_6051)
);

INVxp67_ASAP7_75t_L g6052 ( 
.A(n_5236),
.Y(n_6052)
);

CKINVDCx5p33_ASAP7_75t_R g6053 ( 
.A(n_5706),
.Y(n_6053)
);

CKINVDCx5p33_ASAP7_75t_R g6054 ( 
.A(n_5707),
.Y(n_6054)
);

CKINVDCx5p33_ASAP7_75t_R g6055 ( 
.A(n_5708),
.Y(n_6055)
);

CKINVDCx5p33_ASAP7_75t_R g6056 ( 
.A(n_5710),
.Y(n_6056)
);

INVx1_ASAP7_75t_SL g6057 ( 
.A(n_5408),
.Y(n_6057)
);

NOR2xp33_ASAP7_75t_R g6058 ( 
.A(n_5741),
.B(n_4065),
.Y(n_6058)
);

CKINVDCx20_ASAP7_75t_R g6059 ( 
.A(n_5467),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5532),
.Y(n_6060)
);

CKINVDCx5p33_ASAP7_75t_R g6061 ( 
.A(n_5743),
.Y(n_6061)
);

CKINVDCx20_ASAP7_75t_R g6062 ( 
.A(n_5468),
.Y(n_6062)
);

NOR2xp33_ASAP7_75t_R g6063 ( 
.A(n_5660),
.B(n_4068),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_5630),
.Y(n_6064)
);

CKINVDCx5p33_ASAP7_75t_R g6065 ( 
.A(n_5608),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5394),
.Y(n_6066)
);

INVx3_ASAP7_75t_L g6067 ( 
.A(n_5751),
.Y(n_6067)
);

BUFx6f_ASAP7_75t_L g6068 ( 
.A(n_5260),
.Y(n_6068)
);

INVx2_ASAP7_75t_L g6069 ( 
.A(n_5398),
.Y(n_6069)
);

INVx1_ASAP7_75t_SL g6070 ( 
.A(n_5255),
.Y(n_6070)
);

CKINVDCx5p33_ASAP7_75t_R g6071 ( 
.A(n_5368),
.Y(n_6071)
);

NOR2xp67_ASAP7_75t_L g6072 ( 
.A(n_5513),
.B(n_3071),
.Y(n_6072)
);

INVx3_ASAP7_75t_L g6073 ( 
.A(n_5756),
.Y(n_6073)
);

CKINVDCx5p33_ASAP7_75t_R g6074 ( 
.A(n_5368),
.Y(n_6074)
);

INVx2_ASAP7_75t_L g6075 ( 
.A(n_5420),
.Y(n_6075)
);

INVx2_ASAP7_75t_L g6076 ( 
.A(n_5426),
.Y(n_6076)
);

INVxp67_ASAP7_75t_L g6077 ( 
.A(n_5322),
.Y(n_6077)
);

INVx3_ASAP7_75t_L g6078 ( 
.A(n_5762),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_5432),
.Y(n_6079)
);

CKINVDCx5p33_ASAP7_75t_R g6080 ( 
.A(n_5413),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5533),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5543),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5551),
.Y(n_6083)
);

CKINVDCx5p33_ASAP7_75t_R g6084 ( 
.A(n_5413),
.Y(n_6084)
);

CKINVDCx5p33_ASAP7_75t_R g6085 ( 
.A(n_5619),
.Y(n_6085)
);

INVx2_ASAP7_75t_L g6086 ( 
.A(n_5433),
.Y(n_6086)
);

CKINVDCx5p33_ASAP7_75t_R g6087 ( 
.A(n_5644),
.Y(n_6087)
);

BUFx10_ASAP7_75t_L g6088 ( 
.A(n_5676),
.Y(n_6088)
);

CKINVDCx5p33_ASAP7_75t_R g6089 ( 
.A(n_5598),
.Y(n_6089)
);

INVx3_ASAP7_75t_L g6090 ( 
.A(n_5765),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_5454),
.Y(n_6091)
);

INVx2_ASAP7_75t_L g6092 ( 
.A(n_5455),
.Y(n_6092)
);

INVxp67_ASAP7_75t_SL g6093 ( 
.A(n_5306),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5556),
.Y(n_6094)
);

NOR2xp33_ASAP7_75t_R g6095 ( 
.A(n_5662),
.B(n_4070),
.Y(n_6095)
);

CKINVDCx5p33_ASAP7_75t_R g6096 ( 
.A(n_5600),
.Y(n_6096)
);

CKINVDCx5p33_ASAP7_75t_R g6097 ( 
.A(n_5324),
.Y(n_6097)
);

CKINVDCx5p33_ASAP7_75t_R g6098 ( 
.A(n_5324),
.Y(n_6098)
);

CKINVDCx5p33_ASAP7_75t_R g6099 ( 
.A(n_5693),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5557),
.Y(n_6100)
);

CKINVDCx20_ASAP7_75t_R g6101 ( 
.A(n_5491),
.Y(n_6101)
);

NOR2xp33_ASAP7_75t_L g6102 ( 
.A(n_5723),
.B(n_3073),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_5558),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5559),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_5715),
.Y(n_6105)
);

HB1xp67_ASAP7_75t_L g6106 ( 
.A(n_5631),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_5560),
.Y(n_6107)
);

CKINVDCx5p33_ASAP7_75t_R g6108 ( 
.A(n_5638),
.Y(n_6108)
);

NAND2xp5_ASAP7_75t_SL g6109 ( 
.A(n_5390),
.B(n_3076),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_5562),
.Y(n_6110)
);

BUFx6f_ASAP7_75t_L g6111 ( 
.A(n_5750),
.Y(n_6111)
);

INVx2_ASAP7_75t_L g6112 ( 
.A(n_5457),
.Y(n_6112)
);

BUFx6f_ASAP7_75t_L g6113 ( 
.A(n_5809),
.Y(n_6113)
);

CKINVDCx20_ASAP7_75t_R g6114 ( 
.A(n_5755),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_5638),
.Y(n_6115)
);

OR2x2_ASAP7_75t_L g6116 ( 
.A(n_5342),
.B(n_3077),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5568),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_5504),
.Y(n_6118)
);

CKINVDCx5p33_ASAP7_75t_R g6119 ( 
.A(n_5614),
.Y(n_6119)
);

CKINVDCx5p33_ASAP7_75t_R g6120 ( 
.A(n_5407),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5473),
.Y(n_6121)
);

BUFx10_ASAP7_75t_L g6122 ( 
.A(n_5656),
.Y(n_6122)
);

CKINVDCx20_ASAP7_75t_R g6123 ( 
.A(n_5759),
.Y(n_6123)
);

CKINVDCx20_ASAP7_75t_R g6124 ( 
.A(n_5766),
.Y(n_6124)
);

CKINVDCx20_ASAP7_75t_R g6125 ( 
.A(n_5774),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5580),
.Y(n_6126)
);

NOR2xp33_ASAP7_75t_L g6127 ( 
.A(n_5725),
.B(n_3078),
.Y(n_6127)
);

CKINVDCx5p33_ASAP7_75t_R g6128 ( 
.A(n_5489),
.Y(n_6128)
);

CKINVDCx5p33_ASAP7_75t_R g6129 ( 
.A(n_5525),
.Y(n_6129)
);

CKINVDCx5p33_ASAP7_75t_R g6130 ( 
.A(n_5333),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5584),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_5480),
.Y(n_6132)
);

NOR2xp33_ASAP7_75t_R g6133 ( 
.A(n_5665),
.B(n_4088),
.Y(n_6133)
);

NOR2xp33_ASAP7_75t_R g6134 ( 
.A(n_5651),
.B(n_4116),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_5438),
.Y(n_6135)
);

BUFx10_ASAP7_75t_L g6136 ( 
.A(n_5669),
.Y(n_6136)
);

CKINVDCx5p33_ASAP7_75t_R g6137 ( 
.A(n_5481),
.Y(n_6137)
);

NOR2xp33_ASAP7_75t_R g6138 ( 
.A(n_5652),
.B(n_4130),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_SL g6139 ( 
.A(n_5313),
.B(n_3079),
.Y(n_6139)
);

NOR2xp33_ASAP7_75t_R g6140 ( 
.A(n_5653),
.B(n_4144),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5590),
.Y(n_6141)
);

CKINVDCx20_ASAP7_75t_R g6142 ( 
.A(n_5439),
.Y(n_6142)
);

CKINVDCx20_ASAP7_75t_R g6143 ( 
.A(n_5259),
.Y(n_6143)
);

NAND2xp5_ASAP7_75t_SL g6144 ( 
.A(n_5326),
.B(n_3081),
.Y(n_6144)
);

AND2x2_ASAP7_75t_L g6145 ( 
.A(n_5476),
.B(n_4154),
.Y(n_6145)
);

CKINVDCx5p33_ASAP7_75t_R g6146 ( 
.A(n_5492),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_5486),
.Y(n_6147)
);

NAND2xp5_ASAP7_75t_L g6148 ( 
.A(n_5431),
.B(n_3085),
.Y(n_6148)
);

HB1xp67_ASAP7_75t_L g6149 ( 
.A(n_5334),
.Y(n_6149)
);

INVx1_ASAP7_75t_SL g6150 ( 
.A(n_5542),
.Y(n_6150)
);

BUFx10_ASAP7_75t_L g6151 ( 
.A(n_5634),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5596),
.Y(n_6152)
);

NOR2xp33_ASAP7_75t_R g6153 ( 
.A(n_5621),
.B(n_4166),
.Y(n_6153)
);

CKINVDCx5p33_ASAP7_75t_R g6154 ( 
.A(n_5501),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_5510),
.Y(n_6155)
);

CKINVDCx5p33_ASAP7_75t_R g6156 ( 
.A(n_5691),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_5512),
.Y(n_6157)
);

CKINVDCx5p33_ASAP7_75t_R g6158 ( 
.A(n_5709),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_5597),
.Y(n_6159)
);

AND3x2_ASAP7_75t_L g6160 ( 
.A(n_5405),
.B(n_3422),
.C(n_3421),
.Y(n_6160)
);

CKINVDCx20_ASAP7_75t_R g6161 ( 
.A(n_5353),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5443),
.Y(n_6162)
);

NOR2xp33_ASAP7_75t_SL g6163 ( 
.A(n_5657),
.B(n_4167),
.Y(n_6163)
);

CKINVDCx20_ASAP7_75t_R g6164 ( 
.A(n_5371),
.Y(n_6164)
);

OAI22xp5_ASAP7_75t_L g6165 ( 
.A1(n_5262),
.A2(n_3087),
.B1(n_3092),
.B2(n_3088),
.Y(n_6165)
);

OR2x2_ASAP7_75t_L g6166 ( 
.A(n_5620),
.B(n_3095),
.Y(n_6166)
);

CKINVDCx5p33_ASAP7_75t_R g6167 ( 
.A(n_5671),
.Y(n_6167)
);

CKINVDCx5p33_ASAP7_75t_R g6168 ( 
.A(n_5643),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_5561),
.Y(n_6169)
);

BUFx2_ASAP7_75t_L g6170 ( 
.A(n_5629),
.Y(n_6170)
);

BUFx3_ASAP7_75t_L g6171 ( 
.A(n_5317),
.Y(n_6171)
);

CKINVDCx5p33_ASAP7_75t_R g6172 ( 
.A(n_5663),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5461),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_5506),
.B(n_4175),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5472),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5516),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5474),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5487),
.Y(n_6178)
);

CKINVDCx20_ASAP7_75t_R g6179 ( 
.A(n_5238),
.Y(n_6179)
);

CKINVDCx5p33_ASAP7_75t_R g6180 ( 
.A(n_5667),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_5488),
.Y(n_6181)
);

CKINVDCx5p33_ASAP7_75t_R g6182 ( 
.A(n_5668),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5490),
.Y(n_6183)
);

NOR2xp33_ASAP7_75t_SL g6184 ( 
.A(n_5264),
.B(n_4183),
.Y(n_6184)
);

CKINVDCx20_ASAP7_75t_R g6185 ( 
.A(n_5633),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5496),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5499),
.Y(n_6187)
);

NOR2xp67_ASAP7_75t_L g6188 ( 
.A(n_5763),
.B(n_3099),
.Y(n_6188)
);

INVxp67_ASAP7_75t_L g6189 ( 
.A(n_5548),
.Y(n_6189)
);

CKINVDCx5p33_ASAP7_75t_R g6190 ( 
.A(n_5396),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5503),
.Y(n_6191)
);

CKINVDCx5p33_ASAP7_75t_R g6192 ( 
.A(n_5595),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_5340),
.B(n_4186),
.Y(n_6193)
);

CKINVDCx5p33_ASAP7_75t_R g6194 ( 
.A(n_5601),
.Y(n_6194)
);

CKINVDCx5p33_ASAP7_75t_R g6195 ( 
.A(n_5749),
.Y(n_6195)
);

INVx8_ASAP7_75t_L g6196 ( 
.A(n_5757),
.Y(n_6196)
);

CKINVDCx8_ASAP7_75t_R g6197 ( 
.A(n_5637),
.Y(n_6197)
);

CKINVDCx5p33_ASAP7_75t_R g6198 ( 
.A(n_5757),
.Y(n_6198)
);

CKINVDCx5p33_ASAP7_75t_R g6199 ( 
.A(n_5423),
.Y(n_6199)
);

INVx2_ASAP7_75t_L g6200 ( 
.A(n_5534),
.Y(n_6200)
);

NAND3xp33_ASAP7_75t_L g6201 ( 
.A(n_5401),
.B(n_5565),
.C(n_5528),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_5535),
.Y(n_6202)
);

BUFx6f_ASAP7_75t_L g6203 ( 
.A(n_5343),
.Y(n_6203)
);

CKINVDCx20_ASAP7_75t_R g6204 ( 
.A(n_5636),
.Y(n_6204)
);

CKINVDCx5p33_ASAP7_75t_R g6205 ( 
.A(n_5641),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5536),
.Y(n_6206)
);

INVx1_ASAP7_75t_SL g6207 ( 
.A(n_5588),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_5784),
.B(n_3100),
.Y(n_6208)
);

CKINVDCx5p33_ASAP7_75t_R g6209 ( 
.A(n_5645),
.Y(n_6209)
);

CKINVDCx20_ASAP7_75t_R g6210 ( 
.A(n_5647),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_5537),
.Y(n_6211)
);

CKINVDCx5p33_ASAP7_75t_R g6212 ( 
.A(n_5649),
.Y(n_6212)
);

CKINVDCx5p33_ASAP7_75t_R g6213 ( 
.A(n_5453),
.Y(n_6213)
);

OR2x2_ASAP7_75t_L g6214 ( 
.A(n_5769),
.B(n_3101),
.Y(n_6214)
);

CKINVDCx5p33_ASAP7_75t_R g6215 ( 
.A(n_5625),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5539),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_5541),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_5626),
.Y(n_6218)
);

CKINVDCx5p33_ASAP7_75t_R g6219 ( 
.A(n_5437),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_5295),
.Y(n_6220)
);

NOR2xp33_ASAP7_75t_R g6221 ( 
.A(n_5448),
.B(n_5245),
.Y(n_6221)
);

AND2x2_ASAP7_75t_L g6222 ( 
.A(n_5321),
.B(n_4189),
.Y(n_6222)
);

CKINVDCx5p33_ASAP7_75t_R g6223 ( 
.A(n_5628),
.Y(n_6223)
);

CKINVDCx5p33_ASAP7_75t_R g6224 ( 
.A(n_5440),
.Y(n_6224)
);

CKINVDCx5p33_ASAP7_75t_R g6225 ( 
.A(n_5573),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_5552),
.Y(n_6226)
);

CKINVDCx5p33_ASAP7_75t_R g6227 ( 
.A(n_5607),
.Y(n_6227)
);

NOR2xp33_ASAP7_75t_L g6228 ( 
.A(n_5237),
.B(n_3103),
.Y(n_6228)
);

CKINVDCx5p33_ASAP7_75t_R g6229 ( 
.A(n_5615),
.Y(n_6229)
);

NAND2xp5_ASAP7_75t_SL g6230 ( 
.A(n_5323),
.B(n_3105),
.Y(n_6230)
);

CKINVDCx5p33_ASAP7_75t_R g6231 ( 
.A(n_5624),
.Y(n_6231)
);

INVxp67_ASAP7_75t_L g6232 ( 
.A(n_5605),
.Y(n_6232)
);

HB1xp67_ASAP7_75t_L g6233 ( 
.A(n_5666),
.Y(n_6233)
);

AOI22xp5_ASAP7_75t_L g6234 ( 
.A1(n_5241),
.A2(n_4229),
.B1(n_4231),
.B2(n_4225),
.Y(n_6234)
);

INVx3_ASAP7_75t_L g6235 ( 
.A(n_5775),
.Y(n_6235)
);

NOR2xp67_ASAP7_75t_L g6236 ( 
.A(n_5249),
.B(n_3111),
.Y(n_6236)
);

CKINVDCx5p33_ASAP7_75t_R g6237 ( 
.A(n_5315),
.Y(n_6237)
);

NOR2xp33_ASAP7_75t_R g6238 ( 
.A(n_5745),
.B(n_4244),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_5567),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_5316),
.Y(n_6240)
);

INVx2_ASAP7_75t_L g6241 ( 
.A(n_5569),
.Y(n_6241)
);

CKINVDCx5p33_ASAP7_75t_R g6242 ( 
.A(n_5279),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5575),
.Y(n_6243)
);

CKINVDCx20_ASAP7_75t_R g6244 ( 
.A(n_5391),
.Y(n_6244)
);

CKINVDCx5p33_ASAP7_75t_R g6245 ( 
.A(n_5373),
.Y(n_6245)
);

AND2x6_ASAP7_75t_L g6246 ( 
.A(n_5412),
.B(n_3427),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_5576),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5577),
.Y(n_6248)
);

CKINVDCx5p33_ASAP7_75t_R g6249 ( 
.A(n_5611),
.Y(n_6249)
);

CKINVDCx5p33_ASAP7_75t_R g6250 ( 
.A(n_5424),
.Y(n_6250)
);

CKINVDCx20_ASAP7_75t_R g6251 ( 
.A(n_5509),
.Y(n_6251)
);

CKINVDCx20_ASAP7_75t_R g6252 ( 
.A(n_5566),
.Y(n_6252)
);

INVx2_ASAP7_75t_L g6253 ( 
.A(n_5582),
.Y(n_6253)
);

HB1xp67_ASAP7_75t_L g6254 ( 
.A(n_5682),
.Y(n_6254)
);

INVx3_ASAP7_75t_L g6255 ( 
.A(n_5780),
.Y(n_6255)
);

CKINVDCx16_ASAP7_75t_R g6256 ( 
.A(n_5732),
.Y(n_6256)
);

CKINVDCx5p33_ASAP7_75t_R g6257 ( 
.A(n_5603),
.Y(n_6257)
);

BUFx3_ASAP7_75t_L g6258 ( 
.A(n_5347),
.Y(n_6258)
);

CKINVDCx5p33_ASAP7_75t_R g6259 ( 
.A(n_5609),
.Y(n_6259)
);

CKINVDCx5p33_ASAP7_75t_R g6260 ( 
.A(n_5610),
.Y(n_6260)
);

INVx1_ASAP7_75t_L g6261 ( 
.A(n_5591),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_5746),
.Y(n_6262)
);

AND2x2_ASAP7_75t_L g6263 ( 
.A(n_5469),
.B(n_4249),
.Y(n_6263)
);

NOR2xp33_ASAP7_75t_R g6264 ( 
.A(n_5747),
.B(n_4252),
.Y(n_6264)
);

AOI22xp5_ASAP7_75t_L g6265 ( 
.A1(n_5251),
.A2(n_4295),
.B1(n_3112),
.B2(n_3114),
.Y(n_6265)
);

CKINVDCx20_ASAP7_75t_R g6266 ( 
.A(n_5574),
.Y(n_6266)
);

CKINVDCx5p33_ASAP7_75t_R g6267 ( 
.A(n_5612),
.Y(n_6267)
);

CKINVDCx5p33_ASAP7_75t_R g6268 ( 
.A(n_5547),
.Y(n_6268)
);

CKINVDCx5p33_ASAP7_75t_R g6269 ( 
.A(n_5581),
.Y(n_6269)
);

INVx2_ASAP7_75t_L g6270 ( 
.A(n_5781),
.Y(n_6270)
);

CKINVDCx5p33_ASAP7_75t_R g6271 ( 
.A(n_5586),
.Y(n_6271)
);

CKINVDCx5p33_ASAP7_75t_R g6272 ( 
.A(n_5618),
.Y(n_6272)
);

INVx3_ASAP7_75t_L g6273 ( 
.A(n_5782),
.Y(n_6273)
);

INVx3_ASAP7_75t_L g6274 ( 
.A(n_5788),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5748),
.Y(n_6275)
);

CKINVDCx20_ASAP7_75t_R g6276 ( 
.A(n_5387),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_5792),
.Y(n_6277)
);

CKINVDCx5p33_ASAP7_75t_R g6278 ( 
.A(n_5422),
.Y(n_6278)
);

CKINVDCx16_ASAP7_75t_R g6279 ( 
.A(n_5243),
.Y(n_6279)
);

CKINVDCx5p33_ASAP7_75t_R g6280 ( 
.A(n_5425),
.Y(n_6280)
);

OR2x2_ASAP7_75t_L g6281 ( 
.A(n_5289),
.B(n_3113),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_5752),
.Y(n_6282)
);

CKINVDCx5p33_ASAP7_75t_R g6283 ( 
.A(n_5760),
.Y(n_6283)
);

BUFx6f_ASAP7_75t_L g6284 ( 
.A(n_5352),
.Y(n_6284)
);

AND2x2_ASAP7_75t_L g6285 ( 
.A(n_5266),
.B(n_3115),
.Y(n_6285)
);

BUFx3_ASAP7_75t_L g6286 ( 
.A(n_5761),
.Y(n_6286)
);

CKINVDCx5p33_ASAP7_75t_R g6287 ( 
.A(n_5764),
.Y(n_6287)
);

NOR2xp33_ASAP7_75t_SL g6288 ( 
.A(n_5771),
.B(n_3117),
.Y(n_6288)
);

CKINVDCx5p33_ASAP7_75t_R g6289 ( 
.A(n_5772),
.Y(n_6289)
);

INVx3_ASAP7_75t_L g6290 ( 
.A(n_5797),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5778),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_5789),
.Y(n_6292)
);

CKINVDCx5p33_ASAP7_75t_R g6293 ( 
.A(n_5800),
.Y(n_6293)
);

HB1xp67_ASAP7_75t_L g6294 ( 
.A(n_5804),
.Y(n_6294)
);

NAND2xp5_ASAP7_75t_L g6295 ( 
.A(n_5442),
.B(n_3118),
.Y(n_6295)
);

CKINVDCx5p33_ASAP7_75t_R g6296 ( 
.A(n_5806),
.Y(n_6296)
);

INVx1_ASAP7_75t_SL g6297 ( 
.A(n_5768),
.Y(n_6297)
);

NOR2xp33_ASAP7_75t_L g6298 ( 
.A(n_5336),
.B(n_5346),
.Y(n_6298)
);

HB1xp67_ASAP7_75t_L g6299 ( 
.A(n_5773),
.Y(n_6299)
);

BUFx2_ASAP7_75t_L g6300 ( 
.A(n_5733),
.Y(n_6300)
);

CKINVDCx5p33_ASAP7_75t_R g6301 ( 
.A(n_5441),
.Y(n_6301)
);

AND2x6_ASAP7_75t_L g6302 ( 
.A(n_5545),
.B(n_3430),
.Y(n_6302)
);

NOR2xp33_ASAP7_75t_R g6303 ( 
.A(n_5250),
.B(n_3122),
.Y(n_6303)
);

AND2x4_ASAP7_75t_L g6304 ( 
.A(n_5312),
.B(n_5799),
.Y(n_6304)
);

CKINVDCx5p33_ASAP7_75t_R g6305 ( 
.A(n_5446),
.Y(n_6305)
);

HB1xp67_ASAP7_75t_L g6306 ( 
.A(n_5787),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5519),
.Y(n_6307)
);

CKINVDCx5p33_ASAP7_75t_R g6308 ( 
.A(n_5447),
.Y(n_6308)
);

CKINVDCx5p33_ASAP7_75t_R g6309 ( 
.A(n_5449),
.Y(n_6309)
);

CKINVDCx5p33_ASAP7_75t_R g6310 ( 
.A(n_5450),
.Y(n_6310)
);

CKINVDCx5p33_ASAP7_75t_R g6311 ( 
.A(n_5451),
.Y(n_6311)
);

CKINVDCx5p33_ASAP7_75t_R g6312 ( 
.A(n_5456),
.Y(n_6312)
);

AND3x2_ASAP7_75t_L g6313 ( 
.A(n_5791),
.B(n_3437),
.C(n_3433),
.Y(n_6313)
);

CKINVDCx5p33_ASAP7_75t_R g6314 ( 
.A(n_5464),
.Y(n_6314)
);

CKINVDCx5p33_ASAP7_75t_R g6315 ( 
.A(n_5470),
.Y(n_6315)
);

INVx2_ASAP7_75t_L g6316 ( 
.A(n_5801),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_5529),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_5530),
.Y(n_6318)
);

HB1xp67_ASAP7_75t_L g6319 ( 
.A(n_5807),
.Y(n_6319)
);

CKINVDCx5p33_ASAP7_75t_R g6320 ( 
.A(n_5498),
.Y(n_6320)
);

CKINVDCx5p33_ASAP7_75t_R g6321 ( 
.A(n_5517),
.Y(n_6321)
);

NOR2xp33_ASAP7_75t_R g6322 ( 
.A(n_5261),
.B(n_3128),
.Y(n_6322)
);

INVx2_ASAP7_75t_L g6323 ( 
.A(n_5811),
.Y(n_6323)
);

NAND2xp33_ASAP7_75t_R g6324 ( 
.A(n_5578),
.B(n_3130),
.Y(n_6324)
);

CKINVDCx20_ASAP7_75t_R g6325 ( 
.A(n_5623),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_5555),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5570),
.Y(n_6327)
);

INVx2_ASAP7_75t_L g6328 ( 
.A(n_5399),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5571),
.Y(n_6329)
);

CKINVDCx5p33_ASAP7_75t_R g6330 ( 
.A(n_5549),
.Y(n_6330)
);

NOR2xp67_ASAP7_75t_L g6331 ( 
.A(n_5348),
.B(n_3131),
.Y(n_6331)
);

CKINVDCx5p33_ASAP7_75t_R g6332 ( 
.A(n_5554),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_5579),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_5589),
.Y(n_6334)
);

CKINVDCx5p33_ASAP7_75t_R g6335 ( 
.A(n_5593),
.Y(n_6335)
);

BUFx2_ASAP7_75t_L g6336 ( 
.A(n_5812),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_5485),
.Y(n_6337)
);

BUFx10_ASAP7_75t_L g6338 ( 
.A(n_5622),
.Y(n_6338)
);

BUFx2_ASAP7_75t_L g6339 ( 
.A(n_5303),
.Y(n_6339)
);

INVx3_ASAP7_75t_L g6340 ( 
.A(n_5585),
.Y(n_6340)
);

BUFx8_ASAP7_75t_L g6341 ( 
.A(n_5366),
.Y(n_6341)
);

HB1xp67_ASAP7_75t_L g6342 ( 
.A(n_5383),
.Y(n_6342)
);

CKINVDCx20_ASAP7_75t_R g6343 ( 
.A(n_5523),
.Y(n_6343)
);

CKINVDCx5p33_ASAP7_75t_R g6344 ( 
.A(n_5380),
.Y(n_6344)
);

HB1xp67_ASAP7_75t_L g6345 ( 
.A(n_5385),
.Y(n_6345)
);

BUFx2_ASAP7_75t_L g6346 ( 
.A(n_5395),
.Y(n_6346)
);

CKINVDCx16_ASAP7_75t_R g6347 ( 
.A(n_5404),
.Y(n_6347)
);

CKINVDCx5p33_ASAP7_75t_R g6348 ( 
.A(n_5386),
.Y(n_6348)
);

CKINVDCx5p33_ASAP7_75t_R g6349 ( 
.A(n_5400),
.Y(n_6349)
);

INVx1_ASAP7_75t_SL g6350 ( 
.A(n_5410),
.Y(n_6350)
);

CKINVDCx5p33_ASAP7_75t_R g6351 ( 
.A(n_5421),
.Y(n_6351)
);

CKINVDCx5p33_ASAP7_75t_R g6352 ( 
.A(n_5430),
.Y(n_6352)
);

CKINVDCx5p33_ASAP7_75t_R g6353 ( 
.A(n_5435),
.Y(n_6353)
);

CKINVDCx5p33_ASAP7_75t_R g6354 ( 
.A(n_5444),
.Y(n_6354)
);

NOR2xp33_ASAP7_75t_L g6355 ( 
.A(n_5292),
.B(n_3132),
.Y(n_6355)
);

NAND2xp5_ASAP7_75t_SL g6356 ( 
.A(n_5479),
.B(n_3134),
.Y(n_6356)
);

CKINVDCx5p33_ASAP7_75t_R g6357 ( 
.A(n_5500),
.Y(n_6357)
);

CKINVDCx16_ASAP7_75t_R g6358 ( 
.A(n_5521),
.Y(n_6358)
);

CKINVDCx14_ASAP7_75t_R g6359 ( 
.A(n_5458),
.Y(n_6359)
);

CKINVDCx5p33_ASAP7_75t_R g6360 ( 
.A(n_5802),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5434),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5477),
.Y(n_6362)
);

CKINVDCx5p33_ASAP7_75t_R g6363 ( 
.A(n_5803),
.Y(n_6363)
);

CKINVDCx5p33_ASAP7_75t_R g6364 ( 
.A(n_5270),
.Y(n_6364)
);

NOR2xp33_ASAP7_75t_R g6365 ( 
.A(n_5287),
.B(n_3135),
.Y(n_6365)
);

CKINVDCx5p33_ASAP7_75t_R g6366 ( 
.A(n_5462),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_5463),
.Y(n_6367)
);

CKINVDCx5p33_ASAP7_75t_R g6368 ( 
.A(n_5471),
.Y(n_6368)
);

CKINVDCx5p33_ASAP7_75t_R g6369 ( 
.A(n_5482),
.Y(n_6369)
);

INVx2_ASAP7_75t_L g6370 ( 
.A(n_5300),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_5484),
.Y(n_6371)
);

CKINVDCx5p33_ASAP7_75t_R g6372 ( 
.A(n_5502),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_5507),
.Y(n_6373)
);

NAND2xp5_ASAP7_75t_L g6374 ( 
.A(n_6298),
.B(n_5617),
.Y(n_6374)
);

CKINVDCx5p33_ASAP7_75t_R g6375 ( 
.A(n_5816),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_SL g6376 ( 
.A(n_6269),
.B(n_5627),
.Y(n_6376)
);

NAND2x1p5_ASAP7_75t_L g6377 ( 
.A(n_5959),
.B(n_5583),
.Y(n_6377)
);

NOR2xp33_ASAP7_75t_L g6378 ( 
.A(n_6052),
.B(n_5356),
.Y(n_6378)
);

AND2x4_ASAP7_75t_L g6379 ( 
.A(n_5835),
.B(n_5767),
.Y(n_6379)
);

INVx4_ASAP7_75t_SL g6380 ( 
.A(n_5834),
.Y(n_6380)
);

NOR2xp33_ASAP7_75t_L g6381 ( 
.A(n_5855),
.B(n_5359),
.Y(n_6381)
);

INVx2_ASAP7_75t_L g6382 ( 
.A(n_5829),
.Y(n_6382)
);

BUFx10_ASAP7_75t_L g6383 ( 
.A(n_5817),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_5832),
.Y(n_6384)
);

INVx2_ASAP7_75t_SL g6385 ( 
.A(n_5814),
.Y(n_6385)
);

BUFx4f_ASAP7_75t_L g6386 ( 
.A(n_6025),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_SL g6387 ( 
.A(n_6271),
.B(n_5363),
.Y(n_6387)
);

NAND2xp5_ASAP7_75t_L g6388 ( 
.A(n_6367),
.B(n_5367),
.Y(n_6388)
);

BUFx6f_ASAP7_75t_L g6389 ( 
.A(n_5834),
.Y(n_6389)
);

BUFx2_ASAP7_75t_L g6390 ( 
.A(n_6039),
.Y(n_6390)
);

BUFx3_ASAP7_75t_L g6391 ( 
.A(n_6344),
.Y(n_6391)
);

NAND2xp5_ASAP7_75t_L g6392 ( 
.A(n_6371),
.B(n_5372),
.Y(n_6392)
);

BUFx2_ASAP7_75t_L g6393 ( 
.A(n_5995),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_5833),
.Y(n_6394)
);

BUFx3_ASAP7_75t_L g6395 ( 
.A(n_6348),
.Y(n_6395)
);

INVxp33_ASAP7_75t_L g6396 ( 
.A(n_6238),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_5823),
.Y(n_6397)
);

NOR2xp33_ASAP7_75t_L g6398 ( 
.A(n_6337),
.B(n_5393),
.Y(n_6398)
);

NOR2xp33_ASAP7_75t_L g6399 ( 
.A(n_6156),
.B(n_6158),
.Y(n_6399)
);

BUFx4f_ASAP7_75t_L g6400 ( 
.A(n_5980),
.Y(n_6400)
);

INVx2_ASAP7_75t_SL g6401 ( 
.A(n_6249),
.Y(n_6401)
);

OR2x6_ASAP7_75t_L g6402 ( 
.A(n_5980),
.B(n_5406),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_5864),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_6373),
.B(n_5465),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_6057),
.B(n_5639),
.Y(n_6405)
);

BUFx2_ASAP7_75t_L g6406 ( 
.A(n_5836),
.Y(n_6406)
);

NOR2x1p5_ASAP7_75t_L g6407 ( 
.A(n_5937),
.B(n_3138),
.Y(n_6407)
);

INVx5_ASAP7_75t_L g6408 ( 
.A(n_6088),
.Y(n_6408)
);

INVx5_ASAP7_75t_L g6409 ( 
.A(n_6088),
.Y(n_6409)
);

BUFx2_ASAP7_75t_L g6410 ( 
.A(n_5982),
.Y(n_6410)
);

NAND2xp5_ASAP7_75t_SL g6411 ( 
.A(n_6272),
.B(n_5640),
.Y(n_6411)
);

INVxp67_ASAP7_75t_SL g6412 ( 
.A(n_6106),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_5880),
.Y(n_6413)
);

OAI22xp33_ASAP7_75t_L g6414 ( 
.A1(n_6065),
.A2(n_3139),
.B1(n_3144),
.B2(n_3141),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5826),
.Y(n_6415)
);

INVxp67_ASAP7_75t_SL g6416 ( 
.A(n_5973),
.Y(n_6416)
);

NAND2xp5_ASAP7_75t_L g6417 ( 
.A(n_5875),
.B(n_5483),
.Y(n_6417)
);

INVx6_ASAP7_75t_L g6418 ( 
.A(n_6151),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_6366),
.B(n_5505),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5843),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6368),
.B(n_5283),
.Y(n_6421)
);

INVx4_ASAP7_75t_L g6422 ( 
.A(n_6301),
.Y(n_6422)
);

NOR2xp33_ASAP7_75t_L g6423 ( 
.A(n_5949),
.B(n_3149),
.Y(n_6423)
);

AND2x2_ASAP7_75t_L g6424 ( 
.A(n_5852),
.B(n_3152),
.Y(n_6424)
);

INVx2_ASAP7_75t_L g6425 ( 
.A(n_5889),
.Y(n_6425)
);

NAND2xp5_ASAP7_75t_SL g6426 ( 
.A(n_6369),
.B(n_3153),
.Y(n_6426)
);

BUFx2_ASAP7_75t_L g6427 ( 
.A(n_5872),
.Y(n_6427)
);

INVx2_ASAP7_75t_SL g6428 ( 
.A(n_6267),
.Y(n_6428)
);

INVx2_ASAP7_75t_L g6429 ( 
.A(n_5895),
.Y(n_6429)
);

CKINVDCx5p33_ASAP7_75t_R g6430 ( 
.A(n_5818),
.Y(n_6430)
);

NOR2xp33_ASAP7_75t_L g6431 ( 
.A(n_6372),
.B(n_3158),
.Y(n_6431)
);

INVxp67_ASAP7_75t_L g6432 ( 
.A(n_5815),
.Y(n_6432)
);

NOR2xp33_ASAP7_75t_L g6433 ( 
.A(n_6150),
.B(n_3159),
.Y(n_6433)
);

NAND2xp5_ASAP7_75t_SL g6434 ( 
.A(n_6278),
.B(n_3163),
.Y(n_6434)
);

NAND2xp5_ASAP7_75t_L g6435 ( 
.A(n_6102),
.B(n_5327),
.Y(n_6435)
);

NAND2xp5_ASAP7_75t_SL g6436 ( 
.A(n_6280),
.B(n_3164),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_5844),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5856),
.Y(n_6438)
);

BUFx6f_ASAP7_75t_L g6439 ( 
.A(n_5834),
.Y(n_6439)
);

CKINVDCx5p33_ASAP7_75t_R g6440 ( 
.A(n_5819),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_5901),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_5882),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5884),
.Y(n_6443)
);

AO22x2_ASAP7_75t_L g6444 ( 
.A1(n_5961),
.A2(n_3442),
.B1(n_3448),
.B2(n_3439),
.Y(n_6444)
);

BUFx3_ASAP7_75t_L g6445 ( 
.A(n_6349),
.Y(n_6445)
);

OR2x6_ASAP7_75t_L g6446 ( 
.A(n_6196),
.B(n_5376),
.Y(n_6446)
);

INVx2_ASAP7_75t_L g6447 ( 
.A(n_5912),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_5886),
.Y(n_6448)
);

INVx4_ASAP7_75t_L g6449 ( 
.A(n_6305),
.Y(n_6449)
);

NOR2xp33_ASAP7_75t_L g6450 ( 
.A(n_6207),
.B(n_3165),
.Y(n_6450)
);

INVxp33_ASAP7_75t_L g6451 ( 
.A(n_6264),
.Y(n_6451)
);

INVx3_ASAP7_75t_L g6452 ( 
.A(n_5879),
.Y(n_6452)
);

AND2x6_ASAP7_75t_L g6453 ( 
.A(n_6285),
.B(n_3452),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_5897),
.Y(n_6454)
);

INVx2_ASAP7_75t_SL g6455 ( 
.A(n_6151),
.Y(n_6455)
);

INVx3_ASAP7_75t_L g6456 ( 
.A(n_5879),
.Y(n_6456)
);

INVx1_ASAP7_75t_SL g6457 ( 
.A(n_5865),
.Y(n_6457)
);

NOR2xp33_ASAP7_75t_L g6458 ( 
.A(n_6070),
.B(n_3168),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5900),
.Y(n_6459)
);

AND2x4_ASAP7_75t_L g6460 ( 
.A(n_5866),
.B(n_3460),
.Y(n_6460)
);

INVx2_ASAP7_75t_SL g6461 ( 
.A(n_6286),
.Y(n_6461)
);

BUFx3_ASAP7_75t_L g6462 ( 
.A(n_6351),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5908),
.Y(n_6463)
);

BUFx6f_ASAP7_75t_L g6464 ( 
.A(n_5879),
.Y(n_6464)
);

INVx3_ASAP7_75t_L g6465 ( 
.A(n_5960),
.Y(n_6465)
);

INVx4_ASAP7_75t_L g6466 ( 
.A(n_6308),
.Y(n_6466)
);

INVx2_ASAP7_75t_L g6467 ( 
.A(n_5936),
.Y(n_6467)
);

INVx3_ASAP7_75t_L g6468 ( 
.A(n_5960),
.Y(n_6468)
);

NAND2xp5_ASAP7_75t_L g6469 ( 
.A(n_6127),
.B(n_3169),
.Y(n_6469)
);

INVxp67_ASAP7_75t_SL g6470 ( 
.A(n_6004),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_5943),
.Y(n_6471)
);

BUFx6f_ASAP7_75t_L g6472 ( 
.A(n_5960),
.Y(n_6472)
);

BUFx3_ASAP7_75t_L g6473 ( 
.A(n_6352),
.Y(n_6473)
);

AOI22xp33_ASAP7_75t_L g6474 ( 
.A1(n_6361),
.A2(n_3465),
.B1(n_3469),
.B2(n_3461),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_5915),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_5916),
.Y(n_6476)
);

NAND2xp5_ASAP7_75t_L g6477 ( 
.A(n_5898),
.B(n_3170),
.Y(n_6477)
);

NAND2xp5_ASAP7_75t_L g6478 ( 
.A(n_6050),
.B(n_3172),
.Y(n_6478)
);

INVx2_ASAP7_75t_SL g6479 ( 
.A(n_6309),
.Y(n_6479)
);

INVx4_ASAP7_75t_SL g6480 ( 
.A(n_5983),
.Y(n_6480)
);

INVx2_ASAP7_75t_L g6481 ( 
.A(n_5918),
.Y(n_6481)
);

NOR2xp33_ASAP7_75t_L g6482 ( 
.A(n_6020),
.B(n_3173),
.Y(n_6482)
);

NOR2xp33_ASAP7_75t_L g6483 ( 
.A(n_6044),
.B(n_6077),
.Y(n_6483)
);

AOI22xp33_ASAP7_75t_L g6484 ( 
.A1(n_6201),
.A2(n_3476),
.B1(n_3483),
.B2(n_3475),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6228),
.B(n_3180),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_5919),
.Y(n_6486)
);

OR2x6_ASAP7_75t_L g6487 ( 
.A(n_6196),
.B(n_3490),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_5920),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_5923),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_5926),
.Y(n_6490)
);

NAND2xp5_ASAP7_75t_L g6491 ( 
.A(n_5963),
.B(n_3184),
.Y(n_6491)
);

INVx3_ASAP7_75t_L g6492 ( 
.A(n_5983),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_SL g6493 ( 
.A(n_6089),
.B(n_3187),
.Y(n_6493)
);

INVx5_ASAP7_75t_L g6494 ( 
.A(n_5983),
.Y(n_6494)
);

NAND2xp5_ASAP7_75t_L g6495 ( 
.A(n_6173),
.B(n_3191),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_5931),
.Y(n_6496)
);

INVx5_ASAP7_75t_L g6497 ( 
.A(n_6003),
.Y(n_6497)
);

INVx3_ASAP7_75t_L g6498 ( 
.A(n_6003),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_5933),
.Y(n_6499)
);

OR2x2_ASAP7_75t_L g6500 ( 
.A(n_6116),
.B(n_3193),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_5941),
.Y(n_6501)
);

NOR2xp33_ASAP7_75t_L g6502 ( 
.A(n_6096),
.B(n_3194),
.Y(n_6502)
);

INVx3_ASAP7_75t_L g6503 ( 
.A(n_6003),
.Y(n_6503)
);

INVxp67_ASAP7_75t_L g6504 ( 
.A(n_5839),
.Y(n_6504)
);

HB1xp67_ASAP7_75t_L g6505 ( 
.A(n_5867),
.Y(n_6505)
);

INVx1_ASAP7_75t_L g6506 ( 
.A(n_5951),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5957),
.Y(n_6507)
);

INVx2_ASAP7_75t_SL g6508 ( 
.A(n_6310),
.Y(n_6508)
);

INVx4_ASAP7_75t_SL g6509 ( 
.A(n_6030),
.Y(n_6509)
);

INVx2_ASAP7_75t_L g6510 ( 
.A(n_5962),
.Y(n_6510)
);

NAND2xp5_ASAP7_75t_L g6511 ( 
.A(n_6175),
.B(n_3198),
.Y(n_6511)
);

INVx4_ASAP7_75t_L g6512 ( 
.A(n_6311),
.Y(n_6512)
);

OR2x2_ASAP7_75t_L g6513 ( 
.A(n_5956),
.B(n_3199),
.Y(n_6513)
);

NAND2xp5_ASAP7_75t_L g6514 ( 
.A(n_6177),
.B(n_3201),
.Y(n_6514)
);

NOR2x1p5_ASAP7_75t_L g6515 ( 
.A(n_5953),
.B(n_3203),
.Y(n_6515)
);

INVx5_ASAP7_75t_L g6516 ( 
.A(n_6030),
.Y(n_6516)
);

INVx2_ASAP7_75t_L g6517 ( 
.A(n_5970),
.Y(n_6517)
);

INVx4_ASAP7_75t_L g6518 ( 
.A(n_6312),
.Y(n_6518)
);

AOI22xp33_ASAP7_75t_L g6519 ( 
.A1(n_5902),
.A2(n_3500),
.B1(n_3501),
.B2(n_3497),
.Y(n_6519)
);

BUFx6f_ASAP7_75t_L g6520 ( 
.A(n_6030),
.Y(n_6520)
);

NAND2xp5_ASAP7_75t_L g6521 ( 
.A(n_6178),
.B(n_3210),
.Y(n_6521)
);

NAND2xp5_ASAP7_75t_SL g6522 ( 
.A(n_6085),
.B(n_6354),
.Y(n_6522)
);

OR2x2_ASAP7_75t_L g6523 ( 
.A(n_5869),
.B(n_3211),
.Y(n_6523)
);

BUFx2_ASAP7_75t_L g6524 ( 
.A(n_5876),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_L g6525 ( 
.A(n_6181),
.B(n_3212),
.Y(n_6525)
);

OR2x2_ASAP7_75t_L g6526 ( 
.A(n_6145),
.B(n_6174),
.Y(n_6526)
);

AOI22xp33_ASAP7_75t_L g6527 ( 
.A1(n_5965),
.A2(n_3508),
.B1(n_3510),
.B2(n_3507),
.Y(n_6527)
);

INVx2_ASAP7_75t_SL g6528 ( 
.A(n_6314),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_5964),
.B(n_3217),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_5978),
.Y(n_6530)
);

BUFx6f_ASAP7_75t_L g6531 ( 
.A(n_6068),
.Y(n_6531)
);

BUFx6f_ASAP7_75t_L g6532 ( 
.A(n_6068),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_6183),
.B(n_3222),
.Y(n_6533)
);

NAND2xp5_ASAP7_75t_SL g6534 ( 
.A(n_6135),
.B(n_3223),
.Y(n_6534)
);

BUFx8_ASAP7_75t_SL g6535 ( 
.A(n_5840),
.Y(n_6535)
);

INVx1_ASAP7_75t_SL g6536 ( 
.A(n_6128),
.Y(n_6536)
);

NAND2xp5_ASAP7_75t_L g6537 ( 
.A(n_6186),
.B(n_3226),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_5989),
.Y(n_6538)
);

INVx1_ASAP7_75t_SL g6539 ( 
.A(n_6129),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_6149),
.B(n_3229),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_5990),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_6193),
.B(n_3232),
.Y(n_6542)
);

HB1xp67_ASAP7_75t_L g6543 ( 
.A(n_6294),
.Y(n_6543)
);

AND2x2_ASAP7_75t_L g6544 ( 
.A(n_6037),
.B(n_3235),
.Y(n_6544)
);

INVx3_ASAP7_75t_L g6545 ( 
.A(n_6068),
.Y(n_6545)
);

INVxp67_ASAP7_75t_L g6546 ( 
.A(n_6355),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_5994),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_5996),
.Y(n_6548)
);

AND2x4_ASAP7_75t_L g6549 ( 
.A(n_5924),
.B(n_3514),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_5921),
.B(n_3236),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_6006),
.Y(n_6551)
);

INVx3_ASAP7_75t_L g6552 ( 
.A(n_6111),
.Y(n_6552)
);

AOI22xp5_ASAP7_75t_L g6553 ( 
.A1(n_6325),
.A2(n_3251),
.B1(n_3252),
.B2(n_3240),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6008),
.Y(n_6554)
);

AOI22xp33_ASAP7_75t_L g6555 ( 
.A1(n_6233),
.A2(n_3527),
.B1(n_3531),
.B2(n_3515),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6010),
.Y(n_6556)
);

INVx1_ASAP7_75t_SL g6557 ( 
.A(n_6064),
.Y(n_6557)
);

AOI22xp33_ASAP7_75t_L g6558 ( 
.A1(n_6254),
.A2(n_3533),
.B1(n_3538),
.B2(n_3532),
.Y(n_6558)
);

AND2x6_ASAP7_75t_L g6559 ( 
.A(n_6350),
.B(n_6362),
.Y(n_6559)
);

INVx4_ASAP7_75t_L g6560 ( 
.A(n_6315),
.Y(n_6560)
);

NOR2xp33_ASAP7_75t_L g6561 ( 
.A(n_6189),
.B(n_3256),
.Y(n_6561)
);

BUFx10_ASAP7_75t_L g6562 ( 
.A(n_5820),
.Y(n_6562)
);

BUFx2_ASAP7_75t_L g6563 ( 
.A(n_5892),
.Y(n_6563)
);

NOR2xp33_ASAP7_75t_L g6564 ( 
.A(n_6232),
.B(n_3257),
.Y(n_6564)
);

AND2x6_ASAP7_75t_L g6565 ( 
.A(n_6263),
.B(n_3541),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_6029),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_SL g6567 ( 
.A(n_6137),
.B(n_3259),
.Y(n_6567)
);

INVx4_ASAP7_75t_SL g6568 ( 
.A(n_6111),
.Y(n_6568)
);

INVx2_ASAP7_75t_L g6569 ( 
.A(n_6032),
.Y(n_6569)
);

AND2x4_ASAP7_75t_L g6570 ( 
.A(n_6171),
.B(n_3550),
.Y(n_6570)
);

NOR2xp33_ASAP7_75t_L g6571 ( 
.A(n_6257),
.B(n_6259),
.Y(n_6571)
);

BUFx10_ASAP7_75t_L g6572 ( 
.A(n_5821),
.Y(n_6572)
);

NAND2xp5_ASAP7_75t_L g6573 ( 
.A(n_6187),
.B(n_3260),
.Y(n_6573)
);

BUFx2_ASAP7_75t_L g6574 ( 
.A(n_6018),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6042),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6045),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6046),
.Y(n_6577)
);

INVx6_ASAP7_75t_L g6578 ( 
.A(n_6279),
.Y(n_6578)
);

INVx3_ASAP7_75t_L g6579 ( 
.A(n_6111),
.Y(n_6579)
);

INVx4_ASAP7_75t_L g6580 ( 
.A(n_6320),
.Y(n_6580)
);

NAND2xp33_ASAP7_75t_SL g6581 ( 
.A(n_5878),
.B(n_3267),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6047),
.Y(n_6582)
);

AND2x2_ASAP7_75t_SL g6583 ( 
.A(n_6163),
.B(n_6043),
.Y(n_6583)
);

AOI22xp33_ASAP7_75t_L g6584 ( 
.A1(n_6191),
.A2(n_3561),
.B1(n_3562),
.B2(n_3556),
.Y(n_6584)
);

INVx1_ASAP7_75t_SL g6585 ( 
.A(n_5917),
.Y(n_6585)
);

INVx4_ASAP7_75t_L g6586 ( 
.A(n_6321),
.Y(n_6586)
);

OAI22xp5_ASAP7_75t_L g6587 ( 
.A1(n_6213),
.A2(n_3271),
.B1(n_3272),
.B2(n_3269),
.Y(n_6587)
);

CKINVDCx16_ASAP7_75t_R g6588 ( 
.A(n_5831),
.Y(n_6588)
);

BUFx10_ASAP7_75t_L g6589 ( 
.A(n_5822),
.Y(n_6589)
);

INVx3_ASAP7_75t_L g6590 ( 
.A(n_6113),
.Y(n_6590)
);

INVx1_ASAP7_75t_L g6591 ( 
.A(n_6051),
.Y(n_6591)
);

CKINVDCx20_ASAP7_75t_R g6592 ( 
.A(n_5827),
.Y(n_6592)
);

INVx1_ASAP7_75t_SL g6593 ( 
.A(n_5922),
.Y(n_6593)
);

AOI22xp33_ASAP7_75t_SL g6594 ( 
.A1(n_6021),
.A2(n_3276),
.B1(n_3278),
.B2(n_3275),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6060),
.Y(n_6595)
);

INVx2_ASAP7_75t_SL g6596 ( 
.A(n_6330),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6081),
.Y(n_6597)
);

BUFx3_ASAP7_75t_L g6598 ( 
.A(n_6237),
.Y(n_6598)
);

INVx1_ASAP7_75t_SL g6599 ( 
.A(n_6332),
.Y(n_6599)
);

BUFx10_ASAP7_75t_L g6600 ( 
.A(n_5824),
.Y(n_6600)
);

CKINVDCx5p33_ASAP7_75t_R g6601 ( 
.A(n_5837),
.Y(n_6601)
);

NAND2xp5_ASAP7_75t_L g6602 ( 
.A(n_5913),
.B(n_3283),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6082),
.Y(n_6603)
);

NAND2xp5_ASAP7_75t_L g6604 ( 
.A(n_6208),
.B(n_3285),
.Y(n_6604)
);

BUFx3_ASAP7_75t_L g6605 ( 
.A(n_6240),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6083),
.Y(n_6606)
);

BUFx6f_ASAP7_75t_L g6607 ( 
.A(n_6113),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6094),
.Y(n_6608)
);

INVx4_ASAP7_75t_L g6609 ( 
.A(n_6335),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_SL g6610 ( 
.A(n_6146),
.B(n_3287),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_6100),
.Y(n_6611)
);

NAND2xp5_ASAP7_75t_L g6612 ( 
.A(n_6072),
.B(n_3288),
.Y(n_6612)
);

NAND2xp5_ASAP7_75t_L g6613 ( 
.A(n_6295),
.B(n_3289),
.Y(n_6613)
);

NOR2xp33_ASAP7_75t_L g6614 ( 
.A(n_6260),
.B(n_3291),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6103),
.Y(n_6615)
);

BUFx3_ASAP7_75t_L g6616 ( 
.A(n_5891),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6104),
.Y(n_6617)
);

INVx2_ASAP7_75t_L g6618 ( 
.A(n_6107),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_6110),
.Y(n_6619)
);

NOR2xp33_ASAP7_75t_L g6620 ( 
.A(n_5950),
.B(n_3292),
.Y(n_6620)
);

INVx5_ASAP7_75t_L g6621 ( 
.A(n_6113),
.Y(n_6621)
);

AND2x6_ASAP7_75t_L g6622 ( 
.A(n_6262),
.B(n_3566),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6117),
.Y(n_6623)
);

NOR3xp33_ASAP7_75t_L g6624 ( 
.A(n_6256),
.B(n_6358),
.C(n_6347),
.Y(n_6624)
);

AND2x6_ASAP7_75t_L g6625 ( 
.A(n_6275),
.B(n_3581),
.Y(n_6625)
);

NAND2xp5_ASAP7_75t_SL g6626 ( 
.A(n_6154),
.B(n_3294),
.Y(n_6626)
);

NAND2xp5_ASAP7_75t_SL g6627 ( 
.A(n_5952),
.B(n_3296),
.Y(n_6627)
);

NAND2xp5_ASAP7_75t_L g6628 ( 
.A(n_6126),
.B(n_3297),
.Y(n_6628)
);

INVx3_ASAP7_75t_L g6629 ( 
.A(n_6203),
.Y(n_6629)
);

AOI22xp5_ASAP7_75t_L g6630 ( 
.A1(n_6343),
.A2(n_3301),
.B1(n_3303),
.B2(n_3299),
.Y(n_6630)
);

AND3x2_ASAP7_75t_L g6631 ( 
.A(n_5904),
.B(n_5944),
.C(n_5906),
.Y(n_6631)
);

AND2x4_ASAP7_75t_L g6632 ( 
.A(n_6258),
.B(n_3597),
.Y(n_6632)
);

BUFx6f_ASAP7_75t_L g6633 ( 
.A(n_6203),
.Y(n_6633)
);

NOR2xp33_ASAP7_75t_L g6634 ( 
.A(n_5958),
.B(n_3304),
.Y(n_6634)
);

INVx3_ASAP7_75t_L g6635 ( 
.A(n_6203),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6131),
.Y(n_6636)
);

BUFx3_ASAP7_75t_L g6637 ( 
.A(n_5894),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6141),
.Y(n_6638)
);

NAND2xp33_ASAP7_75t_L g6639 ( 
.A(n_5985),
.B(n_5986),
.Y(n_6639)
);

BUFx10_ASAP7_75t_L g6640 ( 
.A(n_5838),
.Y(n_6640)
);

NAND2xp5_ASAP7_75t_L g6641 ( 
.A(n_6152),
.B(n_3306),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6159),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6162),
.Y(n_6643)
);

AND2x2_ASAP7_75t_L g6644 ( 
.A(n_5825),
.B(n_3313),
.Y(n_6644)
);

CKINVDCx5p33_ASAP7_75t_R g6645 ( 
.A(n_5841),
.Y(n_6645)
);

BUFx6f_ASAP7_75t_L g6646 ( 
.A(n_6284),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6206),
.Y(n_6647)
);

AND2x2_ASAP7_75t_L g6648 ( 
.A(n_6222),
.B(n_3315),
.Y(n_6648)
);

AOI22xp33_ASAP7_75t_L g6649 ( 
.A1(n_6300),
.A2(n_3601),
.B1(n_3602),
.B2(n_3598),
.Y(n_6649)
);

BUFx4f_ASAP7_75t_L g6650 ( 
.A(n_6246),
.Y(n_6650)
);

INVx5_ASAP7_75t_L g6651 ( 
.A(n_6122),
.Y(n_6651)
);

AND2x2_ASAP7_75t_SL g6652 ( 
.A(n_6184),
.B(n_3605),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_L g6653 ( 
.A(n_5945),
.B(n_6026),
.Y(n_6653)
);

NOR2xp33_ASAP7_75t_L g6654 ( 
.A(n_5966),
.B(n_3325),
.Y(n_6654)
);

BUFx3_ASAP7_75t_L g6655 ( 
.A(n_6245),
.Y(n_6655)
);

NAND2xp5_ASAP7_75t_L g6656 ( 
.A(n_6307),
.B(n_3327),
.Y(n_6656)
);

NAND2xp33_ASAP7_75t_L g6657 ( 
.A(n_5987),
.B(n_3328),
.Y(n_6657)
);

NOR2x1p5_ASAP7_75t_L g6658 ( 
.A(n_5849),
.B(n_3329),
.Y(n_6658)
);

BUFx6f_ASAP7_75t_L g6659 ( 
.A(n_6284),
.Y(n_6659)
);

BUFx2_ASAP7_75t_L g6660 ( 
.A(n_6028),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6011),
.B(n_3334),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_SL g6662 ( 
.A(n_5968),
.B(n_3335),
.Y(n_6662)
);

AND2x2_ASAP7_75t_L g6663 ( 
.A(n_5927),
.B(n_3337),
.Y(n_6663)
);

INVx4_ASAP7_75t_L g6664 ( 
.A(n_5850),
.Y(n_6664)
);

AND2x6_ASAP7_75t_L g6665 ( 
.A(n_6282),
.B(n_3606),
.Y(n_6665)
);

INVx4_ASAP7_75t_SL g6666 ( 
.A(n_6302),
.Y(n_6666)
);

AND2x2_ASAP7_75t_L g6667 ( 
.A(n_6223),
.B(n_3339),
.Y(n_6667)
);

AND2x2_ASAP7_75t_L g6668 ( 
.A(n_6339),
.B(n_6346),
.Y(n_6668)
);

BUFx6f_ASAP7_75t_L g6669 ( 
.A(n_6284),
.Y(n_6669)
);

NAND2xp5_ASAP7_75t_L g6670 ( 
.A(n_6317),
.B(n_3340),
.Y(n_6670)
);

INVx5_ASAP7_75t_L g6671 ( 
.A(n_6122),
.Y(n_6671)
);

BUFx3_ASAP7_75t_L g6672 ( 
.A(n_5932),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6211),
.Y(n_6673)
);

NOR2x1p5_ASAP7_75t_L g6674 ( 
.A(n_5853),
.B(n_3343),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_SL g6675 ( 
.A(n_5948),
.B(n_3344),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_L g6676 ( 
.A(n_6318),
.B(n_3348),
.Y(n_6676)
);

NAND2xp5_ASAP7_75t_SL g6677 ( 
.A(n_6012),
.B(n_3351),
.Y(n_6677)
);

OAI22xp33_ASAP7_75t_L g6678 ( 
.A1(n_6250),
.A2(n_3358),
.B1(n_3363),
.B2(n_3352),
.Y(n_6678)
);

INVx3_ASAP7_75t_L g6679 ( 
.A(n_5946),
.Y(n_6679)
);

NOR2xp33_ASAP7_75t_L g6680 ( 
.A(n_6166),
.B(n_3366),
.Y(n_6680)
);

INVxp33_ASAP7_75t_L g6681 ( 
.A(n_6063),
.Y(n_6681)
);

INVx4_ASAP7_75t_L g6682 ( 
.A(n_5857),
.Y(n_6682)
);

INVx4_ASAP7_75t_L g6683 ( 
.A(n_5858),
.Y(n_6683)
);

BUFx6f_ASAP7_75t_L g6684 ( 
.A(n_6136),
.Y(n_6684)
);

AND2x6_ASAP7_75t_L g6685 ( 
.A(n_6291),
.B(n_3609),
.Y(n_6685)
);

INVx3_ASAP7_75t_L g6686 ( 
.A(n_5946),
.Y(n_6686)
);

NOR2xp33_ASAP7_75t_L g6687 ( 
.A(n_6168),
.B(n_3368),
.Y(n_6687)
);

INVx5_ASAP7_75t_L g6688 ( 
.A(n_6136),
.Y(n_6688)
);

NAND2xp5_ASAP7_75t_L g6689 ( 
.A(n_6326),
.B(n_3369),
.Y(n_6689)
);

INVx3_ASAP7_75t_L g6690 ( 
.A(n_6304),
.Y(n_6690)
);

BUFx6f_ASAP7_75t_L g6691 ( 
.A(n_6336),
.Y(n_6691)
);

INVxp67_ASAP7_75t_SL g6692 ( 
.A(n_5903),
.Y(n_6692)
);

AND2x6_ASAP7_75t_L g6693 ( 
.A(n_6292),
.B(n_3610),
.Y(n_6693)
);

BUFx6f_ASAP7_75t_L g6694 ( 
.A(n_6338),
.Y(n_6694)
);

INVx1_ASAP7_75t_SL g6695 ( 
.A(n_5976),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6216),
.Y(n_6696)
);

NAND2xp5_ASAP7_75t_SL g6697 ( 
.A(n_5988),
.B(n_3370),
.Y(n_6697)
);

AND2x2_ASAP7_75t_L g6698 ( 
.A(n_6172),
.B(n_3372),
.Y(n_6698)
);

AOI22xp33_ASAP7_75t_L g6699 ( 
.A1(n_6246),
.A2(n_3617),
.B1(n_3625),
.B2(n_3614),
.Y(n_6699)
);

NAND2xp5_ASAP7_75t_SL g6700 ( 
.A(n_6009),
.B(n_3373),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_5979),
.Y(n_6701)
);

NOR2xp33_ASAP7_75t_L g6702 ( 
.A(n_6220),
.B(n_3374),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6217),
.Y(n_6703)
);

INVx1_ASAP7_75t_L g6704 ( 
.A(n_6226),
.Y(n_6704)
);

INVx1_ASAP7_75t_SL g6705 ( 
.A(n_5977),
.Y(n_6705)
);

INVx4_ASAP7_75t_L g6706 ( 
.A(n_5859),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6239),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_5999),
.Y(n_6708)
);

CKINVDCx5p33_ASAP7_75t_R g6709 ( 
.A(n_5842),
.Y(n_6709)
);

AOI22xp5_ASAP7_75t_L g6710 ( 
.A1(n_6266),
.A2(n_3382),
.B1(n_3383),
.B2(n_3381),
.Y(n_6710)
);

BUFx3_ASAP7_75t_L g6711 ( 
.A(n_5934),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6243),
.Y(n_6712)
);

AND2x2_ASAP7_75t_L g6713 ( 
.A(n_6180),
.B(n_3384),
.Y(n_6713)
);

NAND2xp5_ASAP7_75t_L g6714 ( 
.A(n_6327),
.B(n_3385),
.Y(n_6714)
);

INVx4_ASAP7_75t_L g6715 ( 
.A(n_5870),
.Y(n_6715)
);

BUFx3_ASAP7_75t_L g6716 ( 
.A(n_5877),
.Y(n_6716)
);

AOI22xp5_ASAP7_75t_L g6717 ( 
.A1(n_6246),
.A2(n_3390),
.B1(n_3391),
.B2(n_3388),
.Y(n_6717)
);

INVx4_ASAP7_75t_L g6718 ( 
.A(n_5871),
.Y(n_6718)
);

AND2x2_ASAP7_75t_L g6719 ( 
.A(n_6182),
.B(n_3392),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6247),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_6000),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_SL g6722 ( 
.A(n_5974),
.B(n_3393),
.Y(n_6722)
);

INVx4_ASAP7_75t_L g6723 ( 
.A(n_5873),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6261),
.Y(n_6724)
);

AND3x4_ASAP7_75t_L g6725 ( 
.A(n_6035),
.B(n_3190),
.C(n_3012),
.Y(n_6725)
);

BUFx3_ASAP7_75t_L g6726 ( 
.A(n_5887),
.Y(n_6726)
);

OR2x2_ASAP7_75t_SL g6727 ( 
.A(n_6214),
.B(n_3635),
.Y(n_6727)
);

AND2x6_ASAP7_75t_L g6728 ( 
.A(n_6297),
.B(n_6329),
.Y(n_6728)
);

AO22x2_ASAP7_75t_L g6729 ( 
.A1(n_6109),
.A2(n_3642),
.B1(n_3646),
.B2(n_3640),
.Y(n_6729)
);

INVx5_ASAP7_75t_L g6730 ( 
.A(n_6338),
.Y(n_6730)
);

INVx4_ASAP7_75t_L g6731 ( 
.A(n_5874),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6014),
.Y(n_6732)
);

INVx4_ASAP7_75t_L g6733 ( 
.A(n_5881),
.Y(n_6733)
);

INVx6_ASAP7_75t_L g6734 ( 
.A(n_6341),
.Y(n_6734)
);

NAND2xp5_ASAP7_75t_L g6735 ( 
.A(n_6333),
.B(n_3394),
.Y(n_6735)
);

CKINVDCx20_ASAP7_75t_R g6736 ( 
.A(n_5846),
.Y(n_6736)
);

NAND2xp5_ASAP7_75t_L g6737 ( 
.A(n_6334),
.B(n_6015),
.Y(n_6737)
);

NOR2xp33_ASAP7_75t_L g6738 ( 
.A(n_6224),
.B(n_3398),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_L g6739 ( 
.A(n_6017),
.B(n_3400),
.Y(n_6739)
);

NAND2xp5_ASAP7_75t_SL g6740 ( 
.A(n_5991),
.B(n_3403),
.Y(n_6740)
);

INVx1_ASAP7_75t_SL g6741 ( 
.A(n_5981),
.Y(n_6741)
);

BUFx6f_ASAP7_75t_SL g6742 ( 
.A(n_6246),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_SL g6743 ( 
.A(n_5992),
.B(n_3404),
.Y(n_6743)
);

INVx4_ASAP7_75t_L g6744 ( 
.A(n_5907),
.Y(n_6744)
);

INVxp33_ASAP7_75t_SL g6745 ( 
.A(n_5845),
.Y(n_6745)
);

INVx2_ASAP7_75t_SL g6746 ( 
.A(n_6283),
.Y(n_6746)
);

NOR2x1p5_ASAP7_75t_L g6747 ( 
.A(n_5896),
.B(n_3411),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6027),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6342),
.B(n_3413),
.Y(n_6749)
);

AND2x4_ASAP7_75t_L g6750 ( 
.A(n_6093),
.B(n_3647),
.Y(n_6750)
);

INVx2_ASAP7_75t_L g6751 ( 
.A(n_6066),
.Y(n_6751)
);

BUFx8_ASAP7_75t_SL g6752 ( 
.A(n_5848),
.Y(n_6752)
);

INVx3_ASAP7_75t_L g6753 ( 
.A(n_6304),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6069),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6075),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6076),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_SL g6757 ( 
.A(n_5993),
.B(n_3414),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6079),
.Y(n_6758)
);

BUFx6f_ASAP7_75t_L g6759 ( 
.A(n_6197),
.Y(n_6759)
);

NAND2xp5_ASAP7_75t_L g6760 ( 
.A(n_6086),
.B(n_6091),
.Y(n_6760)
);

NAND2xp5_ASAP7_75t_L g6761 ( 
.A(n_6092),
.B(n_3416),
.Y(n_6761)
);

NOR2xp33_ASAP7_75t_L g6762 ( 
.A(n_6225),
.B(n_3417),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6112),
.B(n_3418),
.Y(n_6763)
);

INVx2_ASAP7_75t_SL g6764 ( 
.A(n_6287),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6121),
.Y(n_6765)
);

AND2x2_ASAP7_75t_L g6766 ( 
.A(n_6345),
.B(n_3419),
.Y(n_6766)
);

INVx1_ASAP7_75t_SL g6767 ( 
.A(n_6289),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6132),
.Y(n_6768)
);

NOR2x1p5_ASAP7_75t_L g6769 ( 
.A(n_5885),
.B(n_3423),
.Y(n_6769)
);

BUFx8_ASAP7_75t_SL g6770 ( 
.A(n_5851),
.Y(n_6770)
);

OR2x2_ASAP7_75t_L g6771 ( 
.A(n_6234),
.B(n_3425),
.Y(n_6771)
);

INVx3_ASAP7_75t_L g6772 ( 
.A(n_6360),
.Y(n_6772)
);

INVxp67_ASAP7_75t_L g6773 ( 
.A(n_6288),
.Y(n_6773)
);

CKINVDCx16_ASAP7_75t_R g6774 ( 
.A(n_5860),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_6147),
.B(n_3429),
.Y(n_6775)
);

NOR2xp33_ASAP7_75t_L g6776 ( 
.A(n_6227),
.B(n_3432),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6155),
.Y(n_6777)
);

NAND2xp5_ASAP7_75t_SL g6778 ( 
.A(n_5997),
.B(n_3434),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6157),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6176),
.Y(n_6780)
);

CKINVDCx5p33_ASAP7_75t_R g6781 ( 
.A(n_5847),
.Y(n_6781)
);

AOI22xp33_ASAP7_75t_L g6782 ( 
.A1(n_6302),
.A2(n_3653),
.B1(n_3654),
.B2(n_3648),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6200),
.Y(n_6783)
);

AO22x2_ASAP7_75t_L g6784 ( 
.A1(n_6139),
.A2(n_3659),
.B1(n_3665),
.B2(n_3656),
.Y(n_6784)
);

NOR2xp33_ASAP7_75t_L g6785 ( 
.A(n_6229),
.B(n_3436),
.Y(n_6785)
);

NAND2xp5_ASAP7_75t_L g6786 ( 
.A(n_6202),
.B(n_3438),
.Y(n_6786)
);

NAND2xp33_ASAP7_75t_L g6787 ( 
.A(n_6130),
.B(n_3440),
.Y(n_6787)
);

NOR2xp33_ASAP7_75t_L g6788 ( 
.A(n_6231),
.B(n_3447),
.Y(n_6788)
);

NOR2xp33_ASAP7_75t_L g6789 ( 
.A(n_6219),
.B(n_3449),
.Y(n_6789)
);

INVx4_ASAP7_75t_L g6790 ( 
.A(n_5890),
.Y(n_6790)
);

AND2x6_ASAP7_75t_L g6791 ( 
.A(n_6265),
.B(n_3667),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_6241),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_SL g6793 ( 
.A(n_5998),
.B(n_6001),
.Y(n_6793)
);

NOR2xp33_ASAP7_75t_L g6794 ( 
.A(n_6099),
.B(n_3450),
.Y(n_6794)
);

BUFx3_ASAP7_75t_L g6795 ( 
.A(n_5893),
.Y(n_6795)
);

OAI22xp33_ASAP7_75t_L g6796 ( 
.A1(n_6190),
.A2(n_3456),
.B1(n_3463),
.B2(n_3454),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_L g6797 ( 
.A(n_6248),
.B(n_6253),
.Y(n_6797)
);

NOR2xp33_ASAP7_75t_L g6798 ( 
.A(n_6105),
.B(n_3464),
.Y(n_6798)
);

INVx4_ASAP7_75t_L g6799 ( 
.A(n_5929),
.Y(n_6799)
);

INVx2_ASAP7_75t_L g6800 ( 
.A(n_5903),
.Y(n_6800)
);

NAND2xp5_ASAP7_75t_SL g6801 ( 
.A(n_6002),
.B(n_3466),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6270),
.Y(n_6802)
);

INVx1_ASAP7_75t_SL g6803 ( 
.A(n_6293),
.Y(n_6803)
);

BUFx6f_ASAP7_75t_L g6804 ( 
.A(n_6363),
.Y(n_6804)
);

INVx2_ASAP7_75t_L g6805 ( 
.A(n_5911),
.Y(n_6805)
);

NAND2xp5_ASAP7_75t_L g6806 ( 
.A(n_6236),
.B(n_3471),
.Y(n_6806)
);

NAND2xp33_ASAP7_75t_L g6807 ( 
.A(n_6167),
.B(n_6195),
.Y(n_6807)
);

NOR2xp33_ASAP7_75t_L g6808 ( 
.A(n_6005),
.B(n_3473),
.Y(n_6808)
);

NAND2xp5_ASAP7_75t_L g6809 ( 
.A(n_6281),
.B(n_3477),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_6277),
.Y(n_6810)
);

NAND2xp5_ASAP7_75t_SL g6811 ( 
.A(n_5984),
.B(n_3481),
.Y(n_6811)
);

NAND2xp5_ASAP7_75t_L g6812 ( 
.A(n_6148),
.B(n_3484),
.Y(n_6812)
);

NAND2xp5_ASAP7_75t_L g6813 ( 
.A(n_5911),
.B(n_6033),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6316),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6033),
.Y(n_6815)
);

AND2x6_ASAP7_75t_L g6816 ( 
.A(n_6323),
.B(n_3674),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6067),
.B(n_3491),
.Y(n_6817)
);

AND2x4_ASAP7_75t_L g6818 ( 
.A(n_6299),
.B(n_3682),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_SL g6819 ( 
.A(n_6007),
.B(n_3492),
.Y(n_6819)
);

NAND2xp5_ASAP7_75t_L g6820 ( 
.A(n_6067),
.B(n_3493),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_SL g6821 ( 
.A(n_6357),
.B(n_3496),
.Y(n_6821)
);

BUFx3_ASAP7_75t_L g6822 ( 
.A(n_5905),
.Y(n_6822)
);

BUFx2_ASAP7_75t_L g6823 ( 
.A(n_5910),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6073),
.Y(n_6824)
);

INVx3_ASAP7_75t_L g6825 ( 
.A(n_6364),
.Y(n_6825)
);

AND2x2_ASAP7_75t_L g6826 ( 
.A(n_5909),
.B(n_3502),
.Y(n_6826)
);

INVxp67_ASAP7_75t_SL g6827 ( 
.A(n_6073),
.Y(n_6827)
);

BUFx10_ASAP7_75t_L g6828 ( 
.A(n_5888),
.Y(n_6828)
);

INVx3_ASAP7_75t_L g6829 ( 
.A(n_6078),
.Y(n_6829)
);

AOI22xp33_ASAP7_75t_L g6830 ( 
.A1(n_6302),
.A2(n_3693),
.B1(n_3696),
.B2(n_3684),
.Y(n_6830)
);

INVx5_ASAP7_75t_L g6831 ( 
.A(n_6302),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_6078),
.B(n_3505),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6090),
.B(n_3506),
.Y(n_6833)
);

OAI22xp33_ASAP7_75t_L g6834 ( 
.A1(n_6242),
.A2(n_3512),
.B1(n_3516),
.B2(n_3511),
.Y(n_6834)
);

INVx6_ASAP7_75t_L g6835 ( 
.A(n_6341),
.Y(n_6835)
);

NOR2xp33_ASAP7_75t_L g6836 ( 
.A(n_6120),
.B(n_6019),
.Y(n_6836)
);

INVx3_ASAP7_75t_L g6837 ( 
.A(n_6090),
.Y(n_6837)
);

NAND2x1p5_ASAP7_75t_L g6838 ( 
.A(n_6235),
.B(n_3698),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6235),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6255),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6255),
.B(n_6273),
.Y(n_6841)
);

INVx3_ASAP7_75t_L g6842 ( 
.A(n_6273),
.Y(n_6842)
);

AND2x6_ASAP7_75t_L g6843 ( 
.A(n_6328),
.B(n_3703),
.Y(n_6843)
);

INVx4_ASAP7_75t_L g6844 ( 
.A(n_5935),
.Y(n_6844)
);

INVxp33_ASAP7_75t_L g6845 ( 
.A(n_6095),
.Y(n_6845)
);

INVx3_ASAP7_75t_L g6846 ( 
.A(n_6274),
.Y(n_6846)
);

AOI22xp33_ASAP7_75t_L g6847 ( 
.A1(n_5947),
.A2(n_3717),
.B1(n_3718),
.B2(n_3712),
.Y(n_6847)
);

INVx2_ASAP7_75t_SL g6848 ( 
.A(n_6296),
.Y(n_6848)
);

NAND2xp5_ASAP7_75t_L g6849 ( 
.A(n_6274),
.B(n_6290),
.Y(n_6849)
);

BUFx10_ASAP7_75t_L g6850 ( 
.A(n_5862),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6290),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_5868),
.B(n_3517),
.Y(n_6852)
);

NOR2xp33_ASAP7_75t_L g6853 ( 
.A(n_6023),
.B(n_3518),
.Y(n_6853)
);

INVx3_ASAP7_75t_L g6854 ( 
.A(n_6370),
.Y(n_6854)
);

INVx2_ASAP7_75t_L g6855 ( 
.A(n_5947),
.Y(n_6855)
);

INVx2_ASAP7_75t_L g6856 ( 
.A(n_6340),
.Y(n_6856)
);

INVx2_ASAP7_75t_L g6857 ( 
.A(n_6340),
.Y(n_6857)
);

AND2x6_ASAP7_75t_L g6858 ( 
.A(n_5972),
.B(n_3727),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6144),
.B(n_3520),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_L g6860 ( 
.A(n_6331),
.B(n_3524),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6306),
.Y(n_6861)
);

INVx2_ASAP7_75t_SL g6862 ( 
.A(n_6221),
.Y(n_6862)
);

BUFx2_ASAP7_75t_L g6863 ( 
.A(n_5914),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6319),
.Y(n_6864)
);

CKINVDCx16_ASAP7_75t_R g6865 ( 
.A(n_5861),
.Y(n_6865)
);

BUFx10_ASAP7_75t_L g6866 ( 
.A(n_5863),
.Y(n_6866)
);

INVx2_ASAP7_75t_L g6867 ( 
.A(n_6313),
.Y(n_6867)
);

INVx2_ASAP7_75t_SL g6868 ( 
.A(n_6303),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_6192),
.B(n_3529),
.Y(n_6869)
);

BUFx3_ASAP7_75t_L g6870 ( 
.A(n_5967),
.Y(n_6870)
);

AOI22xp33_ASAP7_75t_L g6871 ( 
.A1(n_6188),
.A2(n_3738),
.B1(n_3739),
.B2(n_3734),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6230),
.Y(n_6872)
);

INVx1_ASAP7_75t_SL g6873 ( 
.A(n_5942),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6353),
.Y(n_6874)
);

INVx4_ASAP7_75t_SL g6875 ( 
.A(n_5975),
.Y(n_6875)
);

NAND2x1p5_ASAP7_75t_L g6876 ( 
.A(n_6170),
.B(n_3741),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_SL g6877 ( 
.A(n_6194),
.B(n_3530),
.Y(n_6877)
);

BUFx10_ASAP7_75t_L g6878 ( 
.A(n_6160),
.Y(n_6878)
);

INVx2_ASAP7_75t_SL g6879 ( 
.A(n_6322),
.Y(n_6879)
);

INVx5_ASAP7_75t_L g6880 ( 
.A(n_6359),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_SL g6881 ( 
.A(n_5930),
.B(n_3537),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6356),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_5925),
.Y(n_6883)
);

INVx2_ASAP7_75t_L g6884 ( 
.A(n_6031),
.Y(n_6884)
);

NOR2x1_ASAP7_75t_L g6885 ( 
.A(n_6179),
.B(n_3743),
.Y(n_6885)
);

INVx4_ASAP7_75t_L g6886 ( 
.A(n_5928),
.Y(n_6886)
);

NOR2xp33_ASAP7_75t_L g6887 ( 
.A(n_6169),
.B(n_3542),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6034),
.Y(n_6888)
);

NAND2xp5_ASAP7_75t_L g6889 ( 
.A(n_6199),
.B(n_6165),
.Y(n_6889)
);

INVx2_ASAP7_75t_L g6890 ( 
.A(n_6038),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6041),
.Y(n_6891)
);

NAND2xp5_ASAP7_75t_L g6892 ( 
.A(n_6022),
.B(n_3544),
.Y(n_6892)
);

AOI22xp5_ASAP7_75t_L g6893 ( 
.A1(n_6276),
.A2(n_3546),
.B1(n_3548),
.B2(n_3545),
.Y(n_6893)
);

NAND2xp5_ASAP7_75t_SL g6894 ( 
.A(n_6118),
.B(n_3549),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6048),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6198),
.B(n_3552),
.Y(n_6896)
);

INVxp67_ASAP7_75t_SL g6897 ( 
.A(n_6185),
.Y(n_6897)
);

NAND2xp5_ASAP7_75t_SL g6898 ( 
.A(n_6119),
.B(n_3553),
.Y(n_6898)
);

BUFx6f_ASAP7_75t_L g6899 ( 
.A(n_5854),
.Y(n_6899)
);

NOR2xp33_ASAP7_75t_L g6900 ( 
.A(n_6053),
.B(n_3555),
.Y(n_6900)
);

AND2x6_ASAP7_75t_L g6901 ( 
.A(n_6324),
.B(n_3744),
.Y(n_6901)
);

OAI21xp33_ASAP7_75t_SL g6902 ( 
.A1(n_6244),
.A2(n_3754),
.B(n_3750),
.Y(n_6902)
);

INVx4_ASAP7_75t_L g6903 ( 
.A(n_5955),
.Y(n_6903)
);

INVxp67_ASAP7_75t_SL g6904 ( 
.A(n_6204),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6054),
.Y(n_6905)
);

AND2x2_ASAP7_75t_SL g6906 ( 
.A(n_6036),
.B(n_3758),
.Y(n_6906)
);

NAND2xp5_ASAP7_75t_SL g6907 ( 
.A(n_5899),
.B(n_3557),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6055),
.Y(n_6908)
);

NAND2xp5_ASAP7_75t_L g6909 ( 
.A(n_6365),
.B(n_3558),
.Y(n_6909)
);

NAND2xp5_ASAP7_75t_L g6910 ( 
.A(n_6268),
.B(n_3559),
.Y(n_6910)
);

NOR2xp33_ASAP7_75t_L g6911 ( 
.A(n_6056),
.B(n_3564),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_6133),
.B(n_3565),
.Y(n_6912)
);

AOI22xp33_ASAP7_75t_L g6913 ( 
.A1(n_6114),
.A2(n_3761),
.B1(n_3762),
.B2(n_3760),
.Y(n_6913)
);

AOI22xp5_ASAP7_75t_L g6914 ( 
.A1(n_6251),
.A2(n_3569),
.B1(n_3570),
.B2(n_3568),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6205),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6209),
.Y(n_6916)
);

NAND2xp5_ASAP7_75t_SL g6917 ( 
.A(n_6134),
.B(n_3571),
.Y(n_6917)
);

INVx2_ASAP7_75t_SL g6918 ( 
.A(n_6212),
.Y(n_6918)
);

INVx3_ASAP7_75t_L g6919 ( 
.A(n_5938),
.Y(n_6919)
);

NAND2xp5_ASAP7_75t_L g6920 ( 
.A(n_6071),
.B(n_3574),
.Y(n_6920)
);

INVx2_ASAP7_75t_SL g6921 ( 
.A(n_6061),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_6252),
.Y(n_6922)
);

NAND2xp5_ASAP7_75t_L g6923 ( 
.A(n_6378),
.B(n_6074),
.Y(n_6923)
);

BUFx6f_ASAP7_75t_SL g6924 ( 
.A(n_6672),
.Y(n_6924)
);

NAND2xp5_ASAP7_75t_L g6925 ( 
.A(n_6381),
.B(n_6080),
.Y(n_6925)
);

NAND2xp5_ASAP7_75t_SL g6926 ( 
.A(n_6652),
.B(n_6138),
.Y(n_6926)
);

NAND2xp5_ASAP7_75t_SL g6927 ( 
.A(n_6399),
.B(n_6140),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_SL g6928 ( 
.A(n_6398),
.B(n_6084),
.Y(n_6928)
);

AND2x6_ASAP7_75t_SL g6929 ( 
.A(n_6571),
.B(n_5883),
.Y(n_6929)
);

NAND3xp33_ASAP7_75t_L g6930 ( 
.A(n_6680),
.B(n_6049),
.C(n_5954),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_6481),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6397),
.Y(n_6932)
);

NAND2xp5_ASAP7_75t_L g6933 ( 
.A(n_6388),
.B(n_6097),
.Y(n_6933)
);

OAI22xp5_ASAP7_75t_L g6934 ( 
.A1(n_6889),
.A2(n_6653),
.B1(n_6374),
.B2(n_6416),
.Y(n_6934)
);

INVx1_ASAP7_75t_L g6935 ( 
.A(n_6415),
.Y(n_6935)
);

NAND2xp5_ASAP7_75t_L g6936 ( 
.A(n_6392),
.B(n_6098),
.Y(n_6936)
);

INVx2_ASAP7_75t_L g6937 ( 
.A(n_6488),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6420),
.Y(n_6938)
);

NAND2xp5_ASAP7_75t_SL g6939 ( 
.A(n_6401),
.B(n_5939),
.Y(n_6939)
);

NAND2xp5_ASAP7_75t_L g6940 ( 
.A(n_6469),
.B(n_6215),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6477),
.B(n_6218),
.Y(n_6941)
);

INVx2_ASAP7_75t_L g6942 ( 
.A(n_6496),
.Y(n_6942)
);

NOR2xp33_ASAP7_75t_L g6943 ( 
.A(n_6702),
.B(n_5940),
.Y(n_6943)
);

INVxp67_ASAP7_75t_SL g6944 ( 
.A(n_6412),
.Y(n_6944)
);

NAND2xp5_ASAP7_75t_SL g6945 ( 
.A(n_6428),
.B(n_5969),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_SL g6946 ( 
.A(n_6546),
.B(n_5971),
.Y(n_6946)
);

NAND2xp5_ASAP7_75t_L g6947 ( 
.A(n_6478),
.B(n_6153),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_6485),
.B(n_6087),
.Y(n_6948)
);

NAND2xp5_ASAP7_75t_L g6949 ( 
.A(n_6405),
.B(n_6108),
.Y(n_6949)
);

NOR2xp33_ASAP7_75t_L g6950 ( 
.A(n_6789),
.B(n_6210),
.Y(n_6950)
);

BUFx6f_ASAP7_75t_SL g6951 ( 
.A(n_6711),
.Y(n_6951)
);

NAND2xp5_ASAP7_75t_L g6952 ( 
.A(n_6613),
.B(n_6115),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_6437),
.Y(n_6953)
);

CKINVDCx5p33_ASAP7_75t_R g6954 ( 
.A(n_6375),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6687),
.B(n_6040),
.Y(n_6955)
);

INVx2_ASAP7_75t_L g6956 ( 
.A(n_6507),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6604),
.B(n_6058),
.Y(n_6957)
);

NOR2xp33_ASAP7_75t_L g6958 ( 
.A(n_6738),
.B(n_5830),
.Y(n_6958)
);

INVx2_ASAP7_75t_L g6959 ( 
.A(n_6510),
.Y(n_6959)
);

NOR2xp33_ASAP7_75t_L g6960 ( 
.A(n_6762),
.B(n_6143),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6438),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_6517),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_6602),
.B(n_6442),
.Y(n_6963)
);

INVx2_ASAP7_75t_SL g6964 ( 
.A(n_6385),
.Y(n_6964)
);

NAND2xp33_ASAP7_75t_L g6965 ( 
.A(n_6430),
.B(n_6024),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6443),
.Y(n_6966)
);

OAI22xp33_ASAP7_75t_L g6967 ( 
.A1(n_6526),
.A2(n_6773),
.B1(n_6869),
.B2(n_6764),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6448),
.B(n_3575),
.Y(n_6968)
);

INVx2_ASAP7_75t_L g6969 ( 
.A(n_6530),
.Y(n_6969)
);

NOR2xp33_ASAP7_75t_L g6970 ( 
.A(n_6776),
.B(n_6123),
.Y(n_6970)
);

INVx2_ASAP7_75t_L g6971 ( 
.A(n_6547),
.Y(n_6971)
);

INVx2_ASAP7_75t_SL g6972 ( 
.A(n_6406),
.Y(n_6972)
);

OR2x6_ASAP7_75t_L g6973 ( 
.A(n_6479),
.B(n_5828),
.Y(n_6973)
);

INVx2_ASAP7_75t_SL g6974 ( 
.A(n_6427),
.Y(n_6974)
);

NAND2xp5_ASAP7_75t_L g6975 ( 
.A(n_6454),
.B(n_3576),
.Y(n_6975)
);

CKINVDCx14_ASAP7_75t_R g6976 ( 
.A(n_6736),
.Y(n_6976)
);

NAND2xp5_ASAP7_75t_L g6977 ( 
.A(n_6459),
.B(n_6463),
.Y(n_6977)
);

INVx4_ASAP7_75t_L g6978 ( 
.A(n_6494),
.Y(n_6978)
);

OR2x2_ASAP7_75t_L g6979 ( 
.A(n_6767),
.B(n_6013),
.Y(n_6979)
);

INVx4_ASAP7_75t_L g6980 ( 
.A(n_6494),
.Y(n_6980)
);

NAND3xp33_ASAP7_75t_L g6981 ( 
.A(n_6785),
.B(n_6125),
.C(n_6124),
.Y(n_6981)
);

INVx3_ASAP7_75t_L g6982 ( 
.A(n_6655),
.Y(n_6982)
);

INVx2_ASAP7_75t_L g6983 ( 
.A(n_6548),
.Y(n_6983)
);

INVxp67_ASAP7_75t_L g6984 ( 
.A(n_6543),
.Y(n_6984)
);

NAND2xp5_ASAP7_75t_L g6985 ( 
.A(n_6475),
.B(n_3578),
.Y(n_6985)
);

NAND2xp5_ASAP7_75t_L g6986 ( 
.A(n_6476),
.B(n_6486),
.Y(n_6986)
);

NAND2xp5_ASAP7_75t_L g6987 ( 
.A(n_6489),
.B(n_3580),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6490),
.B(n_3582),
.Y(n_6988)
);

NAND2xp33_ASAP7_75t_L g6989 ( 
.A(n_6440),
.B(n_6059),
.Y(n_6989)
);

NAND2xp5_ASAP7_75t_L g6990 ( 
.A(n_6499),
.B(n_3587),
.Y(n_6990)
);

INVx1_ASAP7_75t_L g6991 ( 
.A(n_6501),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6506),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6538),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6541),
.B(n_3590),
.Y(n_6994)
);

NAND2xp5_ASAP7_75t_L g6995 ( 
.A(n_6554),
.B(n_3591),
.Y(n_6995)
);

NAND2xp5_ASAP7_75t_L g6996 ( 
.A(n_6556),
.B(n_3592),
.Y(n_6996)
);

NOR2xp33_ASAP7_75t_L g6997 ( 
.A(n_6788),
.B(n_6161),
.Y(n_6997)
);

AND2x2_ASAP7_75t_L g6998 ( 
.A(n_6794),
.B(n_6164),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6566),
.B(n_6576),
.Y(n_6999)
);

NAND2xp5_ASAP7_75t_L g7000 ( 
.A(n_6577),
.B(n_3595),
.Y(n_7000)
);

O2A1O1Ixp33_ASAP7_75t_L g7001 ( 
.A1(n_6809),
.A2(n_3766),
.B(n_3768),
.C(n_3763),
.Y(n_7001)
);

NAND2xp5_ASAP7_75t_L g7002 ( 
.A(n_6582),
.B(n_3596),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_L g7003 ( 
.A(n_6591),
.B(n_3604),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6551),
.Y(n_7004)
);

NAND2xp5_ASAP7_75t_SL g7005 ( 
.A(n_6583),
.B(n_6062),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_SL g7006 ( 
.A(n_6836),
.B(n_6101),
.Y(n_7006)
);

NAND2xp5_ASAP7_75t_L g7007 ( 
.A(n_6595),
.B(n_3607),
.Y(n_7007)
);

INVx2_ASAP7_75t_L g7008 ( 
.A(n_6569),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_6597),
.B(n_3608),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6603),
.Y(n_7010)
);

NAND2xp5_ASAP7_75t_SL g7011 ( 
.A(n_6746),
.B(n_6142),
.Y(n_7011)
);

NAND2xp5_ASAP7_75t_SL g7012 ( 
.A(n_6848),
.B(n_6016),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6606),
.B(n_3613),
.Y(n_7013)
);

INVxp67_ASAP7_75t_L g7014 ( 
.A(n_6505),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_6608),
.B(n_3616),
.Y(n_7015)
);

NOR2xp67_ASAP7_75t_L g7016 ( 
.A(n_6664),
.B(n_3619),
.Y(n_7016)
);

NOR2xp33_ASAP7_75t_L g7017 ( 
.A(n_6798),
.B(n_3620),
.Y(n_7017)
);

INVx2_ASAP7_75t_SL g7018 ( 
.A(n_6497),
.Y(n_7018)
);

AND2x2_ASAP7_75t_L g7019 ( 
.A(n_6550),
.B(n_3621),
.Y(n_7019)
);

AND2x2_ASAP7_75t_L g7020 ( 
.A(n_6529),
.B(n_3623),
.Y(n_7020)
);

NAND2xp5_ASAP7_75t_L g7021 ( 
.A(n_6611),
.B(n_3629),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_L g7022 ( 
.A(n_6615),
.B(n_3631),
.Y(n_7022)
);

NAND2xp5_ASAP7_75t_L g7023 ( 
.A(n_6617),
.B(n_3634),
.Y(n_7023)
);

NAND2xp5_ASAP7_75t_SL g7024 ( 
.A(n_6884),
.B(n_3638),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6619),
.Y(n_7025)
);

NAND2xp5_ASAP7_75t_L g7026 ( 
.A(n_6636),
.B(n_3639),
.Y(n_7026)
);

O2A1O1Ixp33_ASAP7_75t_L g7027 ( 
.A1(n_6426),
.A2(n_3791),
.B(n_3795),
.C(n_3776),
.Y(n_7027)
);

NOR2xp67_ASAP7_75t_L g7028 ( 
.A(n_6682),
.B(n_3641),
.Y(n_7028)
);

NAND2xp5_ASAP7_75t_SL g7029 ( 
.A(n_6888),
.B(n_3652),
.Y(n_7029)
);

NAND2xp5_ASAP7_75t_L g7030 ( 
.A(n_6638),
.B(n_3655),
.Y(n_7030)
);

INVx2_ASAP7_75t_L g7031 ( 
.A(n_6575),
.Y(n_7031)
);

NOR2xp67_ASAP7_75t_L g7032 ( 
.A(n_6683),
.B(n_3657),
.Y(n_7032)
);

NOR2xp33_ASAP7_75t_L g7033 ( 
.A(n_6423),
.B(n_3658),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_6618),
.Y(n_7034)
);

INVx2_ASAP7_75t_L g7035 ( 
.A(n_6623),
.Y(n_7035)
);

NAND2xp5_ASAP7_75t_L g7036 ( 
.A(n_6642),
.B(n_3660),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6382),
.Y(n_7037)
);

INVx2_ASAP7_75t_SL g7038 ( 
.A(n_6497),
.Y(n_7038)
);

NOR2xp33_ASAP7_75t_L g7039 ( 
.A(n_6431),
.B(n_3662),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_SL g7040 ( 
.A(n_6890),
.B(n_3664),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6643),
.Y(n_7041)
);

NAND2xp5_ASAP7_75t_L g7042 ( 
.A(n_6812),
.B(n_3669),
.Y(n_7042)
);

AND2x2_ASAP7_75t_SL g7043 ( 
.A(n_6906),
.B(n_3797),
.Y(n_7043)
);

NOR3xp33_ASAP7_75t_L g7044 ( 
.A(n_6522),
.B(n_3673),
.C(n_3672),
.Y(n_7044)
);

XOR2xp5_ASAP7_75t_L g7045 ( 
.A(n_6592),
.B(n_3675),
.Y(n_7045)
);

NAND2xp5_ASAP7_75t_L g7046 ( 
.A(n_6387),
.B(n_3677),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_SL g7047 ( 
.A(n_6918),
.B(n_3678),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_6872),
.B(n_3679),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6647),
.Y(n_7049)
);

NAND2xp5_ASAP7_75t_L g7050 ( 
.A(n_6883),
.B(n_3686),
.Y(n_7050)
);

AOI22xp5_ASAP7_75t_L g7051 ( 
.A1(n_6882),
.A2(n_3688),
.B1(n_3691),
.B2(n_3687),
.Y(n_7051)
);

NAND2xp5_ASAP7_75t_L g7052 ( 
.A(n_6491),
.B(n_3694),
.Y(n_7052)
);

NAND2xp5_ASAP7_75t_SL g7053 ( 
.A(n_6921),
.B(n_3697),
.Y(n_7053)
);

NAND2xp5_ASAP7_75t_L g7054 ( 
.A(n_6673),
.B(n_3700),
.Y(n_7054)
);

NOR2xp33_ASAP7_75t_L g7055 ( 
.A(n_6585),
.B(n_3704),
.Y(n_7055)
);

NOR2x1p5_ASAP7_75t_L g7056 ( 
.A(n_6616),
.B(n_3706),
.Y(n_7056)
);

INVx2_ASAP7_75t_L g7057 ( 
.A(n_6384),
.Y(n_7057)
);

AND2x2_ASAP7_75t_L g7058 ( 
.A(n_6542),
.B(n_3707),
.Y(n_7058)
);

INVx2_ASAP7_75t_L g7059 ( 
.A(n_6394),
.Y(n_7059)
);

OR2x2_ASAP7_75t_L g7060 ( 
.A(n_6803),
.B(n_3708),
.Y(n_7060)
);

NAND2xp5_ASAP7_75t_L g7061 ( 
.A(n_6696),
.B(n_6703),
.Y(n_7061)
);

NAND2xp5_ASAP7_75t_L g7062 ( 
.A(n_6704),
.B(n_3711),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6707),
.B(n_3714),
.Y(n_7063)
);

INVx2_ASAP7_75t_SL g7064 ( 
.A(n_6516),
.Y(n_7064)
);

NAND2xp5_ASAP7_75t_L g7065 ( 
.A(n_6712),
.B(n_3715),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_L g7066 ( 
.A(n_6720),
.B(n_3719),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6724),
.B(n_3720),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6760),
.Y(n_7068)
);

NOR2xp33_ASAP7_75t_L g7069 ( 
.A(n_6593),
.B(n_3721),
.Y(n_7069)
);

AND2x2_ASAP7_75t_L g7070 ( 
.A(n_6544),
.B(n_3722),
.Y(n_7070)
);

INVxp67_ASAP7_75t_L g7071 ( 
.A(n_6483),
.Y(n_7071)
);

NAND2xp33_ASAP7_75t_L g7072 ( 
.A(n_6601),
.B(n_3723),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6797),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6732),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_SL g7075 ( 
.A(n_6461),
.B(n_3724),
.Y(n_7075)
);

NOR2xp33_ASAP7_75t_L g7076 ( 
.A(n_6396),
.B(n_3725),
.Y(n_7076)
);

AOI22xp33_ASAP7_75t_L g7077 ( 
.A1(n_6901),
.A2(n_3825),
.B1(n_3827),
.B2(n_3807),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6748),
.Y(n_7078)
);

NOR2xp33_ASAP7_75t_L g7079 ( 
.A(n_6451),
.B(n_3726),
.Y(n_7079)
);

NAND2xp5_ASAP7_75t_L g7080 ( 
.A(n_6901),
.B(n_3730),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6411),
.B(n_3733),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6644),
.B(n_3735),
.Y(n_7082)
);

NAND2xp5_ASAP7_75t_L g7083 ( 
.A(n_6892),
.B(n_3736),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6701),
.B(n_3737),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6758),
.Y(n_7085)
);

NOR2xp33_ASAP7_75t_L g7086 ( 
.A(n_6681),
.B(n_3740),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6765),
.Y(n_7087)
);

INVx2_ASAP7_75t_SL g7088 ( 
.A(n_6516),
.Y(n_7088)
);

INVx2_ASAP7_75t_SL g7089 ( 
.A(n_6621),
.Y(n_7089)
);

NAND2xp33_ASAP7_75t_L g7090 ( 
.A(n_6645),
.B(n_3742),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_SL g7091 ( 
.A(n_6891),
.B(n_3745),
.Y(n_7091)
);

HB1xp67_ASAP7_75t_L g7092 ( 
.A(n_6668),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6777),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_L g7094 ( 
.A(n_6708),
.B(n_3747),
.Y(n_7094)
);

INVxp67_ASAP7_75t_L g7095 ( 
.A(n_6393),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_6721),
.B(n_3748),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_L g7097 ( 
.A(n_6751),
.B(n_3749),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_L g7098 ( 
.A(n_6754),
.B(n_3752),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6779),
.Y(n_7099)
);

NAND2xp33_ASAP7_75t_L g7100 ( 
.A(n_6709),
.B(n_6791),
.Y(n_7100)
);

AND2x2_ASAP7_75t_L g7101 ( 
.A(n_6424),
.B(n_3756),
.Y(n_7101)
);

NOR2xp33_ASAP7_75t_L g7102 ( 
.A(n_6845),
.B(n_3757),
.Y(n_7102)
);

NOR2xp33_ASAP7_75t_R g7103 ( 
.A(n_6781),
.B(n_3759),
.Y(n_7103)
);

BUFx3_ASAP7_75t_L g7104 ( 
.A(n_6637),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6780),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_SL g7106 ( 
.A(n_6895),
.B(n_3765),
.Y(n_7106)
);

NOR2xp33_ASAP7_75t_L g7107 ( 
.A(n_6614),
.B(n_3767),
.Y(n_7107)
);

AOI22xp5_ASAP7_75t_L g7108 ( 
.A1(n_6793),
.A2(n_6877),
.B1(n_6791),
.B2(n_6502),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6783),
.Y(n_7109)
);

NAND2x1p5_ASAP7_75t_L g7110 ( 
.A(n_6621),
.B(n_3832),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6792),
.Y(n_7111)
);

NAND2xp33_ASAP7_75t_L g7112 ( 
.A(n_6804),
.B(n_3769),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6403),
.Y(n_7113)
);

NOR2xp33_ASAP7_75t_L g7114 ( 
.A(n_6808),
.B(n_3771),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_SL g7115 ( 
.A(n_6905),
.B(n_3772),
.Y(n_7115)
);

INVx2_ASAP7_75t_SL g7116 ( 
.A(n_6633),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6755),
.B(n_3773),
.Y(n_7117)
);

INVxp67_ASAP7_75t_L g7118 ( 
.A(n_6885),
.Y(n_7118)
);

NOR2xp33_ASAP7_75t_L g7119 ( 
.A(n_6620),
.B(n_3774),
.Y(n_7119)
);

NAND3xp33_ASAP7_75t_L g7120 ( 
.A(n_6634),
.B(n_3779),
.C(n_3775),
.Y(n_7120)
);

NAND2xp5_ASAP7_75t_L g7121 ( 
.A(n_6756),
.B(n_3780),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6413),
.Y(n_7122)
);

NAND2xp5_ASAP7_75t_SL g7123 ( 
.A(n_6908),
.B(n_3784),
.Y(n_7123)
);

NAND2xp5_ASAP7_75t_L g7124 ( 
.A(n_6768),
.B(n_3787),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_6826),
.B(n_3788),
.Y(n_7125)
);

A2O1A1Ixp33_ASAP7_75t_L g7126 ( 
.A1(n_6482),
.A2(n_6419),
.B(n_6564),
.C(n_6561),
.Y(n_7126)
);

INVxp33_ASAP7_75t_L g7127 ( 
.A(n_6691),
.Y(n_7127)
);

NAND2xp5_ASAP7_75t_L g7128 ( 
.A(n_6425),
.B(n_3789),
.Y(n_7128)
);

AND2x4_ASAP7_75t_L g7129 ( 
.A(n_6598),
.B(n_3834),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_SL g7130 ( 
.A(n_6915),
.B(n_6916),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6429),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6441),
.B(n_3796),
.Y(n_7132)
);

OAI22xp5_ASAP7_75t_L g7133 ( 
.A1(n_6649),
.A2(n_3803),
.B1(n_3804),
.B2(n_3799),
.Y(n_7133)
);

OAI22xp33_ASAP7_75t_L g7134 ( 
.A1(n_6771),
.A2(n_3806),
.B1(n_3808),
.B2(n_3805),
.Y(n_7134)
);

INVxp67_ASAP7_75t_L g7135 ( 
.A(n_6749),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_L g7136 ( 
.A(n_6447),
.B(n_3810),
.Y(n_7136)
);

NAND2xp5_ASAP7_75t_L g7137 ( 
.A(n_6467),
.B(n_3811),
.Y(n_7137)
);

NAND2xp5_ASAP7_75t_L g7138 ( 
.A(n_6471),
.B(n_3815),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_6519),
.B(n_3816),
.Y(n_7139)
);

INVx3_ASAP7_75t_L g7140 ( 
.A(n_6391),
.Y(n_7140)
);

INVx2_ASAP7_75t_L g7141 ( 
.A(n_6800),
.Y(n_7141)
);

NOR2xp33_ASAP7_75t_L g7142 ( 
.A(n_6654),
.B(n_3819),
.Y(n_7142)
);

NOR2xp33_ASAP7_75t_L g7143 ( 
.A(n_6432),
.B(n_3820),
.Y(n_7143)
);

BUFx6f_ASAP7_75t_L g7144 ( 
.A(n_6389),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6805),
.Y(n_7145)
);

INVxp67_ASAP7_75t_L g7146 ( 
.A(n_6766),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6737),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_6527),
.B(n_3823),
.Y(n_7148)
);

NOR2xp33_ASAP7_75t_L g7149 ( 
.A(n_6504),
.B(n_3824),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_SL g7150 ( 
.A(n_6745),
.B(n_3826),
.Y(n_7150)
);

NAND2xp5_ASAP7_75t_L g7151 ( 
.A(n_6555),
.B(n_6558),
.Y(n_7151)
);

INVxp67_ASAP7_75t_L g7152 ( 
.A(n_6574),
.Y(n_7152)
);

AND2x2_ASAP7_75t_L g7153 ( 
.A(n_6648),
.B(n_3828),
.Y(n_7153)
);

INVx8_ASAP7_75t_L g7154 ( 
.A(n_6559),
.Y(n_7154)
);

INVx4_ASAP7_75t_L g7155 ( 
.A(n_6395),
.Y(n_7155)
);

INVxp67_ASAP7_75t_SL g7156 ( 
.A(n_6633),
.Y(n_7156)
);

AND2x4_ASAP7_75t_L g7157 ( 
.A(n_6605),
.B(n_3837),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_6698),
.B(n_3833),
.Y(n_7158)
);

NOR3xp33_ASAP7_75t_L g7159 ( 
.A(n_6902),
.B(n_3836),
.C(n_3835),
.Y(n_7159)
);

AND2x4_ASAP7_75t_L g7160 ( 
.A(n_6445),
.B(n_3846),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6802),
.Y(n_7161)
);

CKINVDCx20_ASAP7_75t_R g7162 ( 
.A(n_6535),
.Y(n_7162)
);

O2A1O1Ixp33_ASAP7_75t_L g7163 ( 
.A1(n_6811),
.A2(n_3864),
.B(n_3878),
.C(n_3847),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_6612),
.B(n_6433),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_SL g7165 ( 
.A(n_6862),
.B(n_3838),
.Y(n_7165)
);

AOI22xp33_ASAP7_75t_L g7166 ( 
.A1(n_6729),
.A2(n_3884),
.B1(n_3886),
.B2(n_3881),
.Y(n_7166)
);

INVx2_ASAP7_75t_L g7167 ( 
.A(n_6815),
.Y(n_7167)
);

NOR2xp33_ASAP7_75t_L g7168 ( 
.A(n_6470),
.B(n_3839),
.Y(n_7168)
);

NAND2xp5_ASAP7_75t_SL g7169 ( 
.A(n_6557),
.B(n_3842),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_SL g7170 ( 
.A(n_6690),
.B(n_6753),
.Y(n_7170)
);

INVx2_ASAP7_75t_L g7171 ( 
.A(n_6810),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_L g7172 ( 
.A(n_6450),
.B(n_3843),
.Y(n_7172)
);

INVx2_ASAP7_75t_L g7173 ( 
.A(n_6814),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_L g7174 ( 
.A(n_6474),
.B(n_6458),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6824),
.Y(n_7175)
);

NOR2x1p5_ASAP7_75t_L g7176 ( 
.A(n_6462),
.B(n_3844),
.Y(n_7176)
);

NAND2xp5_ASAP7_75t_L g7177 ( 
.A(n_6852),
.B(n_6853),
.Y(n_7177)
);

OAI22xp5_ASAP7_75t_L g7178 ( 
.A1(n_6417),
.A2(n_3849),
.B1(n_3850),
.B2(n_3848),
.Y(n_7178)
);

NAND2xp5_ASAP7_75t_L g7179 ( 
.A(n_6900),
.B(n_6911),
.Y(n_7179)
);

AND2x2_ASAP7_75t_SL g7180 ( 
.A(n_6774),
.B(n_3889),
.Y(n_7180)
);

NAND2xp5_ASAP7_75t_L g7181 ( 
.A(n_6829),
.B(n_3851),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_L g7182 ( 
.A(n_6837),
.B(n_3852),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_SL g7183 ( 
.A(n_6919),
.B(n_3853),
.Y(n_7183)
);

A2O1A1Ixp33_ASAP7_75t_L g7184 ( 
.A1(n_6404),
.A2(n_3893),
.B(n_3897),
.C(n_3892),
.Y(n_7184)
);

BUFx3_ASAP7_75t_L g7185 ( 
.A(n_6578),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6839),
.Y(n_7186)
);

NAND2xp5_ASAP7_75t_SL g7187 ( 
.A(n_6536),
.B(n_3854),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_SL g7188 ( 
.A(n_6539),
.B(n_3859),
.Y(n_7188)
);

NOR2xp33_ASAP7_75t_L g7189 ( 
.A(n_6887),
.B(n_3863),
.Y(n_7189)
);

NAND2xp5_ASAP7_75t_L g7190 ( 
.A(n_6842),
.B(n_3866),
.Y(n_7190)
);

AND2x2_ASAP7_75t_SL g7191 ( 
.A(n_6588),
.B(n_3898),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6840),
.Y(n_7192)
);

AND2x2_ASAP7_75t_L g7193 ( 
.A(n_6713),
.B(n_3867),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_6846),
.B(n_3868),
.Y(n_7194)
);

NOR2xp33_ASAP7_75t_L g7195 ( 
.A(n_6705),
.B(n_3869),
.Y(n_7195)
);

NOR2xp33_ASAP7_75t_L g7196 ( 
.A(n_6741),
.B(n_3870),
.Y(n_7196)
);

NAND2xp5_ASAP7_75t_L g7197 ( 
.A(n_6495),
.B(n_3871),
.Y(n_7197)
);

INVx3_ASAP7_75t_L g7198 ( 
.A(n_6473),
.Y(n_7198)
);

NAND2x1p5_ASAP7_75t_L g7199 ( 
.A(n_6408),
.B(n_3900),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_SL g7200 ( 
.A(n_6804),
.B(n_3875),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_SL g7201 ( 
.A(n_6691),
.B(n_6772),
.Y(n_7201)
);

NOR2xp33_ASAP7_75t_L g7202 ( 
.A(n_6920),
.B(n_3876),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_6851),
.Y(n_7203)
);

NAND2xp5_ASAP7_75t_SL g7204 ( 
.A(n_6825),
.B(n_3879),
.Y(n_7204)
);

INVxp67_ASAP7_75t_L g7205 ( 
.A(n_6660),
.Y(n_7205)
);

NOR2xp67_ASAP7_75t_L g7206 ( 
.A(n_6706),
.B(n_3883),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_SL g7207 ( 
.A(n_6679),
.B(n_3887),
.Y(n_7207)
);

INVx2_ASAP7_75t_L g7208 ( 
.A(n_6856),
.Y(n_7208)
);

NAND2xp5_ASAP7_75t_SL g7209 ( 
.A(n_6686),
.B(n_3888),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6511),
.B(n_3890),
.Y(n_7210)
);

INVxp67_ASAP7_75t_L g7211 ( 
.A(n_6823),
.Y(n_7211)
);

BUFx8_ASAP7_75t_L g7212 ( 
.A(n_6410),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6813),
.Y(n_7213)
);

INVx2_ASAP7_75t_SL g7214 ( 
.A(n_6646),
.Y(n_7214)
);

INVx8_ASAP7_75t_L g7215 ( 
.A(n_6559),
.Y(n_7215)
);

NOR2xp33_ASAP7_75t_L g7216 ( 
.A(n_6922),
.B(n_3891),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6841),
.Y(n_7217)
);

NAND2xp33_ASAP7_75t_L g7218 ( 
.A(n_6728),
.B(n_3895),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_6514),
.B(n_3896),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6857),
.Y(n_7220)
);

INVx2_ASAP7_75t_L g7221 ( 
.A(n_6854),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_6849),
.Y(n_7222)
);

INVx2_ASAP7_75t_L g7223 ( 
.A(n_6855),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_6692),
.Y(n_7224)
);

INVx2_ASAP7_75t_L g7225 ( 
.A(n_6377),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_6739),
.Y(n_7226)
);

NAND2xp5_ASAP7_75t_L g7227 ( 
.A(n_6521),
.B(n_3904),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_SL g7228 ( 
.A(n_6868),
.B(n_3905),
.Y(n_7228)
);

BUFx8_ASAP7_75t_L g7229 ( 
.A(n_6524),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_6525),
.B(n_3908),
.Y(n_7230)
);

NOR2xp33_ASAP7_75t_L g7231 ( 
.A(n_6873),
.B(n_3911),
.Y(n_7231)
);

INVx2_ASAP7_75t_L g7232 ( 
.A(n_6761),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_6763),
.Y(n_7233)
);

NAND2xp5_ASAP7_75t_L g7234 ( 
.A(n_6533),
.B(n_6537),
.Y(n_7234)
);

OR2x2_ASAP7_75t_L g7235 ( 
.A(n_6457),
.B(n_3915),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_6573),
.B(n_3916),
.Y(n_7236)
);

OAI22xp5_ASAP7_75t_L g7237 ( 
.A1(n_6827),
.A2(n_3925),
.B1(n_3929),
.B2(n_3924),
.Y(n_7237)
);

OAI221xp5_ASAP7_75t_L g7238 ( 
.A1(n_6913),
.A2(n_3937),
.B1(n_3938),
.B2(n_3936),
.C(n_3930),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_6775),
.Y(n_7239)
);

NOR2xp33_ASAP7_75t_SL g7240 ( 
.A(n_6715),
.B(n_3942),
.Y(n_7240)
);

INVx2_ASAP7_75t_L g7241 ( 
.A(n_6786),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_6628),
.B(n_3945),
.Y(n_7242)
);

NOR2xp33_ASAP7_75t_L g7243 ( 
.A(n_6894),
.B(n_3949),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_6641),
.B(n_3950),
.Y(n_7244)
);

INVx8_ASAP7_75t_L g7245 ( 
.A(n_6880),
.Y(n_7245)
);

NAND2xp5_ASAP7_75t_L g7246 ( 
.A(n_6484),
.B(n_3952),
.Y(n_7246)
);

OR2x6_ASAP7_75t_L g7247 ( 
.A(n_6508),
.B(n_6528),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_6912),
.B(n_3953),
.Y(n_7248)
);

NOR2xp33_ASAP7_75t_L g7249 ( 
.A(n_6898),
.B(n_6434),
.Y(n_7249)
);

NAND2xp5_ASAP7_75t_SL g7250 ( 
.A(n_6879),
.B(n_3954),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_SL g7251 ( 
.A(n_6596),
.B(n_3960),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6817),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6820),
.Y(n_7253)
);

NOR2xp33_ASAP7_75t_L g7254 ( 
.A(n_6436),
.B(n_3962),
.Y(n_7254)
);

BUFx6f_ASAP7_75t_L g7255 ( 
.A(n_6389),
.Y(n_7255)
);

INVx2_ASAP7_75t_L g7256 ( 
.A(n_6629),
.Y(n_7256)
);

AOI22xp33_ASAP7_75t_L g7257 ( 
.A1(n_6784),
.A2(n_3909),
.B1(n_3914),
.B2(n_3903),
.Y(n_7257)
);

INVxp67_ASAP7_75t_L g7258 ( 
.A(n_6863),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_6540),
.B(n_6871),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6719),
.B(n_3963),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_L g7261 ( 
.A(n_6860),
.B(n_3967),
.Y(n_7261)
);

NAND2xp5_ASAP7_75t_SL g7262 ( 
.A(n_6744),
.B(n_3968),
.Y(n_7262)
);

NAND2xp5_ASAP7_75t_L g7263 ( 
.A(n_6663),
.B(n_6832),
.Y(n_7263)
);

NAND2xp5_ASAP7_75t_L g7264 ( 
.A(n_6833),
.B(n_3970),
.Y(n_7264)
);

NAND3xp33_ASAP7_75t_L g7265 ( 
.A(n_6594),
.B(n_3976),
.C(n_3971),
.Y(n_7265)
);

OR2x2_ASAP7_75t_L g7266 ( 
.A(n_6695),
.B(n_3977),
.Y(n_7266)
);

A2O1A1Ixp33_ASAP7_75t_L g7267 ( 
.A1(n_6650),
.A2(n_3923),
.B(n_3928),
.C(n_3917),
.Y(n_7267)
);

NAND2xp5_ASAP7_75t_L g7268 ( 
.A(n_6909),
.B(n_3989),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_6523),
.B(n_3994),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_6861),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_6864),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6656),
.Y(n_7272)
);

NAND2xp33_ASAP7_75t_L g7273 ( 
.A(n_6728),
.B(n_3995),
.Y(n_7273)
);

AND2x2_ASAP7_75t_SL g7274 ( 
.A(n_6865),
.B(n_6639),
.Y(n_7274)
);

INVxp67_ASAP7_75t_L g7275 ( 
.A(n_6897),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_6635),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_L g7277 ( 
.A(n_6500),
.B(n_3998),
.Y(n_7277)
);

NAND2xp5_ASAP7_75t_L g7278 ( 
.A(n_6806),
.B(n_4002),
.Y(n_7278)
);

INVx2_ASAP7_75t_L g7279 ( 
.A(n_6838),
.Y(n_7279)
);

NAND2xp5_ASAP7_75t_L g7280 ( 
.A(n_6513),
.B(n_4003),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_6670),
.Y(n_7281)
);

NAND2xp5_ASAP7_75t_SL g7282 ( 
.A(n_6790),
.B(n_4006),
.Y(n_7282)
);

INVx2_ASAP7_75t_L g7283 ( 
.A(n_6818),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_6452),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_6699),
.B(n_4008),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_SL g7286 ( 
.A(n_6831),
.B(n_4013),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_6676),
.B(n_4016),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_6667),
.B(n_4017),
.Y(n_7288)
);

OR2x2_ASAP7_75t_L g7289 ( 
.A(n_6563),
.B(n_4022),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_L g7290 ( 
.A(n_6689),
.B(n_4023),
.Y(n_7290)
);

NAND2xp5_ASAP7_75t_L g7291 ( 
.A(n_6714),
.B(n_4025),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_6735),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_6456),
.Y(n_7293)
);

NOR2xp33_ASAP7_75t_SL g7294 ( 
.A(n_6718),
.B(n_4028),
.Y(n_7294)
);

NOR3xp33_ASAP7_75t_L g7295 ( 
.A(n_6697),
.B(n_4031),
.C(n_4029),
.Y(n_7295)
);

AO221x1_ASAP7_75t_L g7296 ( 
.A1(n_6796),
.A2(n_6834),
.B1(n_6678),
.B2(n_6414),
.C(n_6587),
.Y(n_7296)
);

NOR2xp67_ASAP7_75t_L g7297 ( 
.A(n_6723),
.B(n_4032),
.Y(n_7297)
);

NAND2xp5_ASAP7_75t_SL g7298 ( 
.A(n_6831),
.B(n_4033),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6816),
.Y(n_7299)
);

NAND2xp5_ASAP7_75t_L g7300 ( 
.A(n_6859),
.B(n_4034),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_SL g7301 ( 
.A(n_6599),
.B(n_4036),
.Y(n_7301)
);

AOI22xp5_ASAP7_75t_L g7302 ( 
.A1(n_6376),
.A2(n_4039),
.B1(n_4041),
.B2(n_4037),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_SL g7303 ( 
.A(n_6646),
.B(n_4045),
.Y(n_7303)
);

INVx2_ASAP7_75t_L g7304 ( 
.A(n_6465),
.Y(n_7304)
);

INVx8_ASAP7_75t_L g7305 ( 
.A(n_6880),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6816),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_6379),
.Y(n_7307)
);

NAND2xp33_ASAP7_75t_SL g7308 ( 
.A(n_6742),
.B(n_4048),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_SL g7309 ( 
.A(n_6659),
.B(n_4050),
.Y(n_7309)
);

INVx2_ASAP7_75t_SL g7310 ( 
.A(n_6659),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_L g7311 ( 
.A(n_6661),
.B(n_4052),
.Y(n_7311)
);

INVx2_ASAP7_75t_SL g7312 ( 
.A(n_6669),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_6468),
.Y(n_7313)
);

NAND2xp5_ASAP7_75t_L g7314 ( 
.A(n_6622),
.B(n_4056),
.Y(n_7314)
);

NOR2xp33_ASAP7_75t_L g7315 ( 
.A(n_6896),
.B(n_4058),
.Y(n_7315)
);

NAND2xp5_ASAP7_75t_SL g7316 ( 
.A(n_6669),
.B(n_4060),
.Y(n_7316)
);

AOI22xp5_ASAP7_75t_L g7317 ( 
.A1(n_6725),
.A2(n_4063),
.B1(n_4078),
.B2(n_4062),
.Y(n_7317)
);

BUFx3_ASAP7_75t_L g7318 ( 
.A(n_6684),
.Y(n_7318)
);

AND2x4_ASAP7_75t_L g7319 ( 
.A(n_6380),
.B(n_3933),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_6622),
.B(n_4080),
.Y(n_7320)
);

NOR2xp67_ASAP7_75t_L g7321 ( 
.A(n_6731),
.B(n_4081),
.Y(n_7321)
);

INVx2_ASAP7_75t_L g7322 ( 
.A(n_6492),
.Y(n_7322)
);

INVx2_ASAP7_75t_L g7323 ( 
.A(n_6498),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_6625),
.B(n_4083),
.Y(n_7324)
);

NOR2xp33_ASAP7_75t_L g7325 ( 
.A(n_6910),
.B(n_4085),
.Y(n_7325)
);

NAND2xp5_ASAP7_75t_SL g7326 ( 
.A(n_6730),
.B(n_4086),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_6503),
.Y(n_7327)
);

NOR2xp33_ASAP7_75t_L g7328 ( 
.A(n_6722),
.B(n_4087),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_6545),
.Y(n_7329)
);

NAND2xp5_ASAP7_75t_L g7330 ( 
.A(n_6625),
.B(n_4093),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_L g7331 ( 
.A(n_6665),
.B(n_4094),
.Y(n_7331)
);

NOR2xp67_ASAP7_75t_L g7332 ( 
.A(n_6733),
.B(n_4100),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_SL g7333 ( 
.A(n_6730),
.B(n_6651),
.Y(n_7333)
);

INVxp33_ASAP7_75t_L g7334 ( 
.A(n_6390),
.Y(n_7334)
);

INVxp67_ASAP7_75t_SL g7335 ( 
.A(n_6439),
.Y(n_7335)
);

AND2x2_ASAP7_75t_L g7336 ( 
.A(n_6876),
.B(n_4101),
.Y(n_7336)
);

INVx2_ASAP7_75t_L g7337 ( 
.A(n_6552),
.Y(n_7337)
);

AND2x2_ASAP7_75t_L g7338 ( 
.A(n_6750),
.B(n_4102),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_6579),
.Y(n_7339)
);

NAND2xp5_ASAP7_75t_SL g7340 ( 
.A(n_6651),
.B(n_6671),
.Y(n_7340)
);

BUFx3_ASAP7_75t_L g7341 ( 
.A(n_6684),
.Y(n_7341)
);

INVx2_ASAP7_75t_L g7342 ( 
.A(n_6590),
.Y(n_7342)
);

BUFx6f_ASAP7_75t_L g7343 ( 
.A(n_6439),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_L g7344 ( 
.A(n_6665),
.B(n_4104),
.Y(n_7344)
);

OR2x2_ASAP7_75t_L g7345 ( 
.A(n_6870),
.B(n_4107),
.Y(n_7345)
);

INVx2_ASAP7_75t_L g7346 ( 
.A(n_6464),
.Y(n_7346)
);

NAND2xp5_ASAP7_75t_L g7347 ( 
.A(n_6685),
.B(n_4110),
.Y(n_7347)
);

AO221x1_ASAP7_75t_L g7348 ( 
.A1(n_6444),
.A2(n_3944),
.B1(n_3947),
.B2(n_3943),
.C(n_3934),
.Y(n_7348)
);

NOR2xp33_ASAP7_75t_L g7349 ( 
.A(n_6740),
.B(n_4114),
.Y(n_7349)
);

NAND2xp5_ASAP7_75t_SL g7350 ( 
.A(n_6671),
.B(n_4118),
.Y(n_7350)
);

AND2x2_ASAP7_75t_L g7351 ( 
.A(n_6553),
.B(n_4121),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6843),
.Y(n_7352)
);

NAND2xp5_ASAP7_75t_L g7353 ( 
.A(n_6685),
.B(n_4122),
.Y(n_7353)
);

INVx2_ASAP7_75t_L g7354 ( 
.A(n_6464),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_6693),
.B(n_4125),
.Y(n_7355)
);

NOR2xp33_ASAP7_75t_L g7356 ( 
.A(n_6743),
.B(n_4126),
.Y(n_7356)
);

BUFx3_ASAP7_75t_L g7357 ( 
.A(n_6694),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_6472),
.Y(n_7358)
);

AND2x4_ASAP7_75t_L g7359 ( 
.A(n_6480),
.B(n_3951),
.Y(n_7359)
);

AOI221xp5_ASAP7_75t_L g7360 ( 
.A1(n_6584),
.A2(n_3961),
.B1(n_3964),
.B2(n_3959),
.C(n_3955),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6843),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6421),
.Y(n_7362)
);

NOR2xp33_ASAP7_75t_L g7363 ( 
.A(n_6757),
.B(n_4127),
.Y(n_7363)
);

NAND2xp5_ASAP7_75t_L g7364 ( 
.A(n_6693),
.B(n_4128),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_SL g7365 ( 
.A(n_6688),
.B(n_4129),
.Y(n_7365)
);

INVx1_ASAP7_75t_SL g7366 ( 
.A(n_6716),
.Y(n_7366)
);

INVx8_ASAP7_75t_L g7367 ( 
.A(n_6688),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_SL g7368 ( 
.A(n_6408),
.B(n_4135),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_6472),
.Y(n_7369)
);

INVx2_ASAP7_75t_L g7370 ( 
.A(n_6520),
.Y(n_7370)
);

NAND2xp5_ASAP7_75t_L g7371 ( 
.A(n_6847),
.B(n_4137),
.Y(n_7371)
);

INVx2_ASAP7_75t_L g7372 ( 
.A(n_6520),
.Y(n_7372)
);

NOR2xp33_ASAP7_75t_L g7373 ( 
.A(n_6778),
.B(n_4140),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_SL g7374 ( 
.A(n_6409),
.B(n_4142),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_6819),
.B(n_6453),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6531),
.Y(n_7376)
);

AND2x2_ASAP7_75t_L g7377 ( 
.A(n_6460),
.B(n_6549),
.Y(n_7377)
);

NAND2xp5_ASAP7_75t_L g7378 ( 
.A(n_6453),
.B(n_4143),
.Y(n_7378)
);

NAND2xp33_ASAP7_75t_SL g7379 ( 
.A(n_6531),
.B(n_4146),
.Y(n_7379)
);

NAND2xp5_ASAP7_75t_SL g7380 ( 
.A(n_6409),
.B(n_4147),
.Y(n_7380)
);

NAND2xp5_ASAP7_75t_L g7381 ( 
.A(n_6565),
.B(n_4148),
.Y(n_7381)
);

NAND2xp5_ASAP7_75t_L g7382 ( 
.A(n_6565),
.B(n_4149),
.Y(n_7382)
);

NAND2xp5_ASAP7_75t_SL g7383 ( 
.A(n_6383),
.B(n_4150),
.Y(n_7383)
);

AND2x2_ASAP7_75t_L g7384 ( 
.A(n_6874),
.B(n_4153),
.Y(n_7384)
);

INVx2_ASAP7_75t_L g7385 ( 
.A(n_6532),
.Y(n_7385)
);

NOR3xp33_ASAP7_75t_L g7386 ( 
.A(n_6700),
.B(n_4157),
.C(n_4155),
.Y(n_7386)
);

BUFx6f_ASAP7_75t_L g7387 ( 
.A(n_6532),
.Y(n_7387)
);

NAND2xp5_ASAP7_75t_L g7388 ( 
.A(n_6782),
.B(n_4158),
.Y(n_7388)
);

NOR2xp33_ASAP7_75t_L g7389 ( 
.A(n_6801),
.B(n_4160),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_L g7390 ( 
.A(n_6830),
.B(n_4161),
.Y(n_7390)
);

NAND2xp5_ASAP7_75t_L g7391 ( 
.A(n_6858),
.B(n_4162),
.Y(n_7391)
);

NAND2xp5_ASAP7_75t_L g7392 ( 
.A(n_6858),
.B(n_4163),
.Y(n_7392)
);

INVx2_ASAP7_75t_SL g7393 ( 
.A(n_6607),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_6607),
.Y(n_7394)
);

OR2x6_ASAP7_75t_L g7395 ( 
.A(n_6422),
.B(n_6449),
.Y(n_7395)
);

NAND2xp33_ASAP7_75t_L g7396 ( 
.A(n_6694),
.B(n_4168),
.Y(n_7396)
);

INVx1_ASAP7_75t_L g7397 ( 
.A(n_6570),
.Y(n_7397)
);

INVx8_ASAP7_75t_L g7398 ( 
.A(n_6402),
.Y(n_7398)
);

INVxp67_ASAP7_75t_SL g7399 ( 
.A(n_6726),
.Y(n_7399)
);

NAND2xp5_ASAP7_75t_SL g7400 ( 
.A(n_6562),
.B(n_4171),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_L g7401 ( 
.A(n_6493),
.B(n_4172),
.Y(n_7401)
);

NOR2xp33_ASAP7_75t_L g7402 ( 
.A(n_6627),
.B(n_6662),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_SL g7403 ( 
.A(n_6572),
.B(n_6589),
.Y(n_7403)
);

NAND2xp5_ASAP7_75t_SL g7404 ( 
.A(n_6600),
.B(n_4173),
.Y(n_7404)
);

NOR2xp33_ASAP7_75t_L g7405 ( 
.A(n_6727),
.B(n_4176),
.Y(n_7405)
);

BUFx6f_ASAP7_75t_L g7406 ( 
.A(n_6759),
.Y(n_7406)
);

AOI22xp33_ASAP7_75t_L g7407 ( 
.A1(n_6446),
.A2(n_3982),
.B1(n_3984),
.B2(n_3978),
.Y(n_7407)
);

NAND2xp33_ASAP7_75t_L g7408 ( 
.A(n_6759),
.B(n_4177),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_6632),
.Y(n_7409)
);

AND2x2_ASAP7_75t_L g7410 ( 
.A(n_6710),
.B(n_4178),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6509),
.Y(n_7411)
);

OAI221xp5_ASAP7_75t_L g7412 ( 
.A1(n_6630),
.A2(n_4184),
.B1(n_4188),
.B2(n_4181),
.C(n_4179),
.Y(n_7412)
);

NOR2xp67_ASAP7_75t_L g7413 ( 
.A(n_6466),
.B(n_4192),
.Y(n_7413)
);

NOR2xp33_ASAP7_75t_L g7414 ( 
.A(n_6534),
.B(n_4194),
.Y(n_7414)
);

NOR3xp33_ASAP7_75t_L g7415 ( 
.A(n_6907),
.B(n_4196),
.C(n_4195),
.Y(n_7415)
);

NAND2xp33_ASAP7_75t_L g7416 ( 
.A(n_6747),
.B(n_4197),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_6568),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6435),
.Y(n_7418)
);

OR2x6_ASAP7_75t_L g7419 ( 
.A(n_6512),
.B(n_3987),
.Y(n_7419)
);

CKINVDCx20_ASAP7_75t_R g7420 ( 
.A(n_6752),
.Y(n_7420)
);

INVxp67_ASAP7_75t_L g7421 ( 
.A(n_6904),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_6666),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6867),
.Y(n_7423)
);

INVxp67_ASAP7_75t_L g7424 ( 
.A(n_6567),
.Y(n_7424)
);

NAND2xp5_ASAP7_75t_SL g7425 ( 
.A(n_6640),
.B(n_4199),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_6717),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6932),
.Y(n_7427)
);

INVx2_ASAP7_75t_L g7428 ( 
.A(n_6935),
.Y(n_7428)
);

NAND2xp5_ASAP7_75t_SL g7429 ( 
.A(n_7179),
.B(n_6518),
.Y(n_7429)
);

INVxp67_ASAP7_75t_L g7430 ( 
.A(n_7092),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_6938),
.Y(n_7431)
);

NAND2x1_ASAP7_75t_L g7432 ( 
.A(n_7208),
.B(n_7220),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_6953),
.Y(n_7433)
);

CKINVDCx20_ASAP7_75t_R g7434 ( 
.A(n_7162),
.Y(n_7434)
);

OAI221xp5_ASAP7_75t_L g7435 ( 
.A1(n_7017),
.A2(n_6893),
.B1(n_6914),
.B2(n_6917),
.C(n_6881),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_6961),
.Y(n_7436)
);

AOI22xp5_ASAP7_75t_L g7437 ( 
.A1(n_6960),
.A2(n_6807),
.B1(n_6624),
.B2(n_6657),
.Y(n_7437)
);

AO22x2_ASAP7_75t_L g7438 ( 
.A1(n_6930),
.A2(n_6677),
.B1(n_6675),
.B2(n_6875),
.Y(n_7438)
);

AOI22xp5_ASAP7_75t_L g7439 ( 
.A1(n_6970),
.A2(n_6560),
.B1(n_6586),
.B2(n_6580),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6966),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_6991),
.Y(n_7441)
);

BUFx8_ASAP7_75t_L g7442 ( 
.A(n_6924),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_6992),
.Y(n_7443)
);

AO22x2_ASAP7_75t_L g7444 ( 
.A1(n_6934),
.A2(n_6626),
.B1(n_6610),
.B2(n_6821),
.Y(n_7444)
);

AND2x4_ASAP7_75t_L g7445 ( 
.A(n_7185),
.B(n_6609),
.Y(n_7445)
);

AO22x1_ASAP7_75t_L g7446 ( 
.A1(n_6997),
.A2(n_6455),
.B1(n_6903),
.B2(n_6899),
.Y(n_7446)
);

INVx4_ASAP7_75t_L g7447 ( 
.A(n_7406),
.Y(n_7447)
);

AO22x2_ASAP7_75t_L g7448 ( 
.A1(n_6926),
.A2(n_4014),
.B1(n_4015),
.B2(n_3992),
.Y(n_7448)
);

BUFx8_ASAP7_75t_L g7449 ( 
.A(n_6951),
.Y(n_7449)
);

BUFx3_ASAP7_75t_L g7450 ( 
.A(n_7104),
.Y(n_7450)
);

AO22x2_ASAP7_75t_L g7451 ( 
.A1(n_7005),
.A2(n_6981),
.B1(n_7362),
.B2(n_7426),
.Y(n_7451)
);

INVx2_ASAP7_75t_L g7452 ( 
.A(n_6993),
.Y(n_7452)
);

AOI22xp5_ASAP7_75t_L g7453 ( 
.A1(n_6943),
.A2(n_6787),
.B1(n_6581),
.B2(n_6658),
.Y(n_7453)
);

INVx2_ASAP7_75t_SL g7454 ( 
.A(n_7406),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_7010),
.Y(n_7455)
);

AO22x2_ASAP7_75t_L g7456 ( 
.A1(n_7174),
.A2(n_4035),
.B1(n_4040),
.B2(n_4021),
.Y(n_7456)
);

AND2x2_ASAP7_75t_L g7457 ( 
.A(n_7043),
.B(n_6407),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7025),
.Y(n_7458)
);

AO22x2_ASAP7_75t_L g7459 ( 
.A1(n_6928),
.A2(n_4047),
.B1(n_4059),
.B2(n_4044),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7041),
.Y(n_7460)
);

NAND2xp33_ASAP7_75t_L g7461 ( 
.A(n_7126),
.B(n_7164),
.Y(n_7461)
);

NAND2x1p5_ASAP7_75t_L g7462 ( 
.A(n_7155),
.B(n_6400),
.Y(n_7462)
);

BUFx2_ASAP7_75t_L g7463 ( 
.A(n_6972),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_6977),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_6986),
.Y(n_7465)
);

INVx2_ASAP7_75t_L g7466 ( 
.A(n_7049),
.Y(n_7466)
);

AO22x2_ASAP7_75t_L g7467 ( 
.A1(n_6923),
.A2(n_4069),
.B1(n_4072),
.B2(n_4061),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6999),
.Y(n_7468)
);

OAI221xp5_ASAP7_75t_L g7469 ( 
.A1(n_7189),
.A2(n_6487),
.B1(n_6386),
.B2(n_6822),
.C(n_6795),
.Y(n_7469)
);

AOI22xp33_ASAP7_75t_L g7470 ( 
.A1(n_7296),
.A2(n_6674),
.B1(n_6515),
.B2(n_6769),
.Y(n_7470)
);

CKINVDCx5p33_ASAP7_75t_R g7471 ( 
.A(n_6954),
.Y(n_7471)
);

BUFx3_ASAP7_75t_L g7472 ( 
.A(n_7245),
.Y(n_7472)
);

NAND2xp5_ASAP7_75t_L g7473 ( 
.A(n_7147),
.B(n_6631),
.Y(n_7473)
);

AO22x2_ASAP7_75t_L g7474 ( 
.A1(n_6925),
.A2(n_4077),
.B1(n_4090),
.B2(n_4076),
.Y(n_7474)
);

INVx2_ASAP7_75t_L g7475 ( 
.A(n_7223),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_7061),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7074),
.Y(n_7477)
);

AO22x2_ASAP7_75t_L g7478 ( 
.A1(n_7006),
.A2(n_4096),
.B1(n_4099),
.B2(n_4091),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_7078),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7085),
.Y(n_7480)
);

AO22x2_ASAP7_75t_L g7481 ( 
.A1(n_7252),
.A2(n_4106),
.B1(n_4112),
.B2(n_4105),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7087),
.Y(n_7482)
);

INVx1_ASAP7_75t_L g7483 ( 
.A(n_7093),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_7099),
.Y(n_7484)
);

NAND2x1p5_ASAP7_75t_L g7485 ( 
.A(n_6982),
.B(n_6886),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7105),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_7109),
.Y(n_7487)
);

AO22x2_ASAP7_75t_L g7488 ( 
.A1(n_7253),
.A2(n_4132),
.B1(n_4133),
.B2(n_4117),
.Y(n_7488)
);

NOR2xp67_ASAP7_75t_L g7489 ( 
.A(n_7140),
.B(n_6799),
.Y(n_7489)
);

INVx3_ASAP7_75t_L g7490 ( 
.A(n_6978),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_7111),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_7177),
.B(n_6844),
.Y(n_7492)
);

INVx1_ASAP7_75t_L g7493 ( 
.A(n_7161),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6931),
.Y(n_7494)
);

BUFx10_ASAP7_75t_L g7495 ( 
.A(n_7076),
.Y(n_7495)
);

INVx1_ASAP7_75t_L g7496 ( 
.A(n_6937),
.Y(n_7496)
);

INVx2_ASAP7_75t_L g7497 ( 
.A(n_6942),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_6956),
.Y(n_7498)
);

BUFx6f_ASAP7_75t_L g7499 ( 
.A(n_7144),
.Y(n_7499)
);

CKINVDCx5p33_ASAP7_75t_R g7500 ( 
.A(n_7420),
.Y(n_7500)
);

OAI221xp5_ASAP7_75t_L g7501 ( 
.A1(n_7119),
.A2(n_6899),
.B1(n_6835),
.B2(n_6734),
.C(n_6418),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_6959),
.Y(n_7502)
);

NAND2x1p5_ASAP7_75t_L g7503 ( 
.A(n_7198),
.B(n_6770),
.Y(n_7503)
);

NAND2xp5_ASAP7_75t_L g7504 ( 
.A(n_7234),
.B(n_6850),
.Y(n_7504)
);

BUFx8_ASAP7_75t_L g7505 ( 
.A(n_6974),
.Y(n_7505)
);

INVx1_ASAP7_75t_L g7506 ( 
.A(n_6962),
.Y(n_7506)
);

AOI22xp5_ASAP7_75t_L g7507 ( 
.A1(n_7033),
.A2(n_7039),
.B1(n_7114),
.B2(n_7107),
.Y(n_7507)
);

AO22x2_ASAP7_75t_L g7508 ( 
.A1(n_7011),
.A2(n_7265),
.B1(n_7418),
.B2(n_6933),
.Y(n_7508)
);

AND2x2_ASAP7_75t_L g7509 ( 
.A(n_6955),
.B(n_6866),
.Y(n_7509)
);

INVx1_ASAP7_75t_L g7510 ( 
.A(n_6969),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_6971),
.Y(n_7511)
);

OAI221xp5_ASAP7_75t_L g7512 ( 
.A1(n_7142),
.A2(n_4152),
.B1(n_4169),
.B2(n_4151),
.C(n_4141),
.Y(n_7512)
);

OAI221xp5_ASAP7_75t_L g7513 ( 
.A1(n_7405),
.A2(n_7325),
.B1(n_7108),
.B2(n_7328),
.C(n_7254),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_6983),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7004),
.Y(n_7515)
);

NOR2xp33_ASAP7_75t_L g7516 ( 
.A(n_6936),
.B(n_6828),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7008),
.Y(n_7517)
);

AND2x6_ASAP7_75t_L g7518 ( 
.A(n_7272),
.B(n_4170),
.Y(n_7518)
);

NAND2x1p5_ASAP7_75t_L g7519 ( 
.A(n_6980),
.B(n_7318),
.Y(n_7519)
);

INVx2_ASAP7_75t_L g7520 ( 
.A(n_7031),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7034),
.Y(n_7521)
);

NOR2xp33_ASAP7_75t_L g7522 ( 
.A(n_7071),
.B(n_6878),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7035),
.Y(n_7523)
);

INVx2_ASAP7_75t_L g7524 ( 
.A(n_7171),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7173),
.Y(n_7525)
);

NAND2x1p5_ASAP7_75t_L g7526 ( 
.A(n_7341),
.B(n_4174),
.Y(n_7526)
);

NOR2xp33_ASAP7_75t_L g7527 ( 
.A(n_6940),
.B(n_4202),
.Y(n_7527)
);

INVx2_ASAP7_75t_L g7528 ( 
.A(n_7037),
.Y(n_7528)
);

INVx2_ASAP7_75t_L g7529 ( 
.A(n_7057),
.Y(n_7529)
);

OAI22xp5_ASAP7_75t_L g7530 ( 
.A1(n_7151),
.A2(n_4207),
.B1(n_4208),
.B2(n_4203),
.Y(n_7530)
);

NOR2xp33_ASAP7_75t_L g7531 ( 
.A(n_6941),
.B(n_4209),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_7113),
.Y(n_7532)
);

INVxp67_ASAP7_75t_L g7533 ( 
.A(n_6964),
.Y(n_7533)
);

AND2x6_ASAP7_75t_L g7534 ( 
.A(n_7281),
.B(n_4182),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_7131),
.Y(n_7535)
);

NAND2xp5_ASAP7_75t_L g7536 ( 
.A(n_7068),
.B(n_4191),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7059),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_7122),
.Y(n_7538)
);

INVx3_ASAP7_75t_L g7539 ( 
.A(n_7357),
.Y(n_7539)
);

AO22x2_ASAP7_75t_L g7540 ( 
.A1(n_7292),
.A2(n_4198),
.B1(n_4205),
.B2(n_4193),
.Y(n_7540)
);

AOI22xp5_ASAP7_75t_L g7541 ( 
.A1(n_6950),
.A2(n_6998),
.B1(n_6958),
.B2(n_6967),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7175),
.Y(n_7542)
);

NOR2xp67_ASAP7_75t_L g7543 ( 
.A(n_7118),
.B(n_1),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7192),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7073),
.Y(n_7545)
);

CKINVDCx5p33_ASAP7_75t_R g7546 ( 
.A(n_6976),
.Y(n_7546)
);

AO22x2_ASAP7_75t_L g7547 ( 
.A1(n_7299),
.A2(n_4217),
.B1(n_4219),
.B2(n_4212),
.Y(n_7547)
);

AO22x2_ASAP7_75t_L g7548 ( 
.A1(n_7306),
.A2(n_4237),
.B1(n_4241),
.B2(n_4227),
.Y(n_7548)
);

CKINVDCx5p33_ASAP7_75t_R g7549 ( 
.A(n_7212),
.Y(n_7549)
);

AND2x6_ASAP7_75t_L g7550 ( 
.A(n_7226),
.B(n_4242),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7270),
.Y(n_7551)
);

AO22x2_ASAP7_75t_L g7552 ( 
.A1(n_6927),
.A2(n_4260),
.B1(n_4262),
.B2(n_4243),
.Y(n_7552)
);

AO22x2_ASAP7_75t_L g7553 ( 
.A1(n_7259),
.A2(n_4265),
.B1(n_4278),
.B2(n_4263),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_6963),
.B(n_4280),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_7271),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7186),
.Y(n_7556)
);

OAI221xp5_ASAP7_75t_L g7557 ( 
.A1(n_7349),
.A2(n_7356),
.B1(n_7389),
.B2(n_7373),
.C(n_7363),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7203),
.Y(n_7558)
);

AO22x2_ASAP7_75t_L g7559 ( 
.A1(n_7352),
.A2(n_4285),
.B1(n_4282),
.B2(n_4),
.Y(n_7559)
);

AND2x4_ASAP7_75t_L g7560 ( 
.A(n_7283),
.B(n_4210),
.Y(n_7560)
);

NAND2xp5_ASAP7_75t_L g7561 ( 
.A(n_6947),
.B(n_4211),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_7141),
.Y(n_7562)
);

AO22x2_ASAP7_75t_L g7563 ( 
.A1(n_7361),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_7563)
);

AOI22xp33_ASAP7_75t_L g7564 ( 
.A1(n_7412),
.A2(n_4214),
.B1(n_4215),
.B2(n_4213),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_7145),
.Y(n_7565)
);

AND2x4_ASAP7_75t_L g7566 ( 
.A(n_7409),
.B(n_4216),
.Y(n_7566)
);

BUFx8_ASAP7_75t_L g7567 ( 
.A(n_7377),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7167),
.Y(n_7568)
);

NAND2xp5_ASAP7_75t_L g7569 ( 
.A(n_7232),
.B(n_4218),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_7213),
.Y(n_7570)
);

AO22x2_ASAP7_75t_L g7571 ( 
.A1(n_7351),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7217),
.Y(n_7572)
);

INVx2_ASAP7_75t_SL g7573 ( 
.A(n_7367),
.Y(n_7573)
);

AND2x4_ASAP7_75t_L g7574 ( 
.A(n_7395),
.B(n_4220),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_L g7575 ( 
.A(n_7233),
.B(n_4221),
.Y(n_7575)
);

OAI221xp5_ASAP7_75t_L g7576 ( 
.A1(n_7243),
.A2(n_4234),
.B1(n_4235),
.B2(n_4226),
.C(n_4222),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7222),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_7224),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7221),
.Y(n_7579)
);

OAI22xp5_ASAP7_75t_SL g7580 ( 
.A1(n_7191),
.A2(n_4240),
.B1(n_4245),
.B2(n_4239),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7423),
.Y(n_7581)
);

AOI22xp5_ASAP7_75t_L g7582 ( 
.A1(n_7249),
.A2(n_4248),
.B1(n_4251),
.B2(n_4246),
.Y(n_7582)
);

INVx2_ASAP7_75t_L g7583 ( 
.A(n_7256),
.Y(n_7583)
);

AOI22xp5_ASAP7_75t_SL g7584 ( 
.A1(n_7045),
.A2(n_4254),
.B1(n_4256),
.B2(n_4253),
.Y(n_7584)
);

INVx2_ASAP7_75t_L g7585 ( 
.A(n_7276),
.Y(n_7585)
);

INVx1_ASAP7_75t_L g7586 ( 
.A(n_7284),
.Y(n_7586)
);

BUFx8_ASAP7_75t_L g7587 ( 
.A(n_7144),
.Y(n_7587)
);

NAND2x1p5_ASAP7_75t_L g7588 ( 
.A(n_7255),
.B(n_413),
.Y(n_7588)
);

NAND2xp5_ASAP7_75t_L g7589 ( 
.A(n_7239),
.B(n_4257),
.Y(n_7589)
);

NAND2x1p5_ASAP7_75t_L g7590 ( 
.A(n_7255),
.B(n_414),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7293),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_7304),
.Y(n_7592)
);

OAI221xp5_ASAP7_75t_L g7593 ( 
.A1(n_7414),
.A2(n_4264),
.B1(n_4266),
.B2(n_4259),
.C(n_4258),
.Y(n_7593)
);

NAND2xp5_ASAP7_75t_L g7594 ( 
.A(n_7241),
.B(n_4267),
.Y(n_7594)
);

OAI221xp5_ASAP7_75t_L g7595 ( 
.A1(n_7077),
.A2(n_4270),
.B1(n_4271),
.B2(n_4269),
.C(n_4268),
.Y(n_7595)
);

NOR3xp33_ASAP7_75t_L g7596 ( 
.A(n_6957),
.B(n_4274),
.C(n_4272),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_7313),
.Y(n_7597)
);

AOI22xp5_ASAP7_75t_L g7598 ( 
.A1(n_7079),
.A2(n_4279),
.B1(n_4281),
.B2(n_4276),
.Y(n_7598)
);

AO22x2_ASAP7_75t_L g7599 ( 
.A1(n_7410),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_7599)
);

AOI22xp5_ASAP7_75t_L g7600 ( 
.A1(n_7086),
.A2(n_7102),
.B1(n_7402),
.B2(n_7196),
.Y(n_7600)
);

AO22x2_ASAP7_75t_L g7601 ( 
.A1(n_7120),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_7601)
);

AND2x4_ASAP7_75t_L g7602 ( 
.A(n_7395),
.B(n_4286),
.Y(n_7602)
);

AND2x6_ASAP7_75t_L g7603 ( 
.A(n_7422),
.B(n_6),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7322),
.Y(n_7604)
);

BUFx8_ASAP7_75t_L g7605 ( 
.A(n_7343),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_7323),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7337),
.Y(n_7607)
);

BUFx2_ASAP7_75t_L g7608 ( 
.A(n_7095),
.Y(n_7608)
);

AO22x2_ASAP7_75t_L g7609 ( 
.A1(n_6949),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_7609)
);

AND2x6_ASAP7_75t_L g7610 ( 
.A(n_7307),
.B(n_7),
.Y(n_7610)
);

AOI22xp33_ASAP7_75t_L g7611 ( 
.A1(n_7135),
.A2(n_4289),
.B1(n_4291),
.B2(n_4288),
.Y(n_7611)
);

INVx2_ASAP7_75t_L g7612 ( 
.A(n_7342),
.Y(n_7612)
);

NAND2xp5_ASAP7_75t_L g7613 ( 
.A(n_7263),
.B(n_7202),
.Y(n_7613)
);

AND2x4_ASAP7_75t_L g7614 ( 
.A(n_7247),
.B(n_4292),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_7315),
.B(n_4297),
.Y(n_7615)
);

AND2x4_ASAP7_75t_L g7616 ( 
.A(n_7247),
.B(n_4298),
.Y(n_7616)
);

NAND2xp5_ASAP7_75t_L g7617 ( 
.A(n_6948),
.B(n_4302),
.Y(n_7617)
);

AOI22xp5_ASAP7_75t_L g7618 ( 
.A1(n_7195),
.A2(n_7069),
.B1(n_7055),
.B2(n_7231),
.Y(n_7618)
);

NAND2xp5_ASAP7_75t_L g7619 ( 
.A(n_7172),
.B(n_4304),
.Y(n_7619)
);

AND2x4_ASAP7_75t_L g7620 ( 
.A(n_7399),
.B(n_4307),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7327),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7329),
.Y(n_7622)
);

AO22x2_ASAP7_75t_L g7623 ( 
.A1(n_7159),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_7623)
);

INVxp67_ASAP7_75t_L g7624 ( 
.A(n_7345),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7339),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_6944),
.Y(n_7626)
);

AO22x2_ASAP7_75t_L g7627 ( 
.A1(n_7130),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7084),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7094),
.Y(n_7629)
);

INVx2_ASAP7_75t_L g7630 ( 
.A(n_7225),
.Y(n_7630)
);

AO22x2_ASAP7_75t_L g7631 ( 
.A1(n_7375),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_7631)
);

AOI22xp5_ASAP7_75t_L g7632 ( 
.A1(n_7146),
.A2(n_416),
.B1(n_417),
.B2(n_415),
.Y(n_7632)
);

OAI221xp5_ASAP7_75t_L g7633 ( 
.A1(n_7311),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.C(n_15),
.Y(n_7633)
);

OR2x6_ASAP7_75t_L g7634 ( 
.A(n_7245),
.B(n_416),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_7096),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7097),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7098),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7117),
.Y(n_7638)
);

INVx2_ASAP7_75t_L g7639 ( 
.A(n_7121),
.Y(n_7639)
);

INVx2_ASAP7_75t_L g7640 ( 
.A(n_7124),
.Y(n_7640)
);

INVx2_ASAP7_75t_L g7641 ( 
.A(n_7128),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_L g7642 ( 
.A(n_6952),
.B(n_12),
.Y(n_7642)
);

AOI22xp5_ASAP7_75t_L g7643 ( 
.A1(n_7275),
.A2(n_418),
.B1(n_419),
.B2(n_417),
.Y(n_7643)
);

OAI221xp5_ASAP7_75t_L g7644 ( 
.A1(n_7277),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_7644)
);

AO22x2_ASAP7_75t_L g7645 ( 
.A1(n_7178),
.A2(n_7421),
.B1(n_7044),
.B2(n_7106),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7132),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_7136),
.Y(n_7647)
);

NAND2x1p5_ASAP7_75t_L g7648 ( 
.A(n_7343),
.B(n_418),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7137),
.Y(n_7649)
);

NAND2xp5_ASAP7_75t_L g7650 ( 
.A(n_7042),
.B(n_7052),
.Y(n_7650)
);

OAI221xp5_ASAP7_75t_L g7651 ( 
.A1(n_7280),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.C(n_17),
.Y(n_7651)
);

AO22x2_ASAP7_75t_L g7652 ( 
.A1(n_7091),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_7652)
);

NAND2xp5_ASAP7_75t_L g7653 ( 
.A(n_7197),
.B(n_17),
.Y(n_7653)
);

INVx2_ASAP7_75t_L g7654 ( 
.A(n_7138),
.Y(n_7654)
);

BUFx6f_ASAP7_75t_SL g7655 ( 
.A(n_6973),
.Y(n_7655)
);

HB1xp67_ASAP7_75t_L g7656 ( 
.A(n_7014),
.Y(n_7656)
);

AOI22xp5_ASAP7_75t_L g7657 ( 
.A1(n_7424),
.A2(n_420),
.B1(n_421),
.B2(n_419),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7346),
.Y(n_7658)
);

AND2x4_ASAP7_75t_L g7659 ( 
.A(n_7397),
.B(n_7366),
.Y(n_7659)
);

AOI22xp5_ASAP7_75t_L g7660 ( 
.A1(n_6946),
.A2(n_421),
.B1(n_422),
.B2(n_420),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_6984),
.B(n_423),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7354),
.Y(n_7662)
);

NAND2xp5_ASAP7_75t_L g7663 ( 
.A(n_7210),
.B(n_18),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7358),
.Y(n_7664)
);

AND2x2_ASAP7_75t_L g7665 ( 
.A(n_7019),
.B(n_424),
.Y(n_7665)
);

NOR2xp67_ASAP7_75t_L g7666 ( 
.A(n_7152),
.B(n_18),
.Y(n_7666)
);

NAND2xp5_ASAP7_75t_L g7667 ( 
.A(n_7219),
.B(n_19),
.Y(n_7667)
);

AO22x2_ASAP7_75t_L g7668 ( 
.A1(n_7115),
.A2(n_7123),
.B1(n_7029),
.B2(n_7040),
.Y(n_7668)
);

OAI221xp5_ASAP7_75t_L g7669 ( 
.A1(n_7248),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.C(n_23),
.Y(n_7669)
);

OAI221xp5_ASAP7_75t_L g7670 ( 
.A1(n_7082),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.C(n_24),
.Y(n_7670)
);

HB1xp67_ASAP7_75t_L g7671 ( 
.A(n_7387),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7370),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7372),
.Y(n_7673)
);

BUFx8_ASAP7_75t_L g7674 ( 
.A(n_7387),
.Y(n_7674)
);

INVx1_ASAP7_75t_L g7675 ( 
.A(n_7385),
.Y(n_7675)
);

INVx2_ASAP7_75t_L g7676 ( 
.A(n_7170),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_6968),
.Y(n_7677)
);

INVx1_ASAP7_75t_L g7678 ( 
.A(n_6975),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_6985),
.Y(n_7679)
);

AO22x2_ASAP7_75t_L g7680 ( 
.A1(n_7024),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_6987),
.Y(n_7681)
);

BUFx8_ASAP7_75t_L g7682 ( 
.A(n_7018),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_6988),
.Y(n_7683)
);

INVx2_ASAP7_75t_L g7684 ( 
.A(n_7279),
.Y(n_7684)
);

BUFx3_ASAP7_75t_L g7685 ( 
.A(n_7305),
.Y(n_7685)
);

AOI22xp5_ASAP7_75t_L g7686 ( 
.A1(n_6939),
.A2(n_426),
.B1(n_427),
.B2(n_425),
.Y(n_7686)
);

OAI221xp5_ASAP7_75t_L g7687 ( 
.A1(n_7269),
.A2(n_7317),
.B1(n_7216),
.B2(n_7048),
.C(n_7050),
.Y(n_7687)
);

NAND2xp5_ASAP7_75t_L g7688 ( 
.A(n_7227),
.B(n_24),
.Y(n_7688)
);

NAND2x1p5_ASAP7_75t_L g7689 ( 
.A(n_7038),
.B(n_425),
.Y(n_7689)
);

BUFx8_ASAP7_75t_L g7690 ( 
.A(n_7064),
.Y(n_7690)
);

AND2x4_ASAP7_75t_L g7691 ( 
.A(n_7156),
.B(n_426),
.Y(n_7691)
);

CKINVDCx11_ASAP7_75t_R g7692 ( 
.A(n_7305),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_6990),
.Y(n_7693)
);

AO22x2_ASAP7_75t_L g7694 ( 
.A1(n_7303),
.A2(n_7316),
.B1(n_7309),
.B2(n_7207),
.Y(n_7694)
);

INVxp67_ASAP7_75t_L g7695 ( 
.A(n_7266),
.Y(n_7695)
);

AND2x4_ASAP7_75t_L g7696 ( 
.A(n_7335),
.B(n_427),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_6994),
.Y(n_7697)
);

INVx1_ASAP7_75t_L g7698 ( 
.A(n_6995),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_6996),
.Y(n_7699)
);

INVx2_ASAP7_75t_L g7700 ( 
.A(n_7369),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_7000),
.Y(n_7701)
);

AO22x2_ASAP7_75t_L g7702 ( 
.A1(n_7209),
.A2(n_7298),
.B1(n_7286),
.B2(n_7211),
.Y(n_7702)
);

AO22x2_ASAP7_75t_L g7703 ( 
.A1(n_7205),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_7703)
);

NAND2xp5_ASAP7_75t_L g7704 ( 
.A(n_7230),
.B(n_25),
.Y(n_7704)
);

AOI22xp5_ASAP7_75t_L g7705 ( 
.A1(n_6989),
.A2(n_429),
.B1(n_430),
.B2(n_428),
.Y(n_7705)
);

INVxp67_ASAP7_75t_SL g7706 ( 
.A(n_7201),
.Y(n_7706)
);

INVxp67_ASAP7_75t_L g7707 ( 
.A(n_7289),
.Y(n_7707)
);

AO22x2_ASAP7_75t_L g7708 ( 
.A1(n_7258),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_7708)
);

NAND2xp5_ASAP7_75t_L g7709 ( 
.A(n_7236),
.B(n_26),
.Y(n_7709)
);

NAND2xp33_ASAP7_75t_L g7710 ( 
.A(n_7367),
.B(n_27),
.Y(n_7710)
);

AO22x2_ASAP7_75t_L g7711 ( 
.A1(n_7133),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7002),
.Y(n_7712)
);

AO22x2_ASAP7_75t_L g7713 ( 
.A1(n_7200),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_7003),
.Y(n_7714)
);

BUFx6f_ASAP7_75t_SL g7715 ( 
.A(n_6973),
.Y(n_7715)
);

NAND2x1p5_ASAP7_75t_L g7716 ( 
.A(n_7088),
.B(n_430),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7007),
.Y(n_7717)
);

INVx1_ASAP7_75t_L g7718 ( 
.A(n_7009),
.Y(n_7718)
);

BUFx8_ASAP7_75t_L g7719 ( 
.A(n_7089),
.Y(n_7719)
);

AO22x2_ASAP7_75t_L g7720 ( 
.A1(n_7139),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_7013),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_7015),
.Y(n_7722)
);

AND2x4_ASAP7_75t_L g7723 ( 
.A(n_7116),
.B(n_431),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7021),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_SL g7725 ( 
.A(n_7274),
.B(n_433),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_7376),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_7022),
.Y(n_7727)
);

BUFx8_ASAP7_75t_L g7728 ( 
.A(n_7129),
.Y(n_7728)
);

AOI22xp5_ASAP7_75t_L g7729 ( 
.A1(n_7125),
.A2(n_434),
.B1(n_435),
.B2(n_433),
.Y(n_7729)
);

INVx1_ASAP7_75t_L g7730 ( 
.A(n_7023),
.Y(n_7730)
);

INVxp67_ASAP7_75t_L g7731 ( 
.A(n_7235),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7026),
.Y(n_7732)
);

AND2x2_ASAP7_75t_L g7733 ( 
.A(n_7020),
.B(n_434),
.Y(n_7733)
);

INVx1_ASAP7_75t_L g7734 ( 
.A(n_7030),
.Y(n_7734)
);

NAND2xp5_ASAP7_75t_L g7735 ( 
.A(n_7242),
.B(n_30),
.Y(n_7735)
);

OAI221xp5_ASAP7_75t_L g7736 ( 
.A1(n_7046),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_7036),
.Y(n_7737)
);

AO22x2_ASAP7_75t_L g7738 ( 
.A1(n_7148),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_7738)
);

INVx1_ASAP7_75t_L g7739 ( 
.A(n_7054),
.Y(n_7739)
);

CKINVDCx11_ASAP7_75t_R g7740 ( 
.A(n_6929),
.Y(n_7740)
);

INVx1_ASAP7_75t_L g7741 ( 
.A(n_7062),
.Y(n_7741)
);

CKINVDCx5p33_ASAP7_75t_R g7742 ( 
.A(n_7229),
.Y(n_7742)
);

AO22x2_ASAP7_75t_L g7743 ( 
.A1(n_7228),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7063),
.Y(n_7744)
);

NOR2xp33_ASAP7_75t_L g7745 ( 
.A(n_7334),
.B(n_435),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_L g7746 ( 
.A(n_7244),
.B(n_35),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7065),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7066),
.Y(n_7748)
);

AO22x2_ASAP7_75t_L g7749 ( 
.A1(n_7250),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7067),
.Y(n_7750)
);

INVxp67_ASAP7_75t_L g7751 ( 
.A(n_7060),
.Y(n_7751)
);

NAND2xp5_ASAP7_75t_L g7752 ( 
.A(n_7083),
.B(n_36),
.Y(n_7752)
);

AO22x2_ASAP7_75t_L g7753 ( 
.A1(n_7371),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_7753)
);

OAI22xp5_ASAP7_75t_SL g7754 ( 
.A1(n_7180),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_7754)
);

AO22x2_ASAP7_75t_L g7755 ( 
.A1(n_7165),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_7755)
);

AND2x2_ASAP7_75t_L g7756 ( 
.A(n_7058),
.B(n_436),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7394),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_7163),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7184),
.Y(n_7759)
);

NAND2x1p5_ASAP7_75t_L g7760 ( 
.A(n_7333),
.B(n_436),
.Y(n_7760)
);

NAND2xp5_ASAP7_75t_L g7761 ( 
.A(n_7300),
.B(n_42),
.Y(n_7761)
);

AOI22xp33_ASAP7_75t_L g7762 ( 
.A1(n_7415),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7027),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7181),
.Y(n_7764)
);

AOI22xp5_ASAP7_75t_L g7765 ( 
.A1(n_7158),
.A2(n_439),
.B1(n_440),
.B2(n_437),
.Y(n_7765)
);

AO22x2_ASAP7_75t_L g7766 ( 
.A1(n_7336),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_7766)
);

CKINVDCx20_ASAP7_75t_R g7767 ( 
.A(n_7103),
.Y(n_7767)
);

CKINVDCx5p33_ASAP7_75t_R g7768 ( 
.A(n_7154),
.Y(n_7768)
);

AO22x2_ASAP7_75t_L g7769 ( 
.A1(n_7080),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_7769)
);

INVx2_ASAP7_75t_L g7770 ( 
.A(n_7182),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7190),
.Y(n_7771)
);

NAND2xp5_ASAP7_75t_L g7772 ( 
.A(n_7287),
.B(n_7290),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7194),
.Y(n_7773)
);

AO22x2_ASAP7_75t_L g7774 ( 
.A1(n_7381),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_7774)
);

AO22x2_ASAP7_75t_L g7775 ( 
.A1(n_7382),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_7246),
.Y(n_7776)
);

BUFx8_ASAP7_75t_L g7777 ( 
.A(n_7157),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7214),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7310),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7312),
.Y(n_7780)
);

AND2x4_ASAP7_75t_L g7781 ( 
.A(n_7393),
.B(n_7340),
.Y(n_7781)
);

INVx8_ASAP7_75t_L g7782 ( 
.A(n_7398),
.Y(n_7782)
);

NAND2x1p5_ASAP7_75t_L g7783 ( 
.A(n_7403),
.B(n_437),
.Y(n_7783)
);

INVx2_ASAP7_75t_L g7784 ( 
.A(n_7264),
.Y(n_7784)
);

BUFx2_ASAP7_75t_L g7785 ( 
.A(n_7160),
.Y(n_7785)
);

AO22x2_ASAP7_75t_L g7786 ( 
.A1(n_7081),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_7786)
);

INVxp67_ASAP7_75t_L g7787 ( 
.A(n_7143),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7001),
.Y(n_7788)
);

OAI221xp5_ASAP7_75t_L g7789 ( 
.A1(n_7051),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_7789)
);

NAND2x1p5_ASAP7_75t_L g7790 ( 
.A(n_6945),
.B(n_440),
.Y(n_7790)
);

NAND2xp5_ASAP7_75t_L g7791 ( 
.A(n_7291),
.B(n_48),
.Y(n_7791)
);

OAI221xp5_ASAP7_75t_L g7792 ( 
.A1(n_7238),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.C(n_52),
.Y(n_7792)
);

OAI221xp5_ASAP7_75t_L g7793 ( 
.A1(n_7401),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_7793)
);

INVx2_ASAP7_75t_L g7794 ( 
.A(n_7261),
.Y(n_7794)
);

AO22x2_ASAP7_75t_L g7795 ( 
.A1(n_7183),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_7795)
);

INVx2_ASAP7_75t_SL g7796 ( 
.A(n_7154),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_L g7797 ( 
.A(n_7070),
.B(n_53),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7285),
.Y(n_7798)
);

AO22x2_ASAP7_75t_L g7799 ( 
.A1(n_7314),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_7799)
);

INVx2_ASAP7_75t_SL g7800 ( 
.A(n_7215),
.Y(n_7800)
);

NAND2xp5_ASAP7_75t_L g7801 ( 
.A(n_7101),
.B(n_55),
.Y(n_7801)
);

AOI22xp5_ASAP7_75t_L g7802 ( 
.A1(n_7193),
.A2(n_7288),
.B1(n_7260),
.B2(n_7072),
.Y(n_7802)
);

INVx1_ASAP7_75t_L g7803 ( 
.A(n_7388),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7390),
.Y(n_7804)
);

INVx1_ASAP7_75t_L g7805 ( 
.A(n_7411),
.Y(n_7805)
);

BUFx8_ASAP7_75t_L g7806 ( 
.A(n_6979),
.Y(n_7806)
);

INVx2_ASAP7_75t_L g7807 ( 
.A(n_7278),
.Y(n_7807)
);

INVx1_ASAP7_75t_L g7808 ( 
.A(n_7417),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_7267),
.Y(n_7809)
);

BUFx8_ASAP7_75t_L g7810 ( 
.A(n_7319),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_7268),
.Y(n_7811)
);

BUFx3_ASAP7_75t_L g7812 ( 
.A(n_7398),
.Y(n_7812)
);

AOI22xp5_ASAP7_75t_L g7813 ( 
.A1(n_7090),
.A2(n_7153),
.B1(n_7386),
.B2(n_7295),
.Y(n_7813)
);

INVx2_ASAP7_75t_L g7814 ( 
.A(n_7215),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7257),
.Y(n_7815)
);

AO22x2_ASAP7_75t_L g7816 ( 
.A1(n_7320),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_7816)
);

INVx2_ASAP7_75t_L g7817 ( 
.A(n_7359),
.Y(n_7817)
);

AO22x2_ASAP7_75t_L g7818 ( 
.A1(n_7324),
.A2(n_7330),
.B1(n_7344),
.B2(n_7331),
.Y(n_7818)
);

AO22x2_ASAP7_75t_L g7819 ( 
.A1(n_7347),
.A2(n_7353),
.B1(n_7364),
.B2(n_7355),
.Y(n_7819)
);

OR2x6_ASAP7_75t_L g7820 ( 
.A(n_7110),
.B(n_7199),
.Y(n_7820)
);

NAND2xp5_ASAP7_75t_L g7821 ( 
.A(n_7168),
.B(n_57),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_7166),
.Y(n_7822)
);

INVx1_ASAP7_75t_L g7823 ( 
.A(n_7391),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_7392),
.Y(n_7824)
);

AND2x6_ASAP7_75t_L g7825 ( 
.A(n_7338),
.B(n_57),
.Y(n_7825)
);

INVx1_ASAP7_75t_L g7826 ( 
.A(n_7237),
.Y(n_7826)
);

AOI22xp5_ASAP7_75t_L g7827 ( 
.A1(n_7100),
.A2(n_7294),
.B1(n_7240),
.B2(n_7149),
.Y(n_7827)
);

INVx4_ASAP7_75t_L g7828 ( 
.A(n_7419),
.Y(n_7828)
);

INVx1_ASAP7_75t_L g7829 ( 
.A(n_7075),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7384),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7407),
.Y(n_7831)
);

INVx1_ASAP7_75t_L g7832 ( 
.A(n_7360),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7218),
.Y(n_7833)
);

CKINVDCx14_ASAP7_75t_R g7834 ( 
.A(n_7308),
.Y(n_7834)
);

AO22x2_ASAP7_75t_L g7835 ( 
.A1(n_7204),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_L g7836 ( 
.A(n_7134),
.B(n_58),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7273),
.Y(n_7837)
);

NOR2xp33_ASAP7_75t_L g7838 ( 
.A(n_7150),
.B(n_441),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7348),
.Y(n_7839)
);

INVxp33_ASAP7_75t_L g7840 ( 
.A(n_7127),
.Y(n_7840)
);

AND2x4_ASAP7_75t_L g7841 ( 
.A(n_7056),
.B(n_442),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_7378),
.Y(n_7842)
);

INVx1_ASAP7_75t_SL g7843 ( 
.A(n_6965),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_7047),
.Y(n_7844)
);

AO22x2_ASAP7_75t_L g7845 ( 
.A1(n_7053),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_7845)
);

NAND2xp33_ASAP7_75t_L g7846 ( 
.A(n_7176),
.B(n_59),
.Y(n_7846)
);

INVx2_ASAP7_75t_L g7847 ( 
.A(n_7251),
.Y(n_7847)
);

AND2x4_ASAP7_75t_L g7848 ( 
.A(n_7012),
.B(n_442),
.Y(n_7848)
);

AND2x2_ASAP7_75t_L g7849 ( 
.A(n_7302),
.B(n_443),
.Y(n_7849)
);

BUFx8_ASAP7_75t_L g7850 ( 
.A(n_7408),
.Y(n_7850)
);

AO22x2_ASAP7_75t_L g7851 ( 
.A1(n_7301),
.A2(n_7169),
.B1(n_7188),
.B2(n_7187),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7379),
.Y(n_7852)
);

AO22x2_ASAP7_75t_L g7853 ( 
.A1(n_7326),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_7350),
.Y(n_7854)
);

AOI22xp5_ASAP7_75t_L g7855 ( 
.A1(n_7016),
.A2(n_444),
.B1(n_445),
.B2(n_443),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7365),
.Y(n_7856)
);

AND2x2_ASAP7_75t_L g7857 ( 
.A(n_7419),
.B(n_444),
.Y(n_7857)
);

BUFx6f_ASAP7_75t_L g7858 ( 
.A(n_7368),
.Y(n_7858)
);

INVx2_ASAP7_75t_L g7859 ( 
.A(n_7262),
.Y(n_7859)
);

NAND2xp5_ASAP7_75t_L g7860 ( 
.A(n_7028),
.B(n_61),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7374),
.Y(n_7861)
);

INVx4_ASAP7_75t_L g7862 ( 
.A(n_7112),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_7380),
.Y(n_7863)
);

INVx1_ASAP7_75t_L g7864 ( 
.A(n_7416),
.Y(n_7864)
);

INVx2_ASAP7_75t_L g7865 ( 
.A(n_7282),
.Y(n_7865)
);

AO22x2_ASAP7_75t_L g7866 ( 
.A1(n_7383),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_7866)
);

NAND2x1p5_ASAP7_75t_L g7867 ( 
.A(n_7032),
.B(n_446),
.Y(n_7867)
);

NAND2xp5_ASAP7_75t_L g7868 ( 
.A(n_7206),
.B(n_63),
.Y(n_7868)
);

A2O1A1Ixp33_ASAP7_75t_L g7869 ( 
.A1(n_7297),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_7869)
);

AND2x4_ASAP7_75t_L g7870 ( 
.A(n_7321),
.B(n_446),
.Y(n_7870)
);

AO22x2_ASAP7_75t_L g7871 ( 
.A1(n_7400),
.A2(n_7404),
.B1(n_7425),
.B2(n_7396),
.Y(n_7871)
);

NAND2xp5_ASAP7_75t_L g7872 ( 
.A(n_7332),
.B(n_64),
.Y(n_7872)
);

NAND2xp5_ASAP7_75t_L g7873 ( 
.A(n_7413),
.B(n_65),
.Y(n_7873)
);

OR2x2_ASAP7_75t_L g7874 ( 
.A(n_7092),
.B(n_66),
.Y(n_7874)
);

NAND2xp5_ASAP7_75t_L g7875 ( 
.A(n_7179),
.B(n_66),
.Y(n_7875)
);

OAI22xp5_ASAP7_75t_L g7876 ( 
.A1(n_7179),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_7876)
);

CKINVDCx5p33_ASAP7_75t_R g7877 ( 
.A(n_6954),
.Y(n_7877)
);

CKINVDCx11_ASAP7_75t_R g7878 ( 
.A(n_7162),
.Y(n_7878)
);

INVx2_ASAP7_75t_L g7879 ( 
.A(n_6932),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_6932),
.Y(n_7880)
);

INVx2_ASAP7_75t_L g7881 ( 
.A(n_6932),
.Y(n_7881)
);

INVx1_ASAP7_75t_SL g7882 ( 
.A(n_6972),
.Y(n_7882)
);

CKINVDCx16_ASAP7_75t_R g7883 ( 
.A(n_7162),
.Y(n_7883)
);

INVxp67_ASAP7_75t_L g7884 ( 
.A(n_7092),
.Y(n_7884)
);

AND2x4_ASAP7_75t_L g7885 ( 
.A(n_7185),
.B(n_447),
.Y(n_7885)
);

OAI221xp5_ASAP7_75t_L g7886 ( 
.A1(n_7179),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_7886)
);

INVx2_ASAP7_75t_SL g7887 ( 
.A(n_7406),
.Y(n_7887)
);

INVx2_ASAP7_75t_L g7888 ( 
.A(n_6932),
.Y(n_7888)
);

AOI22xp5_ASAP7_75t_L g7889 ( 
.A1(n_7017),
.A2(n_449),
.B1(n_450),
.B2(n_448),
.Y(n_7889)
);

AND2x4_ASAP7_75t_L g7890 ( 
.A(n_7185),
.B(n_450),
.Y(n_7890)
);

AO22x2_ASAP7_75t_L g7891 ( 
.A1(n_6930),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_7891)
);

AND2x2_ASAP7_75t_L g7892 ( 
.A(n_7043),
.B(n_451),
.Y(n_7892)
);

NOR2xp33_ASAP7_75t_L g7893 ( 
.A(n_7179),
.B(n_452),
.Y(n_7893)
);

INVx2_ASAP7_75t_L g7894 ( 
.A(n_6932),
.Y(n_7894)
);

AOI22xp5_ASAP7_75t_L g7895 ( 
.A1(n_7017),
.A2(n_453),
.B1(n_454),
.B2(n_452),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_6932),
.Y(n_7896)
);

NAND2xp5_ASAP7_75t_L g7897 ( 
.A(n_7179),
.B(n_67),
.Y(n_7897)
);

AND2x4_ASAP7_75t_L g7898 ( 
.A(n_7185),
.B(n_453),
.Y(n_7898)
);

AND2x4_ASAP7_75t_L g7899 ( 
.A(n_7185),
.B(n_455),
.Y(n_7899)
);

NAND2xp5_ASAP7_75t_L g7900 ( 
.A(n_7179),
.B(n_68),
.Y(n_7900)
);

AO22x2_ASAP7_75t_L g7901 ( 
.A1(n_6930),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_7901)
);

NAND2xp5_ASAP7_75t_L g7902 ( 
.A(n_7179),
.B(n_70),
.Y(n_7902)
);

AOI22xp5_ASAP7_75t_L g7903 ( 
.A1(n_7017),
.A2(n_456),
.B1(n_457),
.B2(n_455),
.Y(n_7903)
);

AO22x2_ASAP7_75t_L g7904 ( 
.A1(n_6930),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_7904)
);

NAND2xp5_ASAP7_75t_L g7905 ( 
.A(n_7179),
.B(n_72),
.Y(n_7905)
);

HB1xp67_ASAP7_75t_L g7906 ( 
.A(n_7092),
.Y(n_7906)
);

INVx1_ASAP7_75t_L g7907 ( 
.A(n_6932),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_6932),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_6932),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_6932),
.Y(n_7910)
);

INVx1_ASAP7_75t_L g7911 ( 
.A(n_6932),
.Y(n_7911)
);

OAI221xp5_ASAP7_75t_L g7912 ( 
.A1(n_7179),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_7912)
);

INVxp67_ASAP7_75t_L g7913 ( 
.A(n_7092),
.Y(n_7913)
);

AND2x6_ASAP7_75t_L g7914 ( 
.A(n_7272),
.B(n_73),
.Y(n_7914)
);

INVx2_ASAP7_75t_L g7915 ( 
.A(n_6932),
.Y(n_7915)
);

AND2x4_ASAP7_75t_L g7916 ( 
.A(n_7185),
.B(n_456),
.Y(n_7916)
);

NAND2xp5_ASAP7_75t_L g7917 ( 
.A(n_7179),
.B(n_75),
.Y(n_7917)
);

AO22x2_ASAP7_75t_L g7918 ( 
.A1(n_6930),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_7918)
);

OAI22xp5_ASAP7_75t_L g7919 ( 
.A1(n_7179),
.A2(n_458),
.B1(n_459),
.B2(n_457),
.Y(n_7919)
);

NAND2xp5_ASAP7_75t_L g7920 ( 
.A(n_7179),
.B(n_76),
.Y(n_7920)
);

AOI22xp5_ASAP7_75t_L g7921 ( 
.A1(n_7017),
.A2(n_460),
.B1(n_461),
.B2(n_459),
.Y(n_7921)
);

AO22x2_ASAP7_75t_L g7922 ( 
.A1(n_6930),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_6932),
.Y(n_7923)
);

NOR2xp33_ASAP7_75t_L g7924 ( 
.A(n_7179),
.B(n_461),
.Y(n_7924)
);

BUFx8_ASAP7_75t_L g7925 ( 
.A(n_6924),
.Y(n_7925)
);

NAND2xp5_ASAP7_75t_L g7926 ( 
.A(n_7507),
.B(n_7613),
.Y(n_7926)
);

NOR2xp33_ASAP7_75t_L g7927 ( 
.A(n_7557),
.B(n_462),
.Y(n_7927)
);

BUFx6f_ASAP7_75t_L g7928 ( 
.A(n_7499),
.Y(n_7928)
);

BUFx3_ASAP7_75t_L g7929 ( 
.A(n_7587),
.Y(n_7929)
);

INVx2_ASAP7_75t_L g7930 ( 
.A(n_7428),
.Y(n_7930)
);

O2A1O1Ixp33_ASAP7_75t_L g7931 ( 
.A1(n_7513),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_7931)
);

NOR2xp33_ASAP7_75t_L g7932 ( 
.A(n_7618),
.B(n_462),
.Y(n_7932)
);

AOI21xp5_ASAP7_75t_L g7933 ( 
.A1(n_7461),
.A2(n_464),
.B(n_463),
.Y(n_7933)
);

CKINVDCx10_ASAP7_75t_R g7934 ( 
.A(n_7883),
.Y(n_7934)
);

NAND2xp5_ASAP7_75t_L g7935 ( 
.A(n_7464),
.B(n_7465),
.Y(n_7935)
);

AOI21xp5_ASAP7_75t_L g7936 ( 
.A1(n_7650),
.A2(n_466),
.B(n_465),
.Y(n_7936)
);

AOI21xp5_ASAP7_75t_L g7937 ( 
.A1(n_7772),
.A2(n_467),
.B(n_465),
.Y(n_7937)
);

OAI22xp5_ASAP7_75t_L g7938 ( 
.A1(n_7600),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_7938)
);

NAND2xp5_ASAP7_75t_SL g7939 ( 
.A(n_7541),
.B(n_468),
.Y(n_7939)
);

AOI21xp5_ASAP7_75t_L g7940 ( 
.A1(n_7687),
.A2(n_7811),
.B(n_7784),
.Y(n_7940)
);

NOR2xp67_ASAP7_75t_L g7941 ( 
.A(n_7862),
.B(n_80),
.Y(n_7941)
);

AOI21x1_ASAP7_75t_L g7942 ( 
.A1(n_7818),
.A2(n_7819),
.B(n_7508),
.Y(n_7942)
);

NAND2xp5_ASAP7_75t_L g7943 ( 
.A(n_7468),
.B(n_81),
.Y(n_7943)
);

AOI21xp5_ASAP7_75t_L g7944 ( 
.A1(n_7794),
.A2(n_470),
.B(n_469),
.Y(n_7944)
);

NAND2xp5_ASAP7_75t_L g7945 ( 
.A(n_7476),
.B(n_7807),
.Y(n_7945)
);

NAND2xp5_ASAP7_75t_L g7946 ( 
.A(n_7677),
.B(n_81),
.Y(n_7946)
);

AOI21x1_ASAP7_75t_L g7947 ( 
.A1(n_7444),
.A2(n_82),
.B(n_83),
.Y(n_7947)
);

OR2x6_ASAP7_75t_L g7948 ( 
.A(n_7782),
.B(n_7462),
.Y(n_7948)
);

NAND2x1_ASAP7_75t_L g7949 ( 
.A(n_7570),
.B(n_471),
.Y(n_7949)
);

NAND2xp5_ASAP7_75t_L g7950 ( 
.A(n_7678),
.B(n_7679),
.Y(n_7950)
);

AOI21xp5_ASAP7_75t_L g7951 ( 
.A1(n_7504),
.A2(n_472),
.B(n_471),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7452),
.Y(n_7952)
);

NOR2xp33_ASAP7_75t_L g7953 ( 
.A(n_7787),
.B(n_472),
.Y(n_7953)
);

AOI21xp5_ASAP7_75t_L g7954 ( 
.A1(n_7435),
.A2(n_475),
.B(n_473),
.Y(n_7954)
);

O2A1O1Ixp5_ASAP7_75t_L g7955 ( 
.A1(n_7893),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_7955)
);

INVx2_ASAP7_75t_L g7956 ( 
.A(n_7466),
.Y(n_7956)
);

NAND2xp5_ASAP7_75t_SL g7957 ( 
.A(n_7492),
.B(n_473),
.Y(n_7957)
);

NAND2xp5_ASAP7_75t_L g7958 ( 
.A(n_7681),
.B(n_82),
.Y(n_7958)
);

NOR2xp33_ASAP7_75t_L g7959 ( 
.A(n_7683),
.B(n_475),
.Y(n_7959)
);

INVx3_ASAP7_75t_L g7960 ( 
.A(n_7450),
.Y(n_7960)
);

AOI21x1_ASAP7_75t_L g7961 ( 
.A1(n_7451),
.A2(n_83),
.B(n_84),
.Y(n_7961)
);

AOI21xp5_ASAP7_75t_L g7962 ( 
.A1(n_7628),
.A2(n_477),
.B(n_476),
.Y(n_7962)
);

BUFx6f_ASAP7_75t_L g7963 ( 
.A(n_7692),
.Y(n_7963)
);

NOR2x1_ASAP7_75t_L g7964 ( 
.A(n_7429),
.B(n_476),
.Y(n_7964)
);

NAND2xp5_ASAP7_75t_L g7965 ( 
.A(n_7693),
.B(n_84),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_7879),
.Y(n_7966)
);

INVx1_ASAP7_75t_SL g7967 ( 
.A(n_7882),
.Y(n_7967)
);

INVx2_ASAP7_75t_L g7968 ( 
.A(n_7881),
.Y(n_7968)
);

A2O1A1Ixp33_ASAP7_75t_L g7969 ( 
.A1(n_7924),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_7969)
);

OAI21xp5_ASAP7_75t_L g7970 ( 
.A1(n_7615),
.A2(n_85),
.B(n_86),
.Y(n_7970)
);

INVx3_ASAP7_75t_L g7971 ( 
.A(n_7445),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_7888),
.Y(n_7972)
);

AOI22xp5_ASAP7_75t_L g7973 ( 
.A1(n_7802),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_7973)
);

AOI22xp5_ASAP7_75t_L g7974 ( 
.A1(n_7457),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_7974)
);

CKINVDCx10_ASAP7_75t_R g7975 ( 
.A(n_7655),
.Y(n_7975)
);

NAND2xp5_ASAP7_75t_SL g7976 ( 
.A(n_7827),
.B(n_477),
.Y(n_7976)
);

AOI21xp5_ASAP7_75t_L g7977 ( 
.A1(n_7629),
.A2(n_479),
.B(n_478),
.Y(n_7977)
);

NOR2xp33_ASAP7_75t_L g7978 ( 
.A(n_7697),
.B(n_478),
.Y(n_7978)
);

NAND2xp5_ASAP7_75t_SL g7979 ( 
.A(n_7495),
.B(n_479),
.Y(n_7979)
);

AOI21xp5_ASAP7_75t_L g7980 ( 
.A1(n_7635),
.A2(n_481),
.B(n_480),
.Y(n_7980)
);

A2O1A1Ixp33_ASAP7_75t_L g7981 ( 
.A1(n_7813),
.A2(n_91),
.B(n_88),
.C(n_90),
.Y(n_7981)
);

NAND2xp5_ASAP7_75t_L g7982 ( 
.A(n_7698),
.B(n_90),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_7894),
.Y(n_7983)
);

O2A1O1Ixp33_ASAP7_75t_L g7984 ( 
.A1(n_7821),
.A2(n_7846),
.B(n_7897),
.C(n_7875),
.Y(n_7984)
);

AOI21xp5_ASAP7_75t_L g7985 ( 
.A1(n_7636),
.A2(n_482),
.B(n_481),
.Y(n_7985)
);

INVx2_ASAP7_75t_L g7986 ( 
.A(n_7915),
.Y(n_7986)
);

AOI21xp5_ASAP7_75t_L g7987 ( 
.A1(n_7637),
.A2(n_483),
.B(n_482),
.Y(n_7987)
);

NAND2x1_ASAP7_75t_L g7988 ( 
.A(n_7572),
.B(n_485),
.Y(n_7988)
);

NAND2xp5_ASAP7_75t_L g7989 ( 
.A(n_7699),
.B(n_91),
.Y(n_7989)
);

A2O1A1Ixp33_ASAP7_75t_L g7990 ( 
.A1(n_7527),
.A2(n_7531),
.B(n_7832),
.C(n_7900),
.Y(n_7990)
);

INVx1_ASAP7_75t_L g7991 ( 
.A(n_7427),
.Y(n_7991)
);

BUFx3_ASAP7_75t_L g7992 ( 
.A(n_7605),
.Y(n_7992)
);

NOR2x1_ASAP7_75t_L g7993 ( 
.A(n_7843),
.B(n_485),
.Y(n_7993)
);

CKINVDCx10_ASAP7_75t_R g7994 ( 
.A(n_7715),
.Y(n_7994)
);

BUFx2_ASAP7_75t_L g7995 ( 
.A(n_7463),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_L g7996 ( 
.A(n_7701),
.B(n_91),
.Y(n_7996)
);

INVx2_ASAP7_75t_L g7997 ( 
.A(n_7524),
.Y(n_7997)
);

AOI21xp5_ASAP7_75t_L g7998 ( 
.A1(n_7638),
.A2(n_487),
.B(n_486),
.Y(n_7998)
);

NOR2xp33_ASAP7_75t_L g7999 ( 
.A(n_7712),
.B(n_486),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_L g8000 ( 
.A(n_7714),
.B(n_93),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7717),
.B(n_93),
.Y(n_8001)
);

INVx1_ASAP7_75t_L g8002 ( 
.A(n_7431),
.Y(n_8002)
);

AOI21xp5_ASAP7_75t_L g8003 ( 
.A1(n_7646),
.A2(n_488),
.B(n_487),
.Y(n_8003)
);

INVx2_ASAP7_75t_L g8004 ( 
.A(n_7497),
.Y(n_8004)
);

AOI22xp5_ASAP7_75t_L g8005 ( 
.A1(n_7668),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_8005)
);

AOI21xp5_ASAP7_75t_L g8006 ( 
.A1(n_7647),
.A2(n_7649),
.B(n_7798),
.Y(n_8006)
);

AND2x4_ASAP7_75t_L g8007 ( 
.A(n_7472),
.B(n_489),
.Y(n_8007)
);

AOI21xp5_ASAP7_75t_L g8008 ( 
.A1(n_7803),
.A2(n_490),
.B(n_489),
.Y(n_8008)
);

A2O1A1Ixp33_ASAP7_75t_L g8009 ( 
.A1(n_7902),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_8009)
);

AOI21xp5_ASAP7_75t_L g8010 ( 
.A1(n_7804),
.A2(n_492),
.B(n_491),
.Y(n_8010)
);

NAND2xp5_ASAP7_75t_L g8011 ( 
.A(n_7718),
.B(n_94),
.Y(n_8011)
);

NAND2xp5_ASAP7_75t_L g8012 ( 
.A(n_7721),
.B(n_95),
.Y(n_8012)
);

AOI21xp5_ASAP7_75t_L g8013 ( 
.A1(n_7764),
.A2(n_7773),
.B(n_7771),
.Y(n_8013)
);

AOI22xp5_ASAP7_75t_L g8014 ( 
.A1(n_7851),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_8014)
);

A2O1A1Ixp33_ASAP7_75t_L g8015 ( 
.A1(n_7905),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_8015)
);

NOR2xp33_ASAP7_75t_L g8016 ( 
.A(n_7722),
.B(n_491),
.Y(n_8016)
);

INVx1_ASAP7_75t_L g8017 ( 
.A(n_7433),
.Y(n_8017)
);

NAND2xp5_ASAP7_75t_SL g8018 ( 
.A(n_7516),
.B(n_492),
.Y(n_8018)
);

INVx3_ASAP7_75t_L g8019 ( 
.A(n_7447),
.Y(n_8019)
);

O2A1O1Ixp33_ASAP7_75t_L g8020 ( 
.A1(n_7917),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_8020)
);

INVx3_ASAP7_75t_L g8021 ( 
.A(n_7539),
.Y(n_8021)
);

INVx3_ASAP7_75t_L g8022 ( 
.A(n_7505),
.Y(n_8022)
);

AO21x2_ASAP7_75t_L g8023 ( 
.A1(n_7761),
.A2(n_99),
.B(n_100),
.Y(n_8023)
);

NAND2xp5_ASAP7_75t_L g8024 ( 
.A(n_7724),
.B(n_101),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7436),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7520),
.Y(n_8026)
);

NAND2xp5_ASAP7_75t_L g8027 ( 
.A(n_7727),
.B(n_101),
.Y(n_8027)
);

NOR2xp33_ASAP7_75t_SL g8028 ( 
.A(n_7471),
.B(n_101),
.Y(n_8028)
);

AOI21x1_ASAP7_75t_L g8029 ( 
.A1(n_7694),
.A2(n_102),
.B(n_103),
.Y(n_8029)
);

INVx1_ASAP7_75t_L g8030 ( 
.A(n_7440),
.Y(n_8030)
);

AO21x1_ASAP7_75t_L g8031 ( 
.A1(n_7839),
.A2(n_494),
.B(n_493),
.Y(n_8031)
);

AOI21xp5_ASAP7_75t_L g8032 ( 
.A1(n_7730),
.A2(n_495),
.B(n_494),
.Y(n_8032)
);

OAI21xp5_ASAP7_75t_L g8033 ( 
.A1(n_7561),
.A2(n_102),
.B(n_103),
.Y(n_8033)
);

AOI21xp5_ASAP7_75t_L g8034 ( 
.A1(n_7732),
.A2(n_496),
.B(n_495),
.Y(n_8034)
);

AOI21xp5_ASAP7_75t_L g8035 ( 
.A1(n_7734),
.A2(n_498),
.B(n_497),
.Y(n_8035)
);

OAI22xp5_ASAP7_75t_L g8036 ( 
.A1(n_7707),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_8036)
);

NOR2xp67_ASAP7_75t_L g8037 ( 
.A(n_7533),
.B(n_104),
.Y(n_8037)
);

OAI21xp5_ASAP7_75t_L g8038 ( 
.A1(n_7619),
.A2(n_104),
.B(n_105),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_L g8039 ( 
.A(n_7737),
.B(n_105),
.Y(n_8039)
);

AOI21xp5_ASAP7_75t_L g8040 ( 
.A1(n_7739),
.A2(n_498),
.B(n_497),
.Y(n_8040)
);

A2O1A1Ixp33_ASAP7_75t_L g8041 ( 
.A1(n_7920),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_8041)
);

NOR3xp33_ASAP7_75t_L g8042 ( 
.A(n_7576),
.B(n_106),
.C(n_107),
.Y(n_8042)
);

O2A1O1Ixp33_ASAP7_75t_L g8043 ( 
.A1(n_7836),
.A2(n_109),
.B(n_106),
.C(n_108),
.Y(n_8043)
);

AOI21xp5_ASAP7_75t_L g8044 ( 
.A1(n_7741),
.A2(n_500),
.B(n_499),
.Y(n_8044)
);

AOI22xp5_ASAP7_75t_SL g8045 ( 
.A1(n_7892),
.A2(n_111),
.B1(n_108),
.B2(n_110),
.Y(n_8045)
);

BUFx6f_ASAP7_75t_L g8046 ( 
.A(n_7499),
.Y(n_8046)
);

NAND2xp5_ASAP7_75t_L g8047 ( 
.A(n_7744),
.B(n_110),
.Y(n_8047)
);

NAND2xp5_ASAP7_75t_SL g8048 ( 
.A(n_7747),
.B(n_500),
.Y(n_8048)
);

O2A1O1Ixp33_ASAP7_75t_L g8049 ( 
.A1(n_7725),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_8049)
);

NAND2xp5_ASAP7_75t_L g8050 ( 
.A(n_7748),
.B(n_111),
.Y(n_8050)
);

NAND2xp5_ASAP7_75t_L g8051 ( 
.A(n_7750),
.B(n_112),
.Y(n_8051)
);

AOI21xp5_ASAP7_75t_L g8052 ( 
.A1(n_7776),
.A2(n_502),
.B(n_501),
.Y(n_8052)
);

NAND2xp5_ASAP7_75t_L g8053 ( 
.A(n_7639),
.B(n_7640),
.Y(n_8053)
);

O2A1O1Ixp33_ASAP7_75t_L g8054 ( 
.A1(n_7710),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_8054)
);

NAND2xp5_ASAP7_75t_L g8055 ( 
.A(n_7641),
.B(n_113),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_7528),
.Y(n_8056)
);

NAND2xp5_ASAP7_75t_L g8057 ( 
.A(n_7654),
.B(n_114),
.Y(n_8057)
);

INVx2_ASAP7_75t_L g8058 ( 
.A(n_7529),
.Y(n_8058)
);

NOR2xp33_ASAP7_75t_L g8059 ( 
.A(n_7840),
.B(n_501),
.Y(n_8059)
);

NAND2xp5_ASAP7_75t_L g8060 ( 
.A(n_7545),
.B(n_114),
.Y(n_8060)
);

NAND2xp5_ASAP7_75t_SL g8061 ( 
.A(n_7437),
.B(n_503),
.Y(n_8061)
);

AND2x2_ASAP7_75t_L g8062 ( 
.A(n_7830),
.B(n_115),
.Y(n_8062)
);

NAND2xp5_ASAP7_75t_L g8063 ( 
.A(n_7815),
.B(n_115),
.Y(n_8063)
);

INVx3_ASAP7_75t_L g8064 ( 
.A(n_7485),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_L g8065 ( 
.A(n_7822),
.B(n_7831),
.Y(n_8065)
);

AOI21xp5_ASAP7_75t_L g8066 ( 
.A1(n_7759),
.A2(n_504),
.B(n_503),
.Y(n_8066)
);

NAND2xp5_ASAP7_75t_L g8067 ( 
.A(n_7770),
.B(n_116),
.Y(n_8067)
);

NOR2xp33_ASAP7_75t_L g8068 ( 
.A(n_7842),
.B(n_504),
.Y(n_8068)
);

NAND2xp5_ASAP7_75t_L g8069 ( 
.A(n_7577),
.B(n_116),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_L g8070 ( 
.A(n_7554),
.B(n_7751),
.Y(n_8070)
);

AOI21xp5_ASAP7_75t_L g8071 ( 
.A1(n_7864),
.A2(n_506),
.B(n_505),
.Y(n_8071)
);

INVx1_ASAP7_75t_L g8072 ( 
.A(n_7441),
.Y(n_8072)
);

AOI21xp5_ASAP7_75t_L g8073 ( 
.A1(n_7833),
.A2(n_507),
.B(n_505),
.Y(n_8073)
);

O2A1O1Ixp33_ASAP7_75t_L g8074 ( 
.A1(n_7838),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_8074)
);

AOI22x1_ASAP7_75t_L g8075 ( 
.A1(n_7645),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_8075)
);

NAND2xp5_ASAP7_75t_L g8076 ( 
.A(n_7695),
.B(n_117),
.Y(n_8076)
);

AOI21xp5_ASAP7_75t_L g8077 ( 
.A1(n_7837),
.A2(n_508),
.B(n_507),
.Y(n_8077)
);

INVx2_ASAP7_75t_L g8078 ( 
.A(n_7525),
.Y(n_8078)
);

OAI21xp33_ASAP7_75t_L g8079 ( 
.A1(n_7564),
.A2(n_118),
.B(n_119),
.Y(n_8079)
);

AOI21xp5_ASAP7_75t_L g8080 ( 
.A1(n_7823),
.A2(n_509),
.B(n_508),
.Y(n_8080)
);

NAND3xp33_ASAP7_75t_L g8081 ( 
.A(n_7762),
.B(n_119),
.C(n_120),
.Y(n_8081)
);

NAND2xp5_ASAP7_75t_SL g8082 ( 
.A(n_7847),
.B(n_510),
.Y(n_8082)
);

AOI21xp33_ASAP7_75t_L g8083 ( 
.A1(n_7788),
.A2(n_120),
.B(n_121),
.Y(n_8083)
);

AOI21xp5_ASAP7_75t_L g8084 ( 
.A1(n_7824),
.A2(n_511),
.B(n_510),
.Y(n_8084)
);

OAI22xp5_ASAP7_75t_L g8085 ( 
.A1(n_7624),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_8085)
);

AOI21xp5_ASAP7_75t_L g8086 ( 
.A1(n_7763),
.A2(n_513),
.B(n_512),
.Y(n_8086)
);

OAI22xp5_ASAP7_75t_L g8087 ( 
.A1(n_7731),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_8087)
);

AOI21xp5_ASAP7_75t_L g8088 ( 
.A1(n_7758),
.A2(n_513),
.B(n_512),
.Y(n_8088)
);

OAI21xp33_ASAP7_75t_L g8089 ( 
.A1(n_7598),
.A2(n_122),
.B(n_123),
.Y(n_8089)
);

NAND3xp33_ASAP7_75t_L g8090 ( 
.A(n_7889),
.B(n_123),
.C(n_124),
.Y(n_8090)
);

OAI21xp5_ASAP7_75t_L g8091 ( 
.A1(n_7617),
.A2(n_124),
.B(n_125),
.Y(n_8091)
);

O2A1O1Ixp33_ASAP7_75t_L g8092 ( 
.A1(n_7789),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_8092)
);

NAND2xp5_ASAP7_75t_L g8093 ( 
.A(n_7653),
.B(n_7663),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_7443),
.Y(n_8094)
);

A2O1A1Ixp33_ASAP7_75t_L g8095 ( 
.A1(n_7667),
.A2(n_7704),
.B(n_7709),
.C(n_7688),
.Y(n_8095)
);

OAI21xp33_ASAP7_75t_L g8096 ( 
.A1(n_7735),
.A2(n_125),
.B(n_127),
.Y(n_8096)
);

NOR2xp33_ASAP7_75t_L g8097 ( 
.A(n_7608),
.B(n_514),
.Y(n_8097)
);

NAND2xp5_ASAP7_75t_SL g8098 ( 
.A(n_7844),
.B(n_514),
.Y(n_8098)
);

AOI21xp5_ASAP7_75t_L g8099 ( 
.A1(n_7626),
.A2(n_517),
.B(n_515),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_7455),
.Y(n_8100)
);

OAI21xp5_ASAP7_75t_L g8101 ( 
.A1(n_7746),
.A2(n_127),
.B(n_128),
.Y(n_8101)
);

INVx1_ASAP7_75t_L g8102 ( 
.A(n_7458),
.Y(n_8102)
);

NOR2xp33_ASAP7_75t_L g8103 ( 
.A(n_7656),
.B(n_515),
.Y(n_8103)
);

OAI21x1_ASAP7_75t_L g8104 ( 
.A1(n_7432),
.A2(n_127),
.B(n_128),
.Y(n_8104)
);

BUFx4f_ASAP7_75t_L g8105 ( 
.A(n_7519),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7460),
.Y(n_8106)
);

AOI21xp5_ASAP7_75t_L g8107 ( 
.A1(n_7791),
.A2(n_519),
.B(n_518),
.Y(n_8107)
);

AOI21xp5_ASAP7_75t_L g8108 ( 
.A1(n_7809),
.A2(n_520),
.B(n_518),
.Y(n_8108)
);

AOI21x1_ASAP7_75t_L g8109 ( 
.A1(n_7438),
.A2(n_129),
.B(n_131),
.Y(n_8109)
);

O2A1O1Ixp33_ASAP7_75t_L g8110 ( 
.A1(n_7792),
.A2(n_132),
.B(n_129),
.C(n_131),
.Y(n_8110)
);

BUFx6f_ASAP7_75t_L g8111 ( 
.A(n_7685),
.Y(n_8111)
);

NAND3xp33_ASAP7_75t_L g8112 ( 
.A(n_7895),
.B(n_129),
.C(n_132),
.Y(n_8112)
);

AOI21xp5_ASAP7_75t_L g8113 ( 
.A1(n_7752),
.A2(n_521),
.B(n_520),
.Y(n_8113)
);

A2O1A1Ixp33_ASAP7_75t_L g8114 ( 
.A1(n_7826),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_8114)
);

INVx2_ASAP7_75t_L g8115 ( 
.A(n_7880),
.Y(n_8115)
);

AOI21xp5_ASAP7_75t_L g8116 ( 
.A1(n_7578),
.A2(n_522),
.B(n_521),
.Y(n_8116)
);

HB1xp67_ASAP7_75t_L g8117 ( 
.A(n_7906),
.Y(n_8117)
);

OAI321xp33_ASAP7_75t_L g8118 ( 
.A1(n_7754),
.A2(n_135),
.A3(n_137),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_8118)
);

O2A1O1Ixp5_ASAP7_75t_L g8119 ( 
.A1(n_7642),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_8119)
);

AOI21xp5_ASAP7_75t_L g8120 ( 
.A1(n_7470),
.A2(n_523),
.B(n_522),
.Y(n_8120)
);

OAI21xp5_ASAP7_75t_L g8121 ( 
.A1(n_7596),
.A2(n_136),
.B(n_137),
.Y(n_8121)
);

AOI21xp5_ASAP7_75t_L g8122 ( 
.A1(n_7536),
.A2(n_524),
.B(n_523),
.Y(n_8122)
);

CKINVDCx8_ASAP7_75t_R g8123 ( 
.A(n_7877),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_L g8124 ( 
.A(n_7550),
.B(n_137),
.Y(n_8124)
);

AOI21xp5_ASAP7_75t_L g8125 ( 
.A1(n_7859),
.A2(n_525),
.B(n_524),
.Y(n_8125)
);

AOI21xp5_ASAP7_75t_L g8126 ( 
.A1(n_7865),
.A2(n_526),
.B(n_525),
.Y(n_8126)
);

NAND3xp33_ASAP7_75t_L g8127 ( 
.A(n_7903),
.B(n_138),
.C(n_139),
.Y(n_8127)
);

AOI21xp5_ASAP7_75t_L g8128 ( 
.A1(n_7702),
.A2(n_528),
.B(n_526),
.Y(n_8128)
);

NAND2xp5_ASAP7_75t_L g8129 ( 
.A(n_7550),
.B(n_138),
.Y(n_8129)
);

OAI21xp5_ASAP7_75t_L g8130 ( 
.A1(n_7569),
.A2(n_139),
.B(n_140),
.Y(n_8130)
);

NOR2xp33_ASAP7_75t_R g8131 ( 
.A(n_7434),
.B(n_529),
.Y(n_8131)
);

INVx1_ASAP7_75t_L g8132 ( 
.A(n_7896),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_7907),
.Y(n_8133)
);

NAND2xp5_ASAP7_75t_L g8134 ( 
.A(n_7550),
.B(n_7706),
.Y(n_8134)
);

AOI22xp5_ASAP7_75t_L g8135 ( 
.A1(n_7518),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_8135)
);

NAND2xp5_ASAP7_75t_L g8136 ( 
.A(n_7430),
.B(n_140),
.Y(n_8136)
);

INVx3_ASAP7_75t_L g8137 ( 
.A(n_7674),
.Y(n_8137)
);

O2A1O1Ixp33_ASAP7_75t_L g8138 ( 
.A1(n_7886),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_8138)
);

BUFx6f_ASAP7_75t_L g8139 ( 
.A(n_7454),
.Y(n_8139)
);

NAND2xp5_ASAP7_75t_L g8140 ( 
.A(n_7884),
.B(n_7913),
.Y(n_8140)
);

INVx3_ASAP7_75t_L g8141 ( 
.A(n_7567),
.Y(n_8141)
);

INVx3_ASAP7_75t_L g8142 ( 
.A(n_7812),
.Y(n_8142)
);

OAI21xp33_ASAP7_75t_L g8143 ( 
.A1(n_7582),
.A2(n_141),
.B(n_142),
.Y(n_8143)
);

AOI21xp5_ASAP7_75t_L g8144 ( 
.A1(n_7475),
.A2(n_530),
.B(n_529),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_7908),
.Y(n_8145)
);

INVx2_ASAP7_75t_L g8146 ( 
.A(n_7909),
.Y(n_8146)
);

AOI21xp5_ASAP7_75t_L g8147 ( 
.A1(n_7871),
.A2(n_531),
.B(n_530),
.Y(n_8147)
);

AND2x2_ASAP7_75t_L g8148 ( 
.A(n_7665),
.B(n_143),
.Y(n_8148)
);

NAND2xp5_ASAP7_75t_L g8149 ( 
.A(n_7509),
.B(n_144),
.Y(n_8149)
);

INVx3_ASAP7_75t_L g8150 ( 
.A(n_7490),
.Y(n_8150)
);

NAND2xp5_ASAP7_75t_L g8151 ( 
.A(n_7518),
.B(n_144),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_7910),
.Y(n_8152)
);

AOI21xp5_ASAP7_75t_L g8153 ( 
.A1(n_7829),
.A2(n_532),
.B(n_531),
.Y(n_8153)
);

OAI22xp5_ASAP7_75t_L g8154 ( 
.A1(n_7473),
.A2(n_7453),
.B1(n_7439),
.B2(n_7522),
.Y(n_8154)
);

AOI21xp5_ASAP7_75t_L g8155 ( 
.A1(n_7575),
.A2(n_533),
.B(n_532),
.Y(n_8155)
);

AO22x1_ASAP7_75t_L g8156 ( 
.A1(n_7914),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7911),
.Y(n_8157)
);

NAND2xp5_ASAP7_75t_L g8158 ( 
.A(n_7518),
.B(n_145),
.Y(n_8158)
);

OR2x2_ASAP7_75t_L g8159 ( 
.A(n_7551),
.B(n_533),
.Y(n_8159)
);

NOR2xp33_ASAP7_75t_L g8160 ( 
.A(n_7854),
.B(n_534),
.Y(n_8160)
);

AOI21x1_ASAP7_75t_L g8161 ( 
.A1(n_7553),
.A2(n_146),
.B(n_147),
.Y(n_8161)
);

NAND2xp5_ASAP7_75t_L g8162 ( 
.A(n_7534),
.B(n_146),
.Y(n_8162)
);

NAND2xp5_ASAP7_75t_L g8163 ( 
.A(n_7534),
.B(n_147),
.Y(n_8163)
);

OAI21xp33_ASAP7_75t_L g8164 ( 
.A1(n_7593),
.A2(n_148),
.B(n_149),
.Y(n_8164)
);

NAND2xp5_ASAP7_75t_L g8165 ( 
.A(n_7534),
.B(n_148),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7589),
.B(n_149),
.Y(n_8166)
);

AOI21xp5_ASAP7_75t_L g8167 ( 
.A1(n_7594),
.A2(n_535),
.B(n_534),
.Y(n_8167)
);

OAI22xp5_ASAP7_75t_L g8168 ( 
.A1(n_7469),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_8168)
);

AO21x1_ASAP7_75t_L g8169 ( 
.A1(n_7876),
.A2(n_7919),
.B(n_7868),
.Y(n_8169)
);

NOR2x1_ASAP7_75t_L g8170 ( 
.A(n_7489),
.B(n_7767),
.Y(n_8170)
);

NAND2xp5_ASAP7_75t_L g8171 ( 
.A(n_7659),
.B(n_150),
.Y(n_8171)
);

AOI21xp5_ASAP7_75t_L g8172 ( 
.A1(n_7923),
.A2(n_7479),
.B(n_7477),
.Y(n_8172)
);

O2A1O1Ixp33_ASAP7_75t_L g8173 ( 
.A1(n_7912),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_8173)
);

AOI21xp5_ASAP7_75t_L g8174 ( 
.A1(n_7480),
.A2(n_536),
.B(n_535),
.Y(n_8174)
);

OAI21xp5_ASAP7_75t_L g8175 ( 
.A1(n_7530),
.A2(n_151),
.B(n_152),
.Y(n_8175)
);

NOR2xp33_ASAP7_75t_L g8176 ( 
.A(n_7856),
.B(n_536),
.Y(n_8176)
);

AND2x2_ASAP7_75t_L g8177 ( 
.A(n_7733),
.B(n_153),
.Y(n_8177)
);

NAND2xp5_ASAP7_75t_L g8178 ( 
.A(n_7797),
.B(n_154),
.Y(n_8178)
);

INVx1_ASAP7_75t_SL g8179 ( 
.A(n_7785),
.Y(n_8179)
);

NAND2xp5_ASAP7_75t_L g8180 ( 
.A(n_7801),
.B(n_154),
.Y(n_8180)
);

AO21x1_ASAP7_75t_L g8181 ( 
.A1(n_7860),
.A2(n_538),
.B(n_537),
.Y(n_8181)
);

AND2x2_ASAP7_75t_L g8182 ( 
.A(n_7756),
.B(n_154),
.Y(n_8182)
);

NAND2xp5_ASAP7_75t_L g8183 ( 
.A(n_7478),
.B(n_155),
.Y(n_8183)
);

AOI22x1_ASAP7_75t_L g8184 ( 
.A1(n_7623),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_8184)
);

INVx3_ASAP7_75t_L g8185 ( 
.A(n_7781),
.Y(n_8185)
);

AND2x2_ASAP7_75t_L g8186 ( 
.A(n_7849),
.B(n_155),
.Y(n_8186)
);

OAI21xp33_ASAP7_75t_L g8187 ( 
.A1(n_7467),
.A2(n_7474),
.B(n_7456),
.Y(n_8187)
);

INVx1_ASAP7_75t_L g8188 ( 
.A(n_7555),
.Y(n_8188)
);

INVx4_ASAP7_75t_L g8189 ( 
.A(n_7768),
.Y(n_8189)
);

INVx1_ASAP7_75t_L g8190 ( 
.A(n_7482),
.Y(n_8190)
);

AOI21xp5_ASAP7_75t_L g8191 ( 
.A1(n_7483),
.A2(n_538),
.B(n_537),
.Y(n_8191)
);

AOI21xp5_ASAP7_75t_L g8192 ( 
.A1(n_7484),
.A2(n_540),
.B(n_539),
.Y(n_8192)
);

AND2x2_ASAP7_75t_L g8193 ( 
.A(n_7743),
.B(n_156),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7486),
.Y(n_8194)
);

INVx1_ASAP7_75t_L g8195 ( 
.A(n_7487),
.Y(n_8195)
);

INVx4_ASAP7_75t_L g8196 ( 
.A(n_7549),
.Y(n_8196)
);

NAND2xp5_ASAP7_75t_L g8197 ( 
.A(n_7446),
.B(n_156),
.Y(n_8197)
);

AOI21x1_ASAP7_75t_L g8198 ( 
.A1(n_7872),
.A2(n_157),
.B(n_158),
.Y(n_8198)
);

AOI21xp5_ASAP7_75t_L g8199 ( 
.A1(n_7491),
.A2(n_542),
.B(n_541),
.Y(n_8199)
);

NOR2xp33_ASAP7_75t_L g8200 ( 
.A(n_7861),
.B(n_541),
.Y(n_8200)
);

AOI21xp5_ASAP7_75t_L g8201 ( 
.A1(n_7493),
.A2(n_544),
.B(n_543),
.Y(n_8201)
);

AOI21xp5_ASAP7_75t_L g8202 ( 
.A1(n_7676),
.A2(n_544),
.B(n_543),
.Y(n_8202)
);

NAND2xp5_ASAP7_75t_L g8203 ( 
.A(n_7448),
.B(n_7494),
.Y(n_8203)
);

O2A1O1Ixp33_ASAP7_75t_L g8204 ( 
.A1(n_7644),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_8204)
);

AOI21xp5_ASAP7_75t_L g8205 ( 
.A1(n_7532),
.A2(n_546),
.B(n_545),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_7542),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_7544),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_7556),
.Y(n_8208)
);

NAND2xp5_ASAP7_75t_L g8209 ( 
.A(n_7496),
.B(n_158),
.Y(n_8209)
);

INVxp67_ASAP7_75t_L g8210 ( 
.A(n_7671),
.Y(n_8210)
);

OAI21xp5_ASAP7_75t_L g8211 ( 
.A1(n_7873),
.A2(n_159),
.B(n_160),
.Y(n_8211)
);

AOI21xp5_ASAP7_75t_L g8212 ( 
.A1(n_7535),
.A2(n_549),
.B(n_548),
.Y(n_8212)
);

OAI21xp5_ASAP7_75t_L g8213 ( 
.A1(n_7651),
.A2(n_160),
.B(n_161),
.Y(n_8213)
);

NOR2xp33_ASAP7_75t_L g8214 ( 
.A(n_7863),
.B(n_549),
.Y(n_8214)
);

OAI21xp5_ASAP7_75t_L g8215 ( 
.A1(n_7670),
.A2(n_160),
.B(n_161),
.Y(n_8215)
);

BUFx2_ASAP7_75t_L g8216 ( 
.A(n_7887),
.Y(n_8216)
);

INVx2_ASAP7_75t_L g8217 ( 
.A(n_7558),
.Y(n_8217)
);

INVxp67_ASAP7_75t_L g8218 ( 
.A(n_7778),
.Y(n_8218)
);

INVx2_ASAP7_75t_L g8219 ( 
.A(n_7498),
.Y(n_8219)
);

AO32x1_ASAP7_75t_L g8220 ( 
.A1(n_7581),
.A2(n_163),
.A3(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_8220)
);

OAI21xp5_ASAP7_75t_L g8221 ( 
.A1(n_7793),
.A2(n_162),
.B(n_163),
.Y(n_8221)
);

NOR2xp33_ASAP7_75t_L g8222 ( 
.A(n_7584),
.B(n_551),
.Y(n_8222)
);

OAI21xp33_ASAP7_75t_L g8223 ( 
.A1(n_7729),
.A2(n_162),
.B(n_163),
.Y(n_8223)
);

AOI21xp5_ASAP7_75t_L g8224 ( 
.A1(n_7852),
.A2(n_7736),
.B(n_7633),
.Y(n_8224)
);

NOR2xp33_ASAP7_75t_L g8225 ( 
.A(n_7546),
.B(n_551),
.Y(n_8225)
);

AOI21xp5_ASAP7_75t_L g8226 ( 
.A1(n_7669),
.A2(n_553),
.B(n_552),
.Y(n_8226)
);

AOI22xp5_ASAP7_75t_L g8227 ( 
.A1(n_7858),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_8227)
);

AOI21xp5_ASAP7_75t_L g8228 ( 
.A1(n_7630),
.A2(n_554),
.B(n_552),
.Y(n_8228)
);

AOI22xp5_ASAP7_75t_L g8229 ( 
.A1(n_7858),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_8229)
);

BUFx3_ASAP7_75t_L g8230 ( 
.A(n_7682),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_7502),
.B(n_165),
.Y(n_8231)
);

AOI21xp5_ASAP7_75t_L g8232 ( 
.A1(n_7537),
.A2(n_555),
.B(n_554),
.Y(n_8232)
);

NAND2xp5_ASAP7_75t_L g8233 ( 
.A(n_7506),
.B(n_167),
.Y(n_8233)
);

OAI22xp5_ASAP7_75t_L g8234 ( 
.A1(n_7834),
.A2(n_7599),
.B1(n_7571),
.B2(n_7501),
.Y(n_8234)
);

OR2x2_ASAP7_75t_L g8235 ( 
.A(n_7874),
.B(n_556),
.Y(n_8235)
);

NAND2xp5_ASAP7_75t_L g8236 ( 
.A(n_7510),
.B(n_7511),
.Y(n_8236)
);

AOI21xp5_ASAP7_75t_L g8237 ( 
.A1(n_7538),
.A2(n_557),
.B(n_556),
.Y(n_8237)
);

AOI21xp5_ASAP7_75t_L g8238 ( 
.A1(n_7514),
.A2(n_558),
.B(n_557),
.Y(n_8238)
);

O2A1O1Ixp33_ASAP7_75t_L g8239 ( 
.A1(n_7869),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_8239)
);

AOI21xp5_ASAP7_75t_L g8240 ( 
.A1(n_7515),
.A2(n_559),
.B(n_558),
.Y(n_8240)
);

AOI21xp5_ASAP7_75t_L g8241 ( 
.A1(n_7517),
.A2(n_561),
.B(n_560),
.Y(n_8241)
);

NAND2xp5_ASAP7_75t_L g8242 ( 
.A(n_7521),
.B(n_167),
.Y(n_8242)
);

HB1xp67_ASAP7_75t_L g8243 ( 
.A(n_7779),
.Y(n_8243)
);

A2O1A1Ixp33_ASAP7_75t_L g8244 ( 
.A1(n_7921),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_8244)
);

INVx2_ASAP7_75t_L g8245 ( 
.A(n_7523),
.Y(n_8245)
);

AND2x2_ASAP7_75t_L g8246 ( 
.A(n_7749),
.B(n_168),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_7755),
.B(n_169),
.Y(n_8247)
);

AOI21xp5_ASAP7_75t_L g8248 ( 
.A1(n_7562),
.A2(n_7568),
.B(n_7565),
.Y(n_8248)
);

A2O1A1Ixp33_ASAP7_75t_L g8249 ( 
.A1(n_7765),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_8249)
);

AND2x2_ASAP7_75t_SL g8250 ( 
.A(n_7705),
.B(n_560),
.Y(n_8250)
);

AOI21xp5_ASAP7_75t_L g8251 ( 
.A1(n_7459),
.A2(n_563),
.B(n_562),
.Y(n_8251)
);

OAI21xp33_ASAP7_75t_L g8252 ( 
.A1(n_7512),
.A2(n_170),
.B(n_171),
.Y(n_8252)
);

NOR2xp33_ASAP7_75t_L g8253 ( 
.A(n_7620),
.B(n_562),
.Y(n_8253)
);

OAI22xp5_ASAP7_75t_L g8254 ( 
.A1(n_7552),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_8254)
);

AOI21xp5_ASAP7_75t_L g8255 ( 
.A1(n_7711),
.A2(n_565),
.B(n_564),
.Y(n_8255)
);

NAND2xp5_ASAP7_75t_L g8256 ( 
.A(n_7540),
.B(n_172),
.Y(n_8256)
);

NOR2xp33_ASAP7_75t_L g8257 ( 
.A(n_7848),
.B(n_564),
.Y(n_8257)
);

BUFx8_ASAP7_75t_L g8258 ( 
.A(n_7814),
.Y(n_8258)
);

AOI22xp5_ASAP7_75t_L g8259 ( 
.A1(n_7825),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_8259)
);

AOI21xp5_ASAP7_75t_L g8260 ( 
.A1(n_7766),
.A2(n_566),
.B(n_565),
.Y(n_8260)
);

INVx2_ASAP7_75t_L g8261 ( 
.A(n_7583),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_L g8262 ( 
.A(n_7481),
.B(n_174),
.Y(n_8262)
);

INVx1_ASAP7_75t_SL g8263 ( 
.A(n_7780),
.Y(n_8263)
);

O2A1O1Ixp33_ASAP7_75t_L g8264 ( 
.A1(n_7790),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_8264)
);

A2O1A1Ixp33_ASAP7_75t_L g8265 ( 
.A1(n_7855),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_8265)
);

AOI21xp5_ASAP7_75t_L g8266 ( 
.A1(n_7684),
.A2(n_567),
.B(n_566),
.Y(n_8266)
);

AND2x2_ASAP7_75t_L g8267 ( 
.A(n_7713),
.B(n_177),
.Y(n_8267)
);

A2O1A1Ixp33_ASAP7_75t_L g8268 ( 
.A1(n_7686),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_8268)
);

AOI21xp5_ASAP7_75t_L g8269 ( 
.A1(n_7563),
.A2(n_568),
.B(n_567),
.Y(n_8269)
);

INVxp67_ASAP7_75t_L g8270 ( 
.A(n_7658),
.Y(n_8270)
);

O2A1O1Ixp33_ASAP7_75t_L g8271 ( 
.A1(n_7745),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_7488),
.B(n_7817),
.Y(n_8272)
);

A2O1A1Ixp33_ASAP7_75t_L g8273 ( 
.A1(n_7660),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_8273)
);

NAND2xp5_ASAP7_75t_L g8274 ( 
.A(n_7560),
.B(n_181),
.Y(n_8274)
);

INVx1_ASAP7_75t_SL g8275 ( 
.A(n_7566),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_7621),
.Y(n_8276)
);

AOI21xp5_ASAP7_75t_L g8277 ( 
.A1(n_7627),
.A2(n_569),
.B(n_568),
.Y(n_8277)
);

INVx11_ASAP7_75t_L g8278 ( 
.A(n_7442),
.Y(n_8278)
);

AND2x2_ASAP7_75t_L g8279 ( 
.A(n_7853),
.B(n_7652),
.Y(n_8279)
);

NOR2xp33_ASAP7_75t_L g8280 ( 
.A(n_7828),
.B(n_7579),
.Y(n_8280)
);

INVx2_ASAP7_75t_L g8281 ( 
.A(n_7585),
.Y(n_8281)
);

INVx11_ASAP7_75t_L g8282 ( 
.A(n_7449),
.Y(n_8282)
);

AOI21xp5_ASAP7_75t_L g8283 ( 
.A1(n_7586),
.A2(n_571),
.B(n_569),
.Y(n_8283)
);

AOI21xp5_ASAP7_75t_L g8284 ( 
.A1(n_7591),
.A2(n_572),
.B(n_571),
.Y(n_8284)
);

AO21x1_ASAP7_75t_L g8285 ( 
.A1(n_7657),
.A2(n_573),
.B(n_572),
.Y(n_8285)
);

AOI21xp5_ASAP7_75t_L g8286 ( 
.A1(n_7592),
.A2(n_7604),
.B(n_7597),
.Y(n_8286)
);

A2O1A1Ixp33_ASAP7_75t_L g8287 ( 
.A1(n_7632),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_8287)
);

OAI22xp5_ASAP7_75t_L g8288 ( 
.A1(n_7611),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_8288)
);

BUFx6f_ASAP7_75t_L g8289 ( 
.A(n_7878),
.Y(n_8289)
);

NOR2x1_ASAP7_75t_L g8290 ( 
.A(n_7820),
.B(n_7574),
.Y(n_8290)
);

NOR2x1_ASAP7_75t_R g8291 ( 
.A(n_7742),
.B(n_573),
.Y(n_8291)
);

AOI21xp5_ASAP7_75t_L g8292 ( 
.A1(n_7606),
.A2(n_576),
.B(n_574),
.Y(n_8292)
);

INVx3_ASAP7_75t_L g8293 ( 
.A(n_7690),
.Y(n_8293)
);

AO21x1_ASAP7_75t_L g8294 ( 
.A1(n_7643),
.A2(n_577),
.B(n_574),
.Y(n_8294)
);

INVx3_ASAP7_75t_L g8295 ( 
.A(n_7719),
.Y(n_8295)
);

INVx3_ASAP7_75t_L g8296 ( 
.A(n_7503),
.Y(n_8296)
);

NAND2xp5_ASAP7_75t_L g8297 ( 
.A(n_7825),
.B(n_182),
.Y(n_8297)
);

NAND2xp5_ASAP7_75t_L g8298 ( 
.A(n_7825),
.B(n_183),
.Y(n_8298)
);

AOI21xp5_ASAP7_75t_L g8299 ( 
.A1(n_7607),
.A2(n_580),
.B(n_577),
.Y(n_8299)
);

AOI21xp5_ASAP7_75t_L g8300 ( 
.A1(n_7612),
.A2(n_581),
.B(n_580),
.Y(n_8300)
);

AND2x4_ASAP7_75t_L g8301 ( 
.A(n_7796),
.B(n_581),
.Y(n_8301)
);

OAI22xp5_ASAP7_75t_L g8302 ( 
.A1(n_7622),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_8302)
);

O2A1O1Ixp33_ASAP7_75t_L g8303 ( 
.A1(n_7783),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_L g8304 ( 
.A(n_7691),
.B(n_186),
.Y(n_8304)
);

AND2x2_ASAP7_75t_L g8305 ( 
.A(n_7680),
.B(n_187),
.Y(n_8305)
);

NOR2xp33_ASAP7_75t_L g8306 ( 
.A(n_7580),
.B(n_7500),
.Y(n_8306)
);

BUFx12f_ASAP7_75t_L g8307 ( 
.A(n_7925),
.Y(n_8307)
);

NAND2xp5_ASAP7_75t_SL g8308 ( 
.A(n_7870),
.B(n_582),
.Y(n_8308)
);

INVx2_ASAP7_75t_SL g8309 ( 
.A(n_7573),
.Y(n_8309)
);

NOR2xp33_ASAP7_75t_L g8310 ( 
.A(n_7696),
.B(n_582),
.Y(n_8310)
);

AND2x4_ASAP7_75t_L g8311 ( 
.A(n_7800),
.B(n_583),
.Y(n_8311)
);

OAI21xp5_ASAP7_75t_L g8312 ( 
.A1(n_7543),
.A2(n_187),
.B(n_188),
.Y(n_8312)
);

NAND3xp33_ASAP7_75t_L g8313 ( 
.A(n_7595),
.B(n_187),
.C(n_188),
.Y(n_8313)
);

NAND2xp5_ASAP7_75t_SL g8314 ( 
.A(n_7614),
.B(n_583),
.Y(n_8314)
);

NAND2xp5_ASAP7_75t_SL g8315 ( 
.A(n_7616),
.B(n_584),
.Y(n_8315)
);

INVx1_ASAP7_75t_L g8316 ( 
.A(n_7625),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7757),
.Y(n_8317)
);

AOI21xp5_ASAP7_75t_L g8318 ( 
.A1(n_7753),
.A2(n_585),
.B(n_584),
.Y(n_8318)
);

AOI21xp5_ASAP7_75t_L g8319 ( 
.A1(n_7891),
.A2(n_586),
.B(n_585),
.Y(n_8319)
);

NAND2xp5_ASAP7_75t_L g8320 ( 
.A(n_7609),
.B(n_189),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7662),
.Y(n_8321)
);

AOI21xp5_ASAP7_75t_L g8322 ( 
.A1(n_7901),
.A2(n_587),
.B(n_586),
.Y(n_8322)
);

OAI21xp5_ASAP7_75t_L g8323 ( 
.A1(n_7666),
.A2(n_189),
.B(n_190),
.Y(n_8323)
);

AOI22xp33_ASAP7_75t_L g8324 ( 
.A1(n_7914),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_7664),
.Y(n_8325)
);

A2O1A1Ixp33_ASAP7_75t_L g8326 ( 
.A1(n_7661),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_8326)
);

INVx2_ASAP7_75t_L g8327 ( 
.A(n_7672),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_L g8328 ( 
.A(n_7673),
.B(n_7675),
.Y(n_8328)
);

O2A1O1Ixp33_ASAP7_75t_L g8329 ( 
.A1(n_7867),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_8329)
);

NAND2xp5_ASAP7_75t_L g8330 ( 
.A(n_7914),
.B(n_192),
.Y(n_8330)
);

NAND2xp5_ASAP7_75t_L g8331 ( 
.A(n_7700),
.B(n_193),
.Y(n_8331)
);

NAND2xp5_ASAP7_75t_SL g8332 ( 
.A(n_7806),
.B(n_587),
.Y(n_8332)
);

AOI21xp5_ASAP7_75t_L g8333 ( 
.A1(n_7904),
.A2(n_589),
.B(n_588),
.Y(n_8333)
);

INVx2_ASAP7_75t_L g8334 ( 
.A(n_7726),
.Y(n_8334)
);

INVx2_ASAP7_75t_L g8335 ( 
.A(n_7805),
.Y(n_8335)
);

BUFx3_ASAP7_75t_L g8336 ( 
.A(n_7810),
.Y(n_8336)
);

NAND2xp5_ASAP7_75t_L g8337 ( 
.A(n_7547),
.B(n_194),
.Y(n_8337)
);

NOR2xp33_ASAP7_75t_L g8338 ( 
.A(n_7760),
.B(n_588),
.Y(n_8338)
);

NAND2xp5_ASAP7_75t_SL g8339 ( 
.A(n_7602),
.B(n_589),
.Y(n_8339)
);

NAND2xp5_ASAP7_75t_L g8340 ( 
.A(n_7548),
.B(n_194),
.Y(n_8340)
);

NAND2xp5_ASAP7_75t_L g8341 ( 
.A(n_7610),
.B(n_195),
.Y(n_8341)
);

AOI21xp33_ASAP7_75t_L g8342 ( 
.A1(n_7601),
.A2(n_7922),
.B(n_7918),
.Y(n_8342)
);

OAI22xp5_ASAP7_75t_L g8343 ( 
.A1(n_7808),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_8343)
);

AOI21x1_ASAP7_75t_L g8344 ( 
.A1(n_7720),
.A2(n_195),
.B(n_196),
.Y(n_8344)
);

OR2x6_ASAP7_75t_SL g8345 ( 
.A(n_7850),
.B(n_196),
.Y(n_8345)
);

NOR2xp67_ASAP7_75t_L g8346 ( 
.A(n_7841),
.B(n_197),
.Y(n_8346)
);

AOI22xp5_ASAP7_75t_L g8347 ( 
.A1(n_7610),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_8347)
);

OAI21xp5_ASAP7_75t_L g8348 ( 
.A1(n_7610),
.A2(n_198),
.B(n_199),
.Y(n_8348)
);

INVx1_ASAP7_75t_L g8349 ( 
.A(n_7738),
.Y(n_8349)
);

AOI22xp5_ASAP7_75t_L g8350 ( 
.A1(n_7866),
.A2(n_201),
.B1(n_198),
.B2(n_200),
.Y(n_8350)
);

NAND3xp33_ASAP7_75t_L g8351 ( 
.A(n_7740),
.B(n_200),
.C(n_201),
.Y(n_8351)
);

AOI21xp5_ASAP7_75t_L g8352 ( 
.A1(n_7795),
.A2(n_591),
.B(n_590),
.Y(n_8352)
);

AND2x2_ASAP7_75t_L g8353 ( 
.A(n_7845),
.B(n_201),
.Y(n_8353)
);

AND2x6_ASAP7_75t_L g8354 ( 
.A(n_7857),
.B(n_590),
.Y(n_8354)
);

OAI21x1_ASAP7_75t_L g8355 ( 
.A1(n_7588),
.A2(n_7648),
.B(n_7590),
.Y(n_8355)
);

AOI21xp5_ASAP7_75t_L g8356 ( 
.A1(n_7835),
.A2(n_592),
.B(n_591),
.Y(n_8356)
);

AO21x1_ASAP7_75t_L g8357 ( 
.A1(n_7786),
.A2(n_593),
.B(n_592),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_7723),
.Y(n_8358)
);

HB1xp67_ASAP7_75t_L g8359 ( 
.A(n_7885),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7631),
.Y(n_8360)
);

A2O1A1Ixp33_ASAP7_75t_L g8361 ( 
.A1(n_7890),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_8361)
);

AOI21xp5_ASAP7_75t_L g8362 ( 
.A1(n_7559),
.A2(n_594),
.B(n_593),
.Y(n_8362)
);

NAND2xp5_ASAP7_75t_L g8363 ( 
.A(n_7769),
.B(n_202),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7799),
.Y(n_8364)
);

AOI21xp5_ASAP7_75t_L g8365 ( 
.A1(n_7816),
.A2(n_596),
.B(n_594),
.Y(n_8365)
);

AOI21xp5_ASAP7_75t_L g8366 ( 
.A1(n_7774),
.A2(n_599),
.B(n_597),
.Y(n_8366)
);

INVx3_ASAP7_75t_L g8367 ( 
.A(n_7728),
.Y(n_8367)
);

CKINVDCx11_ASAP7_75t_R g8368 ( 
.A(n_7634),
.Y(n_8368)
);

O2A1O1Ixp33_ASAP7_75t_L g8369 ( 
.A1(n_7689),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_8369)
);

NAND2xp5_ASAP7_75t_L g8370 ( 
.A(n_7775),
.B(n_203),
.Y(n_8370)
);

AOI22x1_ASAP7_75t_L g8371 ( 
.A1(n_7703),
.A2(n_7708),
.B1(n_7716),
.B2(n_7526),
.Y(n_8371)
);

AOI21xp5_ASAP7_75t_L g8372 ( 
.A1(n_7898),
.A2(n_599),
.B(n_597),
.Y(n_8372)
);

AOI21xp5_ASAP7_75t_L g8373 ( 
.A1(n_7899),
.A2(n_601),
.B(n_600),
.Y(n_8373)
);

NAND2xp5_ASAP7_75t_SL g8374 ( 
.A(n_7916),
.B(n_600),
.Y(n_8374)
);

INVx2_ASAP7_75t_L g8375 ( 
.A(n_7603),
.Y(n_8375)
);

AND2x2_ASAP7_75t_L g8376 ( 
.A(n_7603),
.B(n_204),
.Y(n_8376)
);

INVx2_ASAP7_75t_SL g8377 ( 
.A(n_7777),
.Y(n_8377)
);

OAI22xp5_ASAP7_75t_L g8378 ( 
.A1(n_7603),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_8378)
);

OAI22xp5_ASAP7_75t_L g8379 ( 
.A1(n_7507),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7428),
.Y(n_8380)
);

NAND2xp5_ASAP7_75t_SL g8381 ( 
.A(n_7507),
.B(n_601),
.Y(n_8381)
);

BUFx12f_ASAP7_75t_L g8382 ( 
.A(n_7692),
.Y(n_8382)
);

OR2x2_ASAP7_75t_L g8383 ( 
.A(n_7613),
.B(n_602),
.Y(n_8383)
);

NAND2xp5_ASAP7_75t_SL g8384 ( 
.A(n_7507),
.B(n_602),
.Y(n_8384)
);

AOI21xp5_ASAP7_75t_L g8385 ( 
.A1(n_7461),
.A2(n_605),
.B(n_604),
.Y(n_8385)
);

INVx1_ASAP7_75t_SL g8386 ( 
.A(n_7882),
.Y(n_8386)
);

NOR2xp33_ASAP7_75t_L g8387 ( 
.A(n_7507),
.B(n_604),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7428),
.Y(n_8388)
);

AOI21xp5_ASAP7_75t_L g8389 ( 
.A1(n_7461),
.A2(n_608),
.B(n_606),
.Y(n_8389)
);

NAND3xp33_ASAP7_75t_L g8390 ( 
.A(n_7507),
.B(n_205),
.C(n_206),
.Y(n_8390)
);

OAI22xp5_ASAP7_75t_L g8391 ( 
.A1(n_7507),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_8391)
);

INVx2_ASAP7_75t_L g8392 ( 
.A(n_7428),
.Y(n_8392)
);

AND2x4_ASAP7_75t_L g8393 ( 
.A(n_7450),
.B(n_606),
.Y(n_8393)
);

NAND2xp5_ASAP7_75t_L g8394 ( 
.A(n_7507),
.B(n_208),
.Y(n_8394)
);

NAND2xp5_ASAP7_75t_L g8395 ( 
.A(n_7507),
.B(n_208),
.Y(n_8395)
);

AO21x1_ASAP7_75t_L g8396 ( 
.A1(n_7461),
.A2(n_609),
.B(n_608),
.Y(n_8396)
);

AOI21xp5_ASAP7_75t_L g8397 ( 
.A1(n_7461),
.A2(n_611),
.B(n_610),
.Y(n_8397)
);

NOR2xp33_ASAP7_75t_L g8398 ( 
.A(n_7507),
.B(n_610),
.Y(n_8398)
);

AND2x2_ASAP7_75t_L g8399 ( 
.A(n_7830),
.B(n_209),
.Y(n_8399)
);

NAND2xp5_ASAP7_75t_L g8400 ( 
.A(n_7507),
.B(n_209),
.Y(n_8400)
);

NAND2xp5_ASAP7_75t_L g8401 ( 
.A(n_7507),
.B(n_210),
.Y(n_8401)
);

AOI21xp5_ASAP7_75t_L g8402 ( 
.A1(n_7461),
.A2(n_612),
.B(n_611),
.Y(n_8402)
);

NOR2xp33_ASAP7_75t_L g8403 ( 
.A(n_7507),
.B(n_612),
.Y(n_8403)
);

AOI21xp5_ASAP7_75t_L g8404 ( 
.A1(n_7461),
.A2(n_614),
.B(n_613),
.Y(n_8404)
);

INVx2_ASAP7_75t_L g8405 ( 
.A(n_7428),
.Y(n_8405)
);

NAND2xp5_ASAP7_75t_L g8406 ( 
.A(n_7507),
.B(n_210),
.Y(n_8406)
);

O2A1O1Ixp5_ASAP7_75t_L g8407 ( 
.A1(n_7893),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_8407)
);

AOI21xp5_ASAP7_75t_L g8408 ( 
.A1(n_7461),
.A2(n_615),
.B(n_614),
.Y(n_8408)
);

INVx3_ASAP7_75t_L g8409 ( 
.A(n_7450),
.Y(n_8409)
);

NOR2xp33_ASAP7_75t_L g8410 ( 
.A(n_7507),
.B(n_615),
.Y(n_8410)
);

NOR2xp67_ASAP7_75t_L g8411 ( 
.A(n_7862),
.B(n_211),
.Y(n_8411)
);

NAND2xp5_ASAP7_75t_L g8412 ( 
.A(n_7507),
.B(n_211),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_7428),
.Y(n_8413)
);

AND2x4_ASAP7_75t_L g8414 ( 
.A(n_7450),
.B(n_616),
.Y(n_8414)
);

AO21x1_ASAP7_75t_L g8415 ( 
.A1(n_7461),
.A2(n_618),
.B(n_617),
.Y(n_8415)
);

AOI21xp5_ASAP7_75t_L g8416 ( 
.A1(n_7461),
.A2(n_618),
.B(n_617),
.Y(n_8416)
);

NAND2xp5_ASAP7_75t_L g8417 ( 
.A(n_7507),
.B(n_212),
.Y(n_8417)
);

AOI21xp5_ASAP7_75t_L g8418 ( 
.A1(n_7461),
.A2(n_620),
.B(n_619),
.Y(n_8418)
);

INVx2_ASAP7_75t_L g8419 ( 
.A(n_7428),
.Y(n_8419)
);

AOI21xp5_ASAP7_75t_L g8420 ( 
.A1(n_7461),
.A2(n_620),
.B(n_619),
.Y(n_8420)
);

AND2x4_ASAP7_75t_L g8421 ( 
.A(n_7450),
.B(n_621),
.Y(n_8421)
);

NAND2xp5_ASAP7_75t_SL g8422 ( 
.A(n_7507),
.B(n_622),
.Y(n_8422)
);

INVx1_ASAP7_75t_L g8423 ( 
.A(n_7428),
.Y(n_8423)
);

INVx2_ASAP7_75t_L g8424 ( 
.A(n_7428),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_7507),
.B(n_212),
.Y(n_8425)
);

AOI21xp5_ASAP7_75t_L g8426 ( 
.A1(n_7461),
.A2(n_623),
.B(n_622),
.Y(n_8426)
);

AOI22xp5_ASAP7_75t_L g8427 ( 
.A1(n_7507),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_8427)
);

INVx1_ASAP7_75t_L g8428 ( 
.A(n_7428),
.Y(n_8428)
);

O2A1O1Ixp33_ASAP7_75t_L g8429 ( 
.A1(n_7557),
.A2(n_216),
.B(n_213),
.C(n_214),
.Y(n_8429)
);

NAND2xp5_ASAP7_75t_L g8430 ( 
.A(n_7507),
.B(n_213),
.Y(n_8430)
);

BUFx6f_ASAP7_75t_L g8431 ( 
.A(n_7692),
.Y(n_8431)
);

AOI21xp5_ASAP7_75t_L g8432 ( 
.A1(n_7461),
.A2(n_626),
.B(n_623),
.Y(n_8432)
);

A2O1A1Ixp33_ASAP7_75t_L g8433 ( 
.A1(n_7507),
.A2(n_217),
.B(n_214),
.C(n_216),
.Y(n_8433)
);

NAND2xp5_ASAP7_75t_L g8434 ( 
.A(n_7507),
.B(n_216),
.Y(n_8434)
);

NAND2xp5_ASAP7_75t_L g8435 ( 
.A(n_7507),
.B(n_217),
.Y(n_8435)
);

AOI21xp5_ASAP7_75t_L g8436 ( 
.A1(n_7461),
.A2(n_627),
.B(n_626),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_SL g8437 ( 
.A(n_7507),
.B(n_627),
.Y(n_8437)
);

INVx2_ASAP7_75t_L g8438 ( 
.A(n_7428),
.Y(n_8438)
);

AOI21xp5_ASAP7_75t_L g8439 ( 
.A1(n_7461),
.A2(n_629),
.B(n_628),
.Y(n_8439)
);

OAI22xp5_ASAP7_75t_L g8440 ( 
.A1(n_7507),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_7507),
.B(n_218),
.Y(n_8441)
);

NAND2xp5_ASAP7_75t_L g8442 ( 
.A(n_7507),
.B(n_218),
.Y(n_8442)
);

INVxp67_ASAP7_75t_L g8443 ( 
.A(n_7906),
.Y(n_8443)
);

OAI22xp5_ASAP7_75t_L g8444 ( 
.A1(n_7507),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_8444)
);

OAI22xp5_ASAP7_75t_L g8445 ( 
.A1(n_7507),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_8445)
);

NAND2xp5_ASAP7_75t_SL g8446 ( 
.A(n_7507),
.B(n_628),
.Y(n_8446)
);

AND2x2_ASAP7_75t_L g8447 ( 
.A(n_7830),
.B(n_220),
.Y(n_8447)
);

A2O1A1Ixp33_ASAP7_75t_L g8448 ( 
.A1(n_7507),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_8448)
);

INVx4_ASAP7_75t_L g8449 ( 
.A(n_7471),
.Y(n_8449)
);

INVx2_ASAP7_75t_L g8450 ( 
.A(n_7428),
.Y(n_8450)
);

AND2x4_ASAP7_75t_L g8451 ( 
.A(n_7450),
.B(n_630),
.Y(n_8451)
);

INVx2_ASAP7_75t_SL g8452 ( 
.A(n_7587),
.Y(n_8452)
);

NAND2xp5_ASAP7_75t_L g8453 ( 
.A(n_7507),
.B(n_223),
.Y(n_8453)
);

NOR3xp33_ASAP7_75t_L g8454 ( 
.A(n_7557),
.B(n_223),
.C(n_224),
.Y(n_8454)
);

NAND2xp5_ASAP7_75t_L g8455 ( 
.A(n_7507),
.B(n_224),
.Y(n_8455)
);

O2A1O1Ixp33_ASAP7_75t_L g8456 ( 
.A1(n_7557),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_8456)
);

AND2x2_ASAP7_75t_L g8457 ( 
.A(n_7830),
.B(n_225),
.Y(n_8457)
);

NAND2xp5_ASAP7_75t_SL g8458 ( 
.A(n_7507),
.B(n_630),
.Y(n_8458)
);

NAND2xp5_ASAP7_75t_L g8459 ( 
.A(n_7507),
.B(n_226),
.Y(n_8459)
);

AOI21xp5_ASAP7_75t_L g8460 ( 
.A1(n_7461),
.A2(n_632),
.B(n_631),
.Y(n_8460)
);

OAI21xp33_ASAP7_75t_L g8461 ( 
.A1(n_7507),
.A2(n_227),
.B(n_228),
.Y(n_8461)
);

NOR2xp33_ASAP7_75t_L g8462 ( 
.A(n_7507),
.B(n_632),
.Y(n_8462)
);

HB1xp67_ASAP7_75t_L g8463 ( 
.A(n_7906),
.Y(n_8463)
);

BUFx4f_ASAP7_75t_L g8464 ( 
.A(n_7462),
.Y(n_8464)
);

AO22x1_ASAP7_75t_L g8465 ( 
.A1(n_7893),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_8465)
);

AOI21x1_ASAP7_75t_L g8466 ( 
.A1(n_7818),
.A2(n_228),
.B(n_229),
.Y(n_8466)
);

BUFx4f_ASAP7_75t_L g8467 ( 
.A(n_7462),
.Y(n_8467)
);

OAI321xp33_ASAP7_75t_L g8468 ( 
.A1(n_7507),
.A2(n_232),
.A3(n_234),
.B1(n_230),
.B2(n_231),
.C(n_233),
.Y(n_8468)
);

AND2x4_ASAP7_75t_L g8469 ( 
.A(n_7450),
.B(n_633),
.Y(n_8469)
);

NAND2xp5_ASAP7_75t_L g8470 ( 
.A(n_7926),
.B(n_634),
.Y(n_8470)
);

NOR2xp33_ASAP7_75t_L g8471 ( 
.A(n_7990),
.B(n_634),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_7930),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_7940),
.B(n_635),
.Y(n_8473)
);

OAI22xp5_ASAP7_75t_L g8474 ( 
.A1(n_8387),
.A2(n_8403),
.B1(n_8410),
.B2(n_8398),
.Y(n_8474)
);

AOI21xp5_ASAP7_75t_L g8475 ( 
.A1(n_7935),
.A2(n_636),
.B(n_635),
.Y(n_8475)
);

OAI221xp5_ASAP7_75t_L g8476 ( 
.A1(n_8462),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.C(n_234),
.Y(n_8476)
);

NAND3xp33_ASAP7_75t_SL g8477 ( 
.A(n_8454),
.B(n_231),
.C(n_232),
.Y(n_8477)
);

OAI22xp5_ASAP7_75t_L g8478 ( 
.A1(n_7932),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_8478)
);

BUFx6f_ASAP7_75t_L g8479 ( 
.A(n_7928),
.Y(n_8479)
);

HB1xp67_ASAP7_75t_L g8480 ( 
.A(n_8117),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_7991),
.Y(n_8481)
);

INVx2_ASAP7_75t_L g8482 ( 
.A(n_7956),
.Y(n_8482)
);

AND2x2_ASAP7_75t_L g8483 ( 
.A(n_8186),
.B(n_7927),
.Y(n_8483)
);

AOI21xp5_ASAP7_75t_L g8484 ( 
.A1(n_8006),
.A2(n_637),
.B(n_636),
.Y(n_8484)
);

NAND2xp5_ASAP7_75t_L g8485 ( 
.A(n_7945),
.B(n_7950),
.Y(n_8485)
);

AOI21xp5_ASAP7_75t_L g8486 ( 
.A1(n_7954),
.A2(n_639),
.B(n_638),
.Y(n_8486)
);

INVx2_ASAP7_75t_L g8487 ( 
.A(n_7968),
.Y(n_8487)
);

BUFx6f_ASAP7_75t_L g8488 ( 
.A(n_7928),
.Y(n_8488)
);

O2A1O1Ixp33_ASAP7_75t_L g8489 ( 
.A1(n_7931),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_8002),
.Y(n_8490)
);

NOR2xp67_ASAP7_75t_L g8491 ( 
.A(n_8449),
.B(n_237),
.Y(n_8491)
);

AOI21xp5_ASAP7_75t_L g8492 ( 
.A1(n_8013),
.A2(n_639),
.B(n_638),
.Y(n_8492)
);

CKINVDCx5p33_ASAP7_75t_R g8493 ( 
.A(n_7934),
.Y(n_8493)
);

INVx1_ASAP7_75t_L g8494 ( 
.A(n_8017),
.Y(n_8494)
);

OR2x6_ASAP7_75t_SL g8495 ( 
.A(n_8234),
.B(n_237),
.Y(n_8495)
);

NAND2xp5_ASAP7_75t_SL g8496 ( 
.A(n_8154),
.B(n_640),
.Y(n_8496)
);

AND2x4_ASAP7_75t_L g8497 ( 
.A(n_7948),
.B(n_641),
.Y(n_8497)
);

A2O1A1Ixp33_ASAP7_75t_L g8498 ( 
.A1(n_7984),
.A2(n_642),
.B(n_643),
.C(n_641),
.Y(n_8498)
);

INVx1_ASAP7_75t_L g8499 ( 
.A(n_8025),
.Y(n_8499)
);

NOR2x1_ASAP7_75t_L g8500 ( 
.A(n_8390),
.B(n_642),
.Y(n_8500)
);

INVx2_ASAP7_75t_L g8501 ( 
.A(n_7983),
.Y(n_8501)
);

OAI22xp5_ASAP7_75t_L g8502 ( 
.A1(n_8250),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_8502)
);

AOI21xp5_ASAP7_75t_L g8503 ( 
.A1(n_7933),
.A2(n_645),
.B(n_643),
.Y(n_8503)
);

OAI22xp5_ASAP7_75t_L g8504 ( 
.A1(n_8394),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_8504)
);

INVx1_ASAP7_75t_L g8505 ( 
.A(n_8030),
.Y(n_8505)
);

AND2x2_ASAP7_75t_L g8506 ( 
.A(n_8279),
.B(n_645),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_8072),
.Y(n_8507)
);

NAND3xp33_ASAP7_75t_SL g8508 ( 
.A(n_8042),
.B(n_239),
.C(n_240),
.Y(n_8508)
);

OAI21xp5_ASAP7_75t_L g8509 ( 
.A1(n_8095),
.A2(n_241),
.B(n_242),
.Y(n_8509)
);

INVx2_ASAP7_75t_L g8510 ( 
.A(n_7986),
.Y(n_8510)
);

OAI21xp5_ASAP7_75t_L g8511 ( 
.A1(n_8313),
.A2(n_241),
.B(n_242),
.Y(n_8511)
);

NAND2xp5_ASAP7_75t_L g8512 ( 
.A(n_8093),
.B(n_646),
.Y(n_8512)
);

INVx3_ASAP7_75t_L g8513 ( 
.A(n_8123),
.Y(n_8513)
);

AOI21xp5_ASAP7_75t_L g8514 ( 
.A1(n_8385),
.A2(n_648),
.B(n_647),
.Y(n_8514)
);

NAND2xp5_ASAP7_75t_SL g8515 ( 
.A(n_8134),
.B(n_647),
.Y(n_8515)
);

INVx4_ASAP7_75t_L g8516 ( 
.A(n_7928),
.Y(n_8516)
);

INVx1_ASAP7_75t_SL g8517 ( 
.A(n_7967),
.Y(n_8517)
);

NOR3xp33_ASAP7_75t_L g8518 ( 
.A(n_8121),
.B(n_242),
.C(n_243),
.Y(n_8518)
);

NAND2xp5_ASAP7_75t_L g8519 ( 
.A(n_8053),
.B(n_648),
.Y(n_8519)
);

INVx1_ASAP7_75t_L g8520 ( 
.A(n_8094),
.Y(n_8520)
);

AND2x4_ASAP7_75t_L g8521 ( 
.A(n_7948),
.B(n_649),
.Y(n_8521)
);

BUFx8_ASAP7_75t_L g8522 ( 
.A(n_8289),
.Y(n_8522)
);

INVx2_ASAP7_75t_L g8523 ( 
.A(n_8392),
.Y(n_8523)
);

INVx1_ASAP7_75t_L g8524 ( 
.A(n_8100),
.Y(n_8524)
);

O2A1O1Ixp33_ASAP7_75t_L g8525 ( 
.A1(n_7981),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_8102),
.Y(n_8526)
);

AND2x2_ASAP7_75t_L g8527 ( 
.A(n_8148),
.B(n_649),
.Y(n_8527)
);

NAND2xp5_ASAP7_75t_SL g8528 ( 
.A(n_8070),
.B(n_650),
.Y(n_8528)
);

NAND2xp5_ASAP7_75t_L g8529 ( 
.A(n_8463),
.B(n_650),
.Y(n_8529)
);

NAND2xp5_ASAP7_75t_SL g8530 ( 
.A(n_7964),
.B(n_652),
.Y(n_8530)
);

AND2x2_ASAP7_75t_SL g8531 ( 
.A(n_8005),
.B(n_653),
.Y(n_8531)
);

AND2x4_ASAP7_75t_L g8532 ( 
.A(n_7995),
.B(n_653),
.Y(n_8532)
);

OAI22xp5_ASAP7_75t_L g8533 ( 
.A1(n_8395),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_8533)
);

HB1xp67_ASAP7_75t_L g8534 ( 
.A(n_8243),
.Y(n_8534)
);

AND2x4_ASAP7_75t_L g8535 ( 
.A(n_8290),
.B(n_654),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_8106),
.Y(n_8536)
);

NAND2xp5_ASAP7_75t_L g8537 ( 
.A(n_8065),
.B(n_654),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_8132),
.Y(n_8538)
);

O2A1O1Ixp33_ASAP7_75t_L g8539 ( 
.A1(n_8429),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_8539)
);

NOR2xp33_ASAP7_75t_SL g8540 ( 
.A(n_8382),
.B(n_246),
.Y(n_8540)
);

INVx1_ASAP7_75t_L g8541 ( 
.A(n_8133),
.Y(n_8541)
);

INVx2_ASAP7_75t_L g8542 ( 
.A(n_8405),
.Y(n_8542)
);

A2O1A1Ixp33_ASAP7_75t_L g8543 ( 
.A1(n_8079),
.A2(n_656),
.B(n_657),
.C(n_655),
.Y(n_8543)
);

A2O1A1Ixp33_ASAP7_75t_L g8544 ( 
.A1(n_8110),
.A2(n_656),
.B(n_657),
.C(n_655),
.Y(n_8544)
);

AND2x2_ASAP7_75t_L g8545 ( 
.A(n_8177),
.B(n_658),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_L g8546 ( 
.A(n_8443),
.B(n_8400),
.Y(n_8546)
);

AOI21xp5_ASAP7_75t_L g8547 ( 
.A1(n_8389),
.A2(n_659),
.B(n_658),
.Y(n_8547)
);

AOI21xp33_ASAP7_75t_L g8548 ( 
.A1(n_8169),
.A2(n_246),
.B(n_247),
.Y(n_8548)
);

AOI21xp5_ASAP7_75t_L g8549 ( 
.A1(n_8397),
.A2(n_8404),
.B(n_8402),
.Y(n_8549)
);

NAND2xp5_ASAP7_75t_L g8550 ( 
.A(n_8401),
.B(n_659),
.Y(n_8550)
);

BUFx6f_ASAP7_75t_L g8551 ( 
.A(n_8046),
.Y(n_8551)
);

AOI21xp5_ASAP7_75t_L g8552 ( 
.A1(n_8408),
.A2(n_661),
.B(n_660),
.Y(n_8552)
);

OAI22xp5_ASAP7_75t_L g8553 ( 
.A1(n_8406),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_8553)
);

AOI21xp5_ASAP7_75t_L g8554 ( 
.A1(n_8416),
.A2(n_661),
.B(n_660),
.Y(n_8554)
);

NAND2xp5_ASAP7_75t_L g8555 ( 
.A(n_8412),
.B(n_662),
.Y(n_8555)
);

NAND2xp5_ASAP7_75t_L g8556 ( 
.A(n_8417),
.B(n_662),
.Y(n_8556)
);

INVx3_ASAP7_75t_L g8557 ( 
.A(n_7960),
.Y(n_8557)
);

AOI21x1_ASAP7_75t_L g8558 ( 
.A1(n_7942),
.A2(n_249),
.B(n_250),
.Y(n_8558)
);

OAI21x1_ASAP7_75t_L g8559 ( 
.A1(n_8248),
.A2(n_250),
.B(n_251),
.Y(n_8559)
);

NOR2xp33_ASAP7_75t_L g8560 ( 
.A(n_8386),
.B(n_663),
.Y(n_8560)
);

NOR2xp33_ASAP7_75t_L g8561 ( 
.A(n_8275),
.B(n_663),
.Y(n_8561)
);

NAND2xp5_ASAP7_75t_L g8562 ( 
.A(n_8425),
.B(n_8430),
.Y(n_8562)
);

BUFx2_ASAP7_75t_L g8563 ( 
.A(n_8359),
.Y(n_8563)
);

A2O1A1Ixp33_ASAP7_75t_L g8564 ( 
.A1(n_8175),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_8564)
);

AOI21xp5_ASAP7_75t_L g8565 ( 
.A1(n_8418),
.A2(n_665),
.B(n_664),
.Y(n_8565)
);

BUFx2_ASAP7_75t_L g8566 ( 
.A(n_7971),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_8152),
.Y(n_8567)
);

BUFx2_ASAP7_75t_L g8568 ( 
.A(n_8216),
.Y(n_8568)
);

NOR2xp33_ASAP7_75t_L g8569 ( 
.A(n_8179),
.B(n_666),
.Y(n_8569)
);

AOI21xp5_ASAP7_75t_L g8570 ( 
.A1(n_8420),
.A2(n_668),
.B(n_667),
.Y(n_8570)
);

INVxp67_ASAP7_75t_L g8571 ( 
.A(n_8140),
.Y(n_8571)
);

INVx4_ASAP7_75t_L g8572 ( 
.A(n_8046),
.Y(n_8572)
);

O2A1O1Ixp33_ASAP7_75t_L g8573 ( 
.A1(n_8456),
.A2(n_8381),
.B(n_8422),
.C(n_8384),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_8157),
.Y(n_8574)
);

NAND2xp5_ASAP7_75t_L g8575 ( 
.A(n_8434),
.B(n_668),
.Y(n_8575)
);

AOI21xp5_ASAP7_75t_L g8576 ( 
.A1(n_8426),
.A2(n_670),
.B(n_669),
.Y(n_8576)
);

OAI21xp5_ASAP7_75t_L g8577 ( 
.A1(n_8226),
.A2(n_251),
.B(n_252),
.Y(n_8577)
);

BUFx6f_ASAP7_75t_L g8578 ( 
.A(n_8046),
.Y(n_8578)
);

AOI21xp5_ASAP7_75t_L g8579 ( 
.A1(n_8432),
.A2(n_671),
.B(n_669),
.Y(n_8579)
);

OAI22xp5_ASAP7_75t_SL g8580 ( 
.A1(n_8222),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_8580)
);

NOR2xp33_ASAP7_75t_L g8581 ( 
.A(n_8185),
.B(n_8435),
.Y(n_8581)
);

AND2x4_ASAP7_75t_L g8582 ( 
.A(n_8409),
.B(n_671),
.Y(n_8582)
);

OAI22xp5_ASAP7_75t_L g8583 ( 
.A1(n_8441),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_8583)
);

NAND2xp5_ASAP7_75t_SL g8584 ( 
.A(n_8187),
.B(n_672),
.Y(n_8584)
);

NAND2xp5_ASAP7_75t_SL g8585 ( 
.A(n_7970),
.B(n_673),
.Y(n_8585)
);

INVx1_ASAP7_75t_L g8586 ( 
.A(n_8188),
.Y(n_8586)
);

AOI21xp5_ASAP7_75t_L g8587 ( 
.A1(n_8436),
.A2(n_8460),
.B(n_8439),
.Y(n_8587)
);

AOI21x1_ASAP7_75t_L g8588 ( 
.A1(n_7947),
.A2(n_253),
.B(n_254),
.Y(n_8588)
);

BUFx3_ASAP7_75t_L g8589 ( 
.A(n_8258),
.Y(n_8589)
);

NAND3xp33_ASAP7_75t_SL g8590 ( 
.A(n_8054),
.B(n_255),
.C(n_256),
.Y(n_8590)
);

OR2x6_ASAP7_75t_SL g8591 ( 
.A(n_8442),
.B(n_255),
.Y(n_8591)
);

NOR2xp33_ASAP7_75t_R g8592 ( 
.A(n_7975),
.B(n_255),
.Y(n_8592)
);

AND2x2_ASAP7_75t_L g8593 ( 
.A(n_8182),
.B(n_673),
.Y(n_8593)
);

NAND2xp5_ASAP7_75t_SL g8594 ( 
.A(n_8038),
.B(n_674),
.Y(n_8594)
);

NAND3xp33_ASAP7_75t_L g8595 ( 
.A(n_8091),
.B(n_256),
.C(n_257),
.Y(n_8595)
);

NAND2xp5_ASAP7_75t_L g8596 ( 
.A(n_8453),
.B(n_676),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_8455),
.B(n_676),
.Y(n_8597)
);

NAND2xp5_ASAP7_75t_L g8598 ( 
.A(n_8459),
.B(n_677),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_8190),
.Y(n_8599)
);

OAI22xp5_ASAP7_75t_L g8600 ( 
.A1(n_7939),
.A2(n_260),
.B1(n_257),
.B2(n_258),
.Y(n_8600)
);

AOI21xp5_ASAP7_75t_L g8601 ( 
.A1(n_8061),
.A2(n_678),
.B(n_677),
.Y(n_8601)
);

AOI21xp5_ASAP7_75t_L g8602 ( 
.A1(n_8224),
.A2(n_679),
.B(n_678),
.Y(n_8602)
);

NOR2xp33_ASAP7_75t_L g8603 ( 
.A(n_8306),
.B(n_679),
.Y(n_8603)
);

INVx2_ASAP7_75t_L g8604 ( 
.A(n_8419),
.Y(n_8604)
);

NAND2xp5_ASAP7_75t_SL g8605 ( 
.A(n_8461),
.B(n_680),
.Y(n_8605)
);

BUFx6f_ASAP7_75t_L g8606 ( 
.A(n_8139),
.Y(n_8606)
);

O2A1O1Ixp33_ASAP7_75t_L g8607 ( 
.A1(n_8437),
.A2(n_261),
.B(n_258),
.C(n_260),
.Y(n_8607)
);

OAI22xp5_ASAP7_75t_L g8608 ( 
.A1(n_8090),
.A2(n_261),
.B1(n_258),
.B2(n_260),
.Y(n_8608)
);

BUFx2_ASAP7_75t_L g8609 ( 
.A(n_8375),
.Y(n_8609)
);

AOI21xp5_ASAP7_75t_L g8610 ( 
.A1(n_8172),
.A2(n_682),
.B(n_681),
.Y(n_8610)
);

NAND2xp5_ASAP7_75t_L g8611 ( 
.A(n_8101),
.B(n_681),
.Y(n_8611)
);

NAND2xp5_ASAP7_75t_L g8612 ( 
.A(n_8383),
.B(n_682),
.Y(n_8612)
);

INVxp67_ASAP7_75t_L g8613 ( 
.A(n_8263),
.Y(n_8613)
);

O2A1O1Ixp33_ASAP7_75t_L g8614 ( 
.A1(n_8446),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_8614)
);

AOI21xp5_ASAP7_75t_L g8615 ( 
.A1(n_8130),
.A2(n_684),
.B(n_683),
.Y(n_8615)
);

AOI21xp5_ASAP7_75t_L g8616 ( 
.A1(n_8033),
.A2(n_684),
.B(n_683),
.Y(n_8616)
);

AND2x4_ASAP7_75t_L g8617 ( 
.A(n_8296),
.B(n_685),
.Y(n_8617)
);

NAND2xp5_ASAP7_75t_SL g8618 ( 
.A(n_8164),
.B(n_686),
.Y(n_8618)
);

AND2x2_ASAP7_75t_L g8619 ( 
.A(n_8376),
.B(n_8305),
.Y(n_8619)
);

OAI22xp5_ASAP7_75t_L g8620 ( 
.A1(n_8112),
.A2(n_8127),
.B1(n_7973),
.B2(n_8081),
.Y(n_8620)
);

AOI22xp5_ASAP7_75t_L g8621 ( 
.A1(n_7976),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_8194),
.Y(n_8622)
);

NAND2x1_ASAP7_75t_L g8623 ( 
.A(n_8115),
.B(n_687),
.Y(n_8623)
);

NOR3xp33_ASAP7_75t_SL g8624 ( 
.A(n_8118),
.B(n_262),
.C(n_263),
.Y(n_8624)
);

AND2x2_ASAP7_75t_L g8625 ( 
.A(n_8267),
.B(n_687),
.Y(n_8625)
);

NOR2xp33_ASAP7_75t_SL g8626 ( 
.A(n_8196),
.B(n_264),
.Y(n_8626)
);

NOR2xp33_ASAP7_75t_SL g8627 ( 
.A(n_8464),
.B(n_264),
.Y(n_8627)
);

AOI21xp5_ASAP7_75t_L g8628 ( 
.A1(n_8221),
.A2(n_689),
.B(n_688),
.Y(n_8628)
);

AOI22x1_ASAP7_75t_L g8629 ( 
.A1(n_8213),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_8629)
);

AND2x2_ASAP7_75t_L g8630 ( 
.A(n_8193),
.B(n_690),
.Y(n_8630)
);

AO21x1_ASAP7_75t_L g8631 ( 
.A1(n_8319),
.A2(n_265),
.B(n_266),
.Y(n_8631)
);

AND2x4_ASAP7_75t_L g8632 ( 
.A(n_8064),
.B(n_691),
.Y(n_8632)
);

AOI21xp5_ASAP7_75t_L g8633 ( 
.A1(n_8286),
.A2(n_692),
.B(n_691),
.Y(n_8633)
);

INVx2_ASAP7_75t_L g8634 ( 
.A(n_8424),
.Y(n_8634)
);

INVx2_ASAP7_75t_L g8635 ( 
.A(n_8438),
.Y(n_8635)
);

INVx1_ASAP7_75t_L g8636 ( 
.A(n_8195),
.Y(n_8636)
);

AOI21xp5_ASAP7_75t_L g8637 ( 
.A1(n_8215),
.A2(n_693),
.B(n_692),
.Y(n_8637)
);

A2O1A1Ixp33_ASAP7_75t_L g8638 ( 
.A1(n_8092),
.A2(n_695),
.B(n_696),
.C(n_694),
.Y(n_8638)
);

INVx6_ASAP7_75t_L g8639 ( 
.A(n_8139),
.Y(n_8639)
);

AND2x2_ASAP7_75t_L g8640 ( 
.A(n_8246),
.B(n_694),
.Y(n_8640)
);

OAI22xp5_ASAP7_75t_L g8641 ( 
.A1(n_8458),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_8641)
);

AND2x4_ASAP7_75t_L g8642 ( 
.A(n_8142),
.B(n_695),
.Y(n_8642)
);

NAND2xp5_ASAP7_75t_L g8643 ( 
.A(n_8450),
.B(n_696),
.Y(n_8643)
);

O2A1O1Ixp5_ASAP7_75t_L g8644 ( 
.A1(n_8285),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_SL g8645 ( 
.A(n_7957),
.B(n_697),
.Y(n_8645)
);

NOR2xp33_ASAP7_75t_L g8646 ( 
.A(n_8018),
.B(n_698),
.Y(n_8646)
);

AOI21xp5_ASAP7_75t_L g8647 ( 
.A1(n_8348),
.A2(n_700),
.B(n_699),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8206),
.Y(n_8648)
);

BUFx6f_ASAP7_75t_L g8649 ( 
.A(n_8111),
.Y(n_8649)
);

NAND2xp5_ASAP7_75t_L g8650 ( 
.A(n_8096),
.B(n_700),
.Y(n_8650)
);

NAND2xp5_ASAP7_75t_L g8651 ( 
.A(n_8211),
.B(n_701),
.Y(n_8651)
);

OAI221xp5_ASAP7_75t_L g8652 ( 
.A1(n_8223),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.C(n_271),
.Y(n_8652)
);

BUFx12f_ASAP7_75t_L g8653 ( 
.A(n_8289),
.Y(n_8653)
);

INVx1_ASAP7_75t_L g8654 ( 
.A(n_8207),
.Y(n_8654)
);

OR2x6_ASAP7_75t_L g8655 ( 
.A(n_7963),
.B(n_702),
.Y(n_8655)
);

AOI22xp33_ASAP7_75t_L g8656 ( 
.A1(n_8089),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_8656)
);

NAND2xp5_ASAP7_75t_L g8657 ( 
.A(n_7997),
.B(n_7952),
.Y(n_8657)
);

CKINVDCx20_ASAP7_75t_R g8658 ( 
.A(n_8368),
.Y(n_8658)
);

NAND2xp5_ASAP7_75t_L g8659 ( 
.A(n_7966),
.B(n_703),
.Y(n_8659)
);

INVx2_ASAP7_75t_L g8660 ( 
.A(n_8334),
.Y(n_8660)
);

BUFx6f_ASAP7_75t_L g8661 ( 
.A(n_8111),
.Y(n_8661)
);

NAND3xp33_ASAP7_75t_SL g8662 ( 
.A(n_8028),
.B(n_271),
.C(n_272),
.Y(n_8662)
);

OAI21xp5_ASAP7_75t_L g8663 ( 
.A1(n_8204),
.A2(n_272),
.B(n_273),
.Y(n_8663)
);

INVx2_ASAP7_75t_L g8664 ( 
.A(n_8145),
.Y(n_8664)
);

AOI21xp5_ASAP7_75t_L g8665 ( 
.A1(n_8108),
.A2(n_705),
.B(n_704),
.Y(n_8665)
);

O2A1O1Ixp33_ASAP7_75t_L g8666 ( 
.A1(n_7969),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_8666)
);

OAI22xp5_ASAP7_75t_L g8667 ( 
.A1(n_8427),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_8667)
);

NAND2xp5_ASAP7_75t_SL g8668 ( 
.A(n_8143),
.B(n_704),
.Y(n_8668)
);

AOI21xp5_ASAP7_75t_L g8669 ( 
.A1(n_8066),
.A2(n_706),
.B(n_705),
.Y(n_8669)
);

AOI22xp33_ASAP7_75t_L g8670 ( 
.A1(n_8252),
.A2(n_280),
.B1(n_276),
.B2(n_279),
.Y(n_8670)
);

NAND2xp5_ASAP7_75t_SL g8671 ( 
.A(n_8264),
.B(n_8280),
.Y(n_8671)
);

NOR2xp33_ASAP7_75t_L g8672 ( 
.A(n_8308),
.B(n_706),
.Y(n_8672)
);

OR2x2_ASAP7_75t_L g8673 ( 
.A(n_8349),
.B(n_707),
.Y(n_8673)
);

NAND2xp5_ASAP7_75t_L g8674 ( 
.A(n_7972),
.B(n_708),
.Y(n_8674)
);

A2O1A1Ixp33_ASAP7_75t_L g8675 ( 
.A1(n_8138),
.A2(n_709),
.B(n_710),
.C(n_708),
.Y(n_8675)
);

NAND2x1p5_ASAP7_75t_L g8676 ( 
.A(n_8105),
.B(n_709),
.Y(n_8676)
);

OAI21xp5_ASAP7_75t_L g8677 ( 
.A1(n_8173),
.A2(n_279),
.B(n_280),
.Y(n_8677)
);

AOI21xp5_ASAP7_75t_L g8678 ( 
.A1(n_8239),
.A2(n_712),
.B(n_711),
.Y(n_8678)
);

AOI21x1_ASAP7_75t_L g8679 ( 
.A1(n_7961),
.A2(n_279),
.B(n_281),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8146),
.Y(n_8680)
);

OAI22xp5_ASAP7_75t_L g8681 ( 
.A1(n_8203),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_8681)
);

O2A1O1Ixp33_ASAP7_75t_L g8682 ( 
.A1(n_8074),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_8682)
);

AND2x2_ASAP7_75t_L g8683 ( 
.A(n_8247),
.B(n_712),
.Y(n_8683)
);

INVx2_ASAP7_75t_L g8684 ( 
.A(n_8261),
.Y(n_8684)
);

INVx2_ASAP7_75t_L g8685 ( 
.A(n_8281),
.Y(n_8685)
);

NAND2xp5_ASAP7_75t_L g8686 ( 
.A(n_8380),
.B(n_713),
.Y(n_8686)
);

AND2x4_ASAP7_75t_L g8687 ( 
.A(n_8170),
.B(n_713),
.Y(n_8687)
);

INVx2_ASAP7_75t_L g8688 ( 
.A(n_8078),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_8276),
.Y(n_8689)
);

AO22x1_ASAP7_75t_L g8690 ( 
.A1(n_8323),
.A2(n_8354),
.B1(n_8312),
.B2(n_7993),
.Y(n_8690)
);

INVx2_ASAP7_75t_L g8691 ( 
.A(n_8208),
.Y(n_8691)
);

AOI21xp5_ASAP7_75t_L g8692 ( 
.A1(n_8086),
.A2(n_715),
.B(n_714),
.Y(n_8692)
);

BUFx6f_ASAP7_75t_L g8693 ( 
.A(n_8467),
.Y(n_8693)
);

NOR2xp33_ASAP7_75t_L g8694 ( 
.A(n_8021),
.B(n_714),
.Y(n_8694)
);

AOI21xp5_ASAP7_75t_L g8695 ( 
.A1(n_8088),
.A2(n_717),
.B(n_716),
.Y(n_8695)
);

BUFx8_ASAP7_75t_SL g8696 ( 
.A(n_8307),
.Y(n_8696)
);

BUFx2_ASAP7_75t_L g8697 ( 
.A(n_8210),
.Y(n_8697)
);

INVx1_ASAP7_75t_L g8698 ( 
.A(n_8316),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_L g8699 ( 
.A(n_8388),
.B(n_716),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8317),
.Y(n_8700)
);

NAND2xp5_ASAP7_75t_SL g8701 ( 
.A(n_8197),
.B(n_718),
.Y(n_8701)
);

AOI21xp5_ASAP7_75t_L g8702 ( 
.A1(n_8156),
.A2(n_719),
.B(n_718),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_8413),
.Y(n_8703)
);

INVx3_ASAP7_75t_L g8704 ( 
.A(n_8019),
.Y(n_8704)
);

OAI21xp5_ASAP7_75t_L g8705 ( 
.A1(n_8120),
.A2(n_282),
.B(n_284),
.Y(n_8705)
);

NAND2xp5_ASAP7_75t_L g8706 ( 
.A(n_8423),
.B(n_720),
.Y(n_8706)
);

INVx2_ASAP7_75t_SL g8707 ( 
.A(n_7994),
.Y(n_8707)
);

NOR2xp33_ASAP7_75t_L g8708 ( 
.A(n_8149),
.B(n_720),
.Y(n_8708)
);

O2A1O1Ixp33_ASAP7_75t_L g8709 ( 
.A1(n_8244),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_8709)
);

O2A1O1Ixp33_ASAP7_75t_L g8710 ( 
.A1(n_8433),
.A2(n_288),
.B(n_285),
.C(n_287),
.Y(n_8710)
);

INVxp67_ASAP7_75t_L g8711 ( 
.A(n_8097),
.Y(n_8711)
);

HB1xp67_ASAP7_75t_L g8712 ( 
.A(n_8428),
.Y(n_8712)
);

AOI21xp5_ASAP7_75t_L g8713 ( 
.A1(n_8220),
.A2(n_722),
.B(n_721),
.Y(n_8713)
);

NAND2xp5_ASAP7_75t_SL g8714 ( 
.A(n_8303),
.B(n_722),
.Y(n_8714)
);

O2A1O1Ixp33_ASAP7_75t_L g8715 ( 
.A1(n_8448),
.A2(n_288),
.B(n_285),
.C(n_287),
.Y(n_8715)
);

OR2x6_ASAP7_75t_L g8716 ( 
.A(n_7963),
.B(n_724),
.Y(n_8716)
);

A2O1A1Ixp33_ASAP7_75t_L g8717 ( 
.A1(n_8273),
.A2(n_726),
.B(n_727),
.C(n_725),
.Y(n_8717)
);

O2A1O1Ixp33_ASAP7_75t_L g8718 ( 
.A1(n_8265),
.A2(n_290),
.B(n_288),
.C(n_289),
.Y(n_8718)
);

NAND2xp5_ASAP7_75t_L g8719 ( 
.A(n_8219),
.B(n_8245),
.Y(n_8719)
);

INVx2_ASAP7_75t_L g8720 ( 
.A(n_8217),
.Y(n_8720)
);

AOI21xp5_ASAP7_75t_L g8721 ( 
.A1(n_8220),
.A2(n_8236),
.B(n_7937),
.Y(n_8721)
);

O2A1O1Ixp5_ASAP7_75t_L g8722 ( 
.A1(n_8294),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_8722)
);

NAND2xp5_ASAP7_75t_SL g8723 ( 
.A(n_8014),
.B(n_725),
.Y(n_8723)
);

NAND2xp5_ASAP7_75t_L g8724 ( 
.A(n_8004),
.B(n_726),
.Y(n_8724)
);

AOI22xp33_ASAP7_75t_L g8725 ( 
.A1(n_8184),
.A2(n_292),
.B1(n_289),
.B2(n_291),
.Y(n_8725)
);

INVx3_ASAP7_75t_SL g8726 ( 
.A(n_8431),
.Y(n_8726)
);

NOR2xp33_ASAP7_75t_L g8727 ( 
.A(n_8339),
.B(n_727),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_8321),
.Y(n_8728)
);

INVx2_ASAP7_75t_L g8729 ( 
.A(n_8026),
.Y(n_8729)
);

BUFx6f_ASAP7_75t_L g8730 ( 
.A(n_8431),
.Y(n_8730)
);

OAI21xp5_ASAP7_75t_L g8731 ( 
.A1(n_8268),
.A2(n_292),
.B(n_293),
.Y(n_8731)
);

HB1xp67_ASAP7_75t_L g8732 ( 
.A(n_8335),
.Y(n_8732)
);

INVx4_ASAP7_75t_L g8733 ( 
.A(n_8278),
.Y(n_8733)
);

NAND2xp5_ASAP7_75t_L g8734 ( 
.A(n_8056),
.B(n_728),
.Y(n_8734)
);

AOI22xp33_ASAP7_75t_L g8735 ( 
.A1(n_8075),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_8735)
);

NOR3xp33_ASAP7_75t_SL g8736 ( 
.A(n_8128),
.B(n_295),
.C(n_296),
.Y(n_8736)
);

AND2x2_ASAP7_75t_L g8737 ( 
.A(n_8353),
.B(n_728),
.Y(n_8737)
);

INVx2_ASAP7_75t_L g8738 ( 
.A(n_8058),
.Y(n_8738)
);

NOR2x1_ASAP7_75t_R g8739 ( 
.A(n_7929),
.B(n_296),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_8325),
.Y(n_8740)
);

AOI21xp5_ASAP7_75t_L g8741 ( 
.A1(n_7936),
.A2(n_731),
.B(n_730),
.Y(n_8741)
);

OAI22xp5_ASAP7_75t_L g8742 ( 
.A1(n_8350),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_8328),
.Y(n_8743)
);

NAND2x1p5_ASAP7_75t_L g8744 ( 
.A(n_8137),
.B(n_730),
.Y(n_8744)
);

INVx1_ASAP7_75t_L g8745 ( 
.A(n_8327),
.Y(n_8745)
);

AOI221xp5_ASAP7_75t_L g8746 ( 
.A1(n_8271),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.C(n_300),
.Y(n_8746)
);

AOI21xp5_ASAP7_75t_L g8747 ( 
.A1(n_8468),
.A2(n_733),
.B(n_731),
.Y(n_8747)
);

INVx2_ASAP7_75t_L g8748 ( 
.A(n_8270),
.Y(n_8748)
);

A2O1A1Ixp33_ASAP7_75t_L g8749 ( 
.A1(n_8147),
.A2(n_8167),
.B(n_8155),
.C(n_8249),
.Y(n_8749)
);

AOI21xp5_ASAP7_75t_L g8750 ( 
.A1(n_8396),
.A2(n_735),
.B(n_734),
.Y(n_8750)
);

INVx1_ASAP7_75t_L g8751 ( 
.A(n_8466),
.Y(n_8751)
);

AOI21xp33_ASAP7_75t_L g8752 ( 
.A1(n_8043),
.A2(n_297),
.B(n_298),
.Y(n_8752)
);

NOR2xp33_ASAP7_75t_R g8753 ( 
.A(n_8141),
.B(n_299),
.Y(n_8753)
);

INVx2_ASAP7_75t_L g8754 ( 
.A(n_8218),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_8360),
.Y(n_8755)
);

INVx1_ASAP7_75t_L g8756 ( 
.A(n_8364),
.Y(n_8756)
);

OR2x2_ASAP7_75t_L g8757 ( 
.A(n_8272),
.B(n_734),
.Y(n_8757)
);

BUFx2_ASAP7_75t_L g8758 ( 
.A(n_8358),
.Y(n_8758)
);

BUFx4f_ASAP7_75t_L g8759 ( 
.A(n_8293),
.Y(n_8759)
);

NAND2xp5_ASAP7_75t_L g8760 ( 
.A(n_8063),
.B(n_735),
.Y(n_8760)
);

AOI21xp5_ASAP7_75t_L g8761 ( 
.A1(n_8415),
.A2(n_737),
.B(n_736),
.Y(n_8761)
);

INVx2_ASAP7_75t_SL g8762 ( 
.A(n_7992),
.Y(n_8762)
);

AOI21x1_ASAP7_75t_L g8763 ( 
.A1(n_8029),
.A2(n_299),
.B(n_300),
.Y(n_8763)
);

AOI21xp5_ASAP7_75t_L g8764 ( 
.A1(n_8073),
.A2(n_738),
.B(n_737),
.Y(n_8764)
);

OAI22xp5_ASAP7_75t_L g8765 ( 
.A1(n_8287),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_8765)
);

A2O1A1Ixp33_ASAP7_75t_L g8766 ( 
.A1(n_8107),
.A2(n_739),
.B(n_740),
.C(n_738),
.Y(n_8766)
);

AOI21xp5_ASAP7_75t_L g8767 ( 
.A1(n_8077),
.A2(n_741),
.B(n_740),
.Y(n_8767)
);

INVx4_ASAP7_75t_L g8768 ( 
.A(n_8282),
.Y(n_8768)
);

NOR2xp33_ASAP7_75t_L g8769 ( 
.A(n_8374),
.B(n_741),
.Y(n_8769)
);

OAI22xp5_ASAP7_75t_L g8770 ( 
.A1(n_8371),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_8770)
);

INVx3_ASAP7_75t_L g8771 ( 
.A(n_8189),
.Y(n_8771)
);

NOR2xp33_ASAP7_75t_L g8772 ( 
.A(n_8314),
.B(n_742),
.Y(n_8772)
);

BUFx2_ASAP7_75t_L g8773 ( 
.A(n_8150),
.Y(n_8773)
);

INVx2_ASAP7_75t_L g8774 ( 
.A(n_8104),
.Y(n_8774)
);

NAND2xp5_ASAP7_75t_L g8775 ( 
.A(n_7943),
.B(n_743),
.Y(n_8775)
);

HB1xp67_ASAP7_75t_L g8776 ( 
.A(n_8109),
.Y(n_8776)
);

INVx4_ASAP7_75t_L g8777 ( 
.A(n_8022),
.Y(n_8777)
);

INVx2_ASAP7_75t_L g8778 ( 
.A(n_8209),
.Y(n_8778)
);

INVx2_ASAP7_75t_L g8779 ( 
.A(n_8231),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_SL g8780 ( 
.A(n_8049),
.B(n_743),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_8233),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_L g8782 ( 
.A(n_8048),
.B(n_744),
.Y(n_8782)
);

XNOR2xp5_ASAP7_75t_L g8783 ( 
.A(n_8377),
.B(n_301),
.Y(n_8783)
);

AOI21xp5_ASAP7_75t_L g8784 ( 
.A1(n_7944),
.A2(n_8010),
.B(n_8008),
.Y(n_8784)
);

NAND2xp5_ASAP7_75t_SL g8785 ( 
.A(n_8168),
.B(n_744),
.Y(n_8785)
);

INVx2_ASAP7_75t_L g8786 ( 
.A(n_8242),
.Y(n_8786)
);

O2A1O1Ixp33_ASAP7_75t_L g8787 ( 
.A1(n_8326),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_8787)
);

AND2x2_ASAP7_75t_L g8788 ( 
.A(n_8330),
.B(n_745),
.Y(n_8788)
);

BUFx2_ASAP7_75t_L g8789 ( 
.A(n_8309),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_7959),
.B(n_745),
.Y(n_8790)
);

NOR2xp33_ASAP7_75t_L g8791 ( 
.A(n_8315),
.B(n_746),
.Y(n_8791)
);

INVx1_ASAP7_75t_L g8792 ( 
.A(n_8060),
.Y(n_8792)
);

OAI22xp5_ASAP7_75t_L g8793 ( 
.A1(n_8259),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_8793)
);

HB1xp67_ASAP7_75t_L g8794 ( 
.A(n_8023),
.Y(n_8794)
);

BUFx6f_ASAP7_75t_L g8795 ( 
.A(n_8230),
.Y(n_8795)
);

NOR2xp33_ASAP7_75t_L g8796 ( 
.A(n_8166),
.B(n_746),
.Y(n_8796)
);

NAND2xp5_ASAP7_75t_SL g8797 ( 
.A(n_8329),
.B(n_747),
.Y(n_8797)
);

INVx1_ASAP7_75t_L g8798 ( 
.A(n_8069),
.Y(n_8798)
);

NAND2xp5_ASAP7_75t_L g8799 ( 
.A(n_7978),
.B(n_747),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_8198),
.Y(n_8800)
);

NAND2xp5_ASAP7_75t_L g8801 ( 
.A(n_7999),
.B(n_748),
.Y(n_8801)
);

INVx1_ASAP7_75t_L g8802 ( 
.A(n_8331),
.Y(n_8802)
);

BUFx2_ASAP7_75t_R g8803 ( 
.A(n_8336),
.Y(n_8803)
);

NAND2xp5_ASAP7_75t_L g8804 ( 
.A(n_8016),
.B(n_748),
.Y(n_8804)
);

INVx2_ASAP7_75t_L g8805 ( 
.A(n_8159),
.Y(n_8805)
);

NOR2xp33_ASAP7_75t_L g8806 ( 
.A(n_8297),
.B(n_749),
.Y(n_8806)
);

BUFx12f_ASAP7_75t_L g8807 ( 
.A(n_8452),
.Y(n_8807)
);

AOI21xp5_ASAP7_75t_L g8808 ( 
.A1(n_8052),
.A2(n_751),
.B(n_750),
.Y(n_8808)
);

INVx1_ASAP7_75t_L g8809 ( 
.A(n_8344),
.Y(n_8809)
);

INVx5_ASAP7_75t_L g8810 ( 
.A(n_8354),
.Y(n_8810)
);

BUFx3_ASAP7_75t_L g8811 ( 
.A(n_8295),
.Y(n_8811)
);

AOI22xp5_ASAP7_75t_L g8812 ( 
.A1(n_8068),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_SL g8813 ( 
.A(n_7941),
.B(n_750),
.Y(n_8813)
);

INVx1_ASAP7_75t_L g8814 ( 
.A(n_8067),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8055),
.Y(n_8815)
);

INVx3_ASAP7_75t_L g8816 ( 
.A(n_8367),
.Y(n_8816)
);

AOI21xp5_ASAP7_75t_L g8817 ( 
.A1(n_8071),
.A2(n_752),
.B(n_751),
.Y(n_8817)
);

AOI21xp5_ASAP7_75t_L g8818 ( 
.A1(n_8202),
.A2(n_754),
.B(n_753),
.Y(n_8818)
);

AND2x4_ASAP7_75t_L g8819 ( 
.A(n_8355),
.B(n_753),
.Y(n_8819)
);

OR2x6_ASAP7_75t_L g8820 ( 
.A(n_8372),
.B(n_755),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_SL g8821 ( 
.A(n_8411),
.B(n_755),
.Y(n_8821)
);

INVx3_ASAP7_75t_L g8822 ( 
.A(n_8393),
.Y(n_8822)
);

INVx3_ASAP7_75t_SL g8823 ( 
.A(n_8414),
.Y(n_8823)
);

A2O1A1Ixp33_ASAP7_75t_L g8824 ( 
.A1(n_8113),
.A2(n_8122),
.B(n_7951),
.C(n_8020),
.Y(n_8824)
);

NOR2xp33_ASAP7_75t_L g8825 ( 
.A(n_8298),
.B(n_756),
.Y(n_8825)
);

OAI22xp5_ASAP7_75t_L g8826 ( 
.A1(n_7974),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_8826)
);

A2O1A1Ixp33_ASAP7_75t_L g8827 ( 
.A1(n_8369),
.A2(n_757),
.B(n_758),
.C(n_756),
.Y(n_8827)
);

OAI22xp5_ASAP7_75t_L g8828 ( 
.A1(n_8324),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_8828)
);

NOR2xp33_ASAP7_75t_L g8829 ( 
.A(n_8253),
.B(n_757),
.Y(n_8829)
);

NOR2xp33_ASAP7_75t_L g8830 ( 
.A(n_8257),
.B(n_758),
.Y(n_8830)
);

INVx2_ASAP7_75t_L g8831 ( 
.A(n_8057),
.Y(n_8831)
);

BUFx4f_ASAP7_75t_L g8832 ( 
.A(n_8421),
.Y(n_8832)
);

INVx1_ASAP7_75t_L g8833 ( 
.A(n_8161),
.Y(n_8833)
);

AOI21xp5_ASAP7_75t_L g8834 ( 
.A1(n_8125),
.A2(n_760),
.B(n_759),
.Y(n_8834)
);

AOI21xp5_ASAP7_75t_L g8835 ( 
.A1(n_8126),
.A2(n_760),
.B(n_759),
.Y(n_8835)
);

INVx3_ASAP7_75t_L g8836 ( 
.A(n_8451),
.Y(n_8836)
);

CKINVDCx10_ASAP7_75t_R g8837 ( 
.A(n_8345),
.Y(n_8837)
);

NAND2xp5_ASAP7_75t_L g8838 ( 
.A(n_7946),
.B(n_761),
.Y(n_8838)
);

NOR2xp67_ASAP7_75t_L g8839 ( 
.A(n_7958),
.B(n_308),
.Y(n_8839)
);

AND2x2_ASAP7_75t_L g8840 ( 
.A(n_8160),
.B(n_762),
.Y(n_8840)
);

NAND2xp5_ASAP7_75t_L g8841 ( 
.A(n_7965),
.B(n_762),
.Y(n_8841)
);

OR2x2_ASAP7_75t_L g8842 ( 
.A(n_7982),
.B(n_763),
.Y(n_8842)
);

O2A1O1Ixp33_ASAP7_75t_L g8843 ( 
.A1(n_7979),
.A2(n_312),
.B(n_309),
.C(n_311),
.Y(n_8843)
);

AND2x4_ASAP7_75t_L g8844 ( 
.A(n_8469),
.B(n_763),
.Y(n_8844)
);

HB1xp67_ASAP7_75t_L g8845 ( 
.A(n_8171),
.Y(n_8845)
);

NAND2xp5_ASAP7_75t_SL g8846 ( 
.A(n_8176),
.B(n_764),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_7989),
.Y(n_8847)
);

CKINVDCx14_ASAP7_75t_R g8848 ( 
.A(n_8131),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_7996),
.Y(n_8849)
);

NOR2xp33_ASAP7_75t_L g8850 ( 
.A(n_8341),
.B(n_765),
.Y(n_8850)
);

AOI21xp5_ASAP7_75t_L g8851 ( 
.A1(n_8144),
.A2(n_767),
.B(n_766),
.Y(n_8851)
);

INVx1_ASAP7_75t_L g8852 ( 
.A(n_8000),
.Y(n_8852)
);

AO31x2_ASAP7_75t_L g8853 ( 
.A1(n_8031),
.A2(n_313),
.A3(n_311),
.B(n_312),
.Y(n_8853)
);

NOR2xp33_ASAP7_75t_SL g8854 ( 
.A(n_8291),
.B(n_311),
.Y(n_8854)
);

INVx2_ASAP7_75t_L g8855 ( 
.A(n_8001),
.Y(n_8855)
);

O2A1O1Ixp33_ASAP7_75t_L g8856 ( 
.A1(n_8009),
.A2(n_315),
.B(n_312),
.C(n_314),
.Y(n_8856)
);

INVx1_ASAP7_75t_L g8857 ( 
.A(n_8011),
.Y(n_8857)
);

INVx2_ASAP7_75t_L g8858 ( 
.A(n_8012),
.Y(n_8858)
);

HB1xp67_ASAP7_75t_L g8859 ( 
.A(n_8098),
.Y(n_8859)
);

OAI22xp5_ASAP7_75t_L g8860 ( 
.A1(n_8045),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_8860)
);

CKINVDCx5p33_ASAP7_75t_R g8861 ( 
.A(n_8225),
.Y(n_8861)
);

NAND2xp5_ASAP7_75t_L g8862 ( 
.A(n_8024),
.B(n_767),
.Y(n_8862)
);

NAND2xp5_ASAP7_75t_SL g8863 ( 
.A(n_8200),
.B(n_768),
.Y(n_8863)
);

A2O1A1Ixp33_ASAP7_75t_L g8864 ( 
.A1(n_8338),
.A2(n_771),
.B(n_772),
.C(n_768),
.Y(n_8864)
);

OAI22xp5_ASAP7_75t_L g8865 ( 
.A1(n_8347),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_8865)
);

AOI21xp5_ASAP7_75t_L g8866 ( 
.A1(n_8228),
.A2(n_772),
.B(n_771),
.Y(n_8866)
);

NAND2xp5_ASAP7_75t_SL g8867 ( 
.A(n_8214),
.B(n_773),
.Y(n_8867)
);

AND2x4_ASAP7_75t_L g8868 ( 
.A(n_8007),
.B(n_773),
.Y(n_8868)
);

INVx5_ASAP7_75t_L g8869 ( 
.A(n_8354),
.Y(n_8869)
);

AOI22xp5_ASAP7_75t_L g8870 ( 
.A1(n_8346),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_8870)
);

NOR2xp33_ASAP7_75t_R g8871 ( 
.A(n_8076),
.B(n_317),
.Y(n_8871)
);

O2A1O1Ixp33_ASAP7_75t_L g8872 ( 
.A1(n_8015),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_8872)
);

BUFx12f_ASAP7_75t_L g8873 ( 
.A(n_8235),
.Y(n_8873)
);

OAI22xp5_ASAP7_75t_L g8874 ( 
.A1(n_8351),
.A2(n_8227),
.B1(n_8229),
.B2(n_8135),
.Y(n_8874)
);

INVxp67_ASAP7_75t_L g8875 ( 
.A(n_8059),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_L g8876 ( 
.A(n_8027),
.B(n_774),
.Y(n_8876)
);

INVx3_ASAP7_75t_L g8877 ( 
.A(n_8301),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_SL g8878 ( 
.A(n_8082),
.B(n_774),
.Y(n_8878)
);

CKINVDCx14_ASAP7_75t_R g8879 ( 
.A(n_8310),
.Y(n_8879)
);

AND2x2_ASAP7_75t_L g8880 ( 
.A(n_8062),
.B(n_775),
.Y(n_8880)
);

INVx2_ASAP7_75t_L g8881 ( 
.A(n_8039),
.Y(n_8881)
);

OAI22xp5_ASAP7_75t_L g8882 ( 
.A1(n_8361),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_8882)
);

OAI22xp33_ASAP7_75t_L g8883 ( 
.A1(n_8260),
.A2(n_776),
.B1(n_777),
.B2(n_775),
.Y(n_8883)
);

INVx2_ASAP7_75t_L g8884 ( 
.A(n_8047),
.Y(n_8884)
);

OAI21xp5_ASAP7_75t_L g8885 ( 
.A1(n_7955),
.A2(n_321),
.B(n_322),
.Y(n_8885)
);

AOI21xp5_ASAP7_75t_L g8886 ( 
.A1(n_8266),
.A2(n_8153),
.B(n_8034),
.Y(n_8886)
);

CKINVDCx5p33_ASAP7_75t_R g8887 ( 
.A(n_8332),
.Y(n_8887)
);

NOR2xp33_ASAP7_75t_R g8888 ( 
.A(n_8050),
.B(n_321),
.Y(n_8888)
);

A2O1A1Ixp33_ASAP7_75t_L g8889 ( 
.A1(n_8407),
.A2(n_777),
.B(n_779),
.C(n_776),
.Y(n_8889)
);

NAND2xp5_ASAP7_75t_L g8890 ( 
.A(n_8051),
.B(n_779),
.Y(n_8890)
);

BUFx3_ASAP7_75t_L g8891 ( 
.A(n_8311),
.Y(n_8891)
);

AND2x2_ASAP7_75t_L g8892 ( 
.A(n_8399),
.B(n_780),
.Y(n_8892)
);

INVx4_ASAP7_75t_L g8893 ( 
.A(n_8447),
.Y(n_8893)
);

INVx2_ASAP7_75t_L g8894 ( 
.A(n_7949),
.Y(n_8894)
);

A2O1A1Ixp33_ASAP7_75t_L g8895 ( 
.A1(n_8080),
.A2(n_782),
.B(n_783),
.C(n_781),
.Y(n_8895)
);

AOI21xp5_ASAP7_75t_L g8896 ( 
.A1(n_8032),
.A2(n_8040),
.B(n_8035),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8181),
.Y(n_8897)
);

INVx1_ASAP7_75t_SL g8898 ( 
.A(n_8304),
.Y(n_8898)
);

NOR2xp33_ASAP7_75t_L g8899 ( 
.A(n_8151),
.B(n_781),
.Y(n_8899)
);

OAI22xp5_ASAP7_75t_L g8900 ( 
.A1(n_8041),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_8900)
);

AOI22xp33_ASAP7_75t_L g8901 ( 
.A1(n_8357),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_8901)
);

AND2x2_ASAP7_75t_L g8902 ( 
.A(n_8457),
.B(n_782),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_SL g8903 ( 
.A(n_8158),
.B(n_783),
.Y(n_8903)
);

O2A1O1Ixp33_ASAP7_75t_SL g8904 ( 
.A1(n_8114),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8178),
.B(n_8180),
.Y(n_8905)
);

INVx2_ASAP7_75t_L g8906 ( 
.A(n_7988),
.Y(n_8906)
);

HB1xp67_ASAP7_75t_L g8907 ( 
.A(n_8136),
.Y(n_8907)
);

OA21x2_ASAP7_75t_L g8908 ( 
.A1(n_8119),
.A2(n_325),
.B(n_326),
.Y(n_8908)
);

INVx1_ASAP7_75t_SL g8909 ( 
.A(n_8274),
.Y(n_8909)
);

HB1xp67_ASAP7_75t_L g8910 ( 
.A(n_8183),
.Y(n_8910)
);

NOR2xp33_ASAP7_75t_R g8911 ( 
.A(n_7953),
.B(n_325),
.Y(n_8911)
);

NAND2xp5_ASAP7_75t_L g8912 ( 
.A(n_8342),
.B(n_785),
.Y(n_8912)
);

NAND2xp5_ASAP7_75t_L g8913 ( 
.A(n_8322),
.B(n_785),
.Y(n_8913)
);

NAND2xp5_ASAP7_75t_L g8914 ( 
.A(n_8333),
.B(n_787),
.Y(n_8914)
);

NOR2xp33_ASAP7_75t_L g8915 ( 
.A(n_8162),
.B(n_787),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_SL g8916 ( 
.A(n_8163),
.B(n_788),
.Y(n_8916)
);

NAND2xp5_ASAP7_75t_L g8917 ( 
.A(n_8269),
.B(n_788),
.Y(n_8917)
);

INVx3_ASAP7_75t_L g8918 ( 
.A(n_8165),
.Y(n_8918)
);

NOR2xp33_ASAP7_75t_L g8919 ( 
.A(n_8124),
.B(n_8129),
.Y(n_8919)
);

NAND3xp33_ASAP7_75t_L g8920 ( 
.A(n_8084),
.B(n_326),
.C(n_327),
.Y(n_8920)
);

AOI21xp5_ASAP7_75t_L g8921 ( 
.A1(n_8044),
.A2(n_790),
.B(n_789),
.Y(n_8921)
);

OAI22xp5_ASAP7_75t_L g8922 ( 
.A1(n_8320),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_8922)
);

NOR2xp33_ASAP7_75t_L g8923 ( 
.A(n_8256),
.B(n_790),
.Y(n_8923)
);

NAND2xp5_ASAP7_75t_L g8924 ( 
.A(n_8255),
.B(n_791),
.Y(n_8924)
);

INVx2_ASAP7_75t_L g8925 ( 
.A(n_8262),
.Y(n_8925)
);

NAND2x1p5_ASAP7_75t_L g8926 ( 
.A(n_8037),
.B(n_792),
.Y(n_8926)
);

INVx3_ASAP7_75t_L g8927 ( 
.A(n_8337),
.Y(n_8927)
);

INVx2_ASAP7_75t_L g8928 ( 
.A(n_8340),
.Y(n_8928)
);

BUFx6f_ASAP7_75t_L g8929 ( 
.A(n_8363),
.Y(n_8929)
);

AND2x4_ASAP7_75t_L g8930 ( 
.A(n_8373),
.B(n_793),
.Y(n_8930)
);

A2O1A1Ixp33_ASAP7_75t_L g8931 ( 
.A1(n_7962),
.A2(n_795),
.B(n_796),
.C(n_793),
.Y(n_8931)
);

INVx3_ASAP7_75t_L g8932 ( 
.A(n_8370),
.Y(n_8932)
);

OAI22xp5_ASAP7_75t_L g8933 ( 
.A1(n_8362),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8277),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8318),
.B(n_795),
.Y(n_8935)
);

NAND2xp5_ASAP7_75t_L g8936 ( 
.A(n_8352),
.B(n_796),
.Y(n_8936)
);

INVx1_ASAP7_75t_SL g8937 ( 
.A(n_8103),
.Y(n_8937)
);

OAI22xp5_ASAP7_75t_L g8938 ( 
.A1(n_8379),
.A2(n_331),
.B1(n_328),
.B2(n_330),
.Y(n_8938)
);

OR2x2_ASAP7_75t_L g8939 ( 
.A(n_8365),
.B(n_8366),
.Y(n_8939)
);

NOR2xp33_ASAP7_75t_L g8940 ( 
.A(n_8087),
.B(n_797),
.Y(n_8940)
);

INVx3_ASAP7_75t_L g8941 ( 
.A(n_8465),
.Y(n_8941)
);

AOI21xp5_ASAP7_75t_L g8942 ( 
.A1(n_7977),
.A2(n_798),
.B(n_797),
.Y(n_8942)
);

INVx2_ASAP7_75t_L g8943 ( 
.A(n_8343),
.Y(n_8943)
);

NAND2xp5_ASAP7_75t_SL g8944 ( 
.A(n_8251),
.B(n_798),
.Y(n_8944)
);

NAND2xp5_ASAP7_75t_L g8945 ( 
.A(n_8356),
.B(n_799),
.Y(n_8945)
);

NAND2xp5_ASAP7_75t_L g8946 ( 
.A(n_8254),
.B(n_799),
.Y(n_8946)
);

INVx2_ASAP7_75t_L g8947 ( 
.A(n_8302),
.Y(n_8947)
);

INVx1_ASAP7_75t_L g8948 ( 
.A(n_8099),
.Y(n_8948)
);

INVx2_ASAP7_75t_SL g8949 ( 
.A(n_8036),
.Y(n_8949)
);

NAND2x1p5_ASAP7_75t_L g8950 ( 
.A(n_8300),
.B(n_800),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_SL g8951 ( 
.A(n_8083),
.B(n_802),
.Y(n_8951)
);

INVx2_ASAP7_75t_L g8952 ( 
.A(n_8288),
.Y(n_8952)
);

OAI22xp5_ASAP7_75t_L g8953 ( 
.A1(n_8391),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_8953)
);

INVx1_ASAP7_75t_L g8954 ( 
.A(n_8116),
.Y(n_8954)
);

INVx2_ASAP7_75t_L g8955 ( 
.A(n_7938),
.Y(n_8955)
);

NAND2xp5_ASAP7_75t_L g8956 ( 
.A(n_8440),
.B(n_8444),
.Y(n_8956)
);

INVx3_ASAP7_75t_L g8957 ( 
.A(n_8085),
.Y(n_8957)
);

INVx3_ASAP7_75t_L g8958 ( 
.A(n_8378),
.Y(n_8958)
);

AND2x2_ASAP7_75t_L g8959 ( 
.A(n_7980),
.B(n_802),
.Y(n_8959)
);

NAND2xp5_ASAP7_75t_SL g8960 ( 
.A(n_8445),
.B(n_803),
.Y(n_8960)
);

BUFx2_ASAP7_75t_L g8961 ( 
.A(n_8283),
.Y(n_8961)
);

AO22x1_ASAP7_75t_L g8962 ( 
.A1(n_7985),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_8962)
);

HB1xp67_ASAP7_75t_L g8963 ( 
.A(n_8284),
.Y(n_8963)
);

INVxp67_ASAP7_75t_L g8964 ( 
.A(n_7987),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8292),
.Y(n_8965)
);

NAND2xp5_ASAP7_75t_SL g8966 ( 
.A(n_7998),
.B(n_803),
.Y(n_8966)
);

AOI21xp5_ASAP7_75t_L g8967 ( 
.A1(n_8003),
.A2(n_805),
.B(n_804),
.Y(n_8967)
);

NAND2xp5_ASAP7_75t_SL g8968 ( 
.A(n_8299),
.B(n_805),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_SL g8969 ( 
.A(n_8205),
.B(n_806),
.Y(n_8969)
);

OAI22xp5_ASAP7_75t_L g8970 ( 
.A1(n_8174),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_8970)
);

INVx1_ASAP7_75t_SL g8971 ( 
.A(n_8232),
.Y(n_8971)
);

NAND2xp5_ASAP7_75t_L g8972 ( 
.A(n_8212),
.B(n_8191),
.Y(n_8972)
);

NOR2xp33_ASAP7_75t_L g8973 ( 
.A(n_8237),
.B(n_807),
.Y(n_8973)
);

A2O1A1Ixp33_ASAP7_75t_L g8974 ( 
.A1(n_8192),
.A2(n_808),
.B(n_809),
.C(n_807),
.Y(n_8974)
);

O2A1O1Ixp5_ASAP7_75t_L g8975 ( 
.A1(n_8199),
.A2(n_8201),
.B(n_8240),
.C(n_8238),
.Y(n_8975)
);

INVx4_ASAP7_75t_L g8976 ( 
.A(n_8241),
.Y(n_8976)
);

INVx1_ASAP7_75t_L g8977 ( 
.A(n_7991),
.Y(n_8977)
);

INVxp67_ASAP7_75t_L g8978 ( 
.A(n_8117),
.Y(n_8978)
);

O2A1O1Ixp33_ASAP7_75t_L g8979 ( 
.A1(n_7990),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_8979)
);

O2A1O1Ixp5_ASAP7_75t_L g8980 ( 
.A1(n_7954),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_8980)
);

AND2x4_ASAP7_75t_L g8981 ( 
.A(n_7948),
.B(n_808),
.Y(n_8981)
);

INVx2_ASAP7_75t_L g8982 ( 
.A(n_7930),
.Y(n_8982)
);

BUFx12f_ASAP7_75t_L g8983 ( 
.A(n_8289),
.Y(n_8983)
);

AOI21xp5_ASAP7_75t_L g8984 ( 
.A1(n_7940),
.A2(n_810),
.B(n_809),
.Y(n_8984)
);

BUFx6f_ASAP7_75t_L g8985 ( 
.A(n_7928),
.Y(n_8985)
);

A2O1A1Ixp33_ASAP7_75t_SL g8986 ( 
.A1(n_7927),
.A2(n_338),
.B(n_335),
.C(n_337),
.Y(n_8986)
);

HB1xp67_ASAP7_75t_L g8987 ( 
.A(n_8117),
.Y(n_8987)
);

OAI21x1_ASAP7_75t_L g8988 ( 
.A1(n_7942),
.A2(n_337),
.B(n_339),
.Y(n_8988)
);

CKINVDCx5p33_ASAP7_75t_R g8989 ( 
.A(n_7934),
.Y(n_8989)
);

AND2x2_ASAP7_75t_L g8990 ( 
.A(n_8186),
.B(n_810),
.Y(n_8990)
);

NAND2xp5_ASAP7_75t_L g8991 ( 
.A(n_7926),
.B(n_811),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_7991),
.Y(n_8992)
);

O2A1O1Ixp33_ASAP7_75t_L g8993 ( 
.A1(n_7990),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_8993)
);

INVxp67_ASAP7_75t_L g8994 ( 
.A(n_8117),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_7991),
.Y(n_8995)
);

HB1xp67_ASAP7_75t_L g8996 ( 
.A(n_8117),
.Y(n_8996)
);

OAI22xp5_ASAP7_75t_L g8997 ( 
.A1(n_7990),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_8997)
);

NAND2xp5_ASAP7_75t_L g8998 ( 
.A(n_7926),
.B(n_811),
.Y(n_8998)
);

INVx2_ASAP7_75t_L g8999 ( 
.A(n_7930),
.Y(n_8999)
);

NAND2xp5_ASAP7_75t_SL g9000 ( 
.A(n_7940),
.B(n_812),
.Y(n_9000)
);

INVx2_ASAP7_75t_L g9001 ( 
.A(n_7930),
.Y(n_9001)
);

NOR2xp33_ASAP7_75t_L g9002 ( 
.A(n_7926),
.B(n_812),
.Y(n_9002)
);

O2A1O1Ixp33_ASAP7_75t_L g9003 ( 
.A1(n_7990),
.A2(n_343),
.B(n_340),
.C(n_342),
.Y(n_9003)
);

INVx1_ASAP7_75t_L g9004 ( 
.A(n_7991),
.Y(n_9004)
);

INVx4_ASAP7_75t_L g9005 ( 
.A(n_7928),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_7991),
.Y(n_9006)
);

NOR2xp33_ASAP7_75t_L g9007 ( 
.A(n_7926),
.B(n_813),
.Y(n_9007)
);

NAND2xp5_ASAP7_75t_L g9008 ( 
.A(n_7926),
.B(n_813),
.Y(n_9008)
);

AOI21xp5_ASAP7_75t_L g9009 ( 
.A1(n_7940),
.A2(n_815),
.B(n_814),
.Y(n_9009)
);

INVx3_ASAP7_75t_L g9010 ( 
.A(n_8123),
.Y(n_9010)
);

INVx2_ASAP7_75t_SL g9011 ( 
.A(n_7928),
.Y(n_9011)
);

NAND2xp5_ASAP7_75t_L g9012 ( 
.A(n_7926),
.B(n_814),
.Y(n_9012)
);

NOR2xp33_ASAP7_75t_R g9013 ( 
.A(n_7934),
.B(n_343),
.Y(n_9013)
);

BUFx6f_ASAP7_75t_L g9014 ( 
.A(n_7928),
.Y(n_9014)
);

CKINVDCx5p33_ASAP7_75t_R g9015 ( 
.A(n_7934),
.Y(n_9015)
);

OAI21xp5_ASAP7_75t_L g9016 ( 
.A1(n_7990),
.A2(n_343),
.B(n_344),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_7991),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_7991),
.Y(n_9018)
);

AOI21xp5_ASAP7_75t_L g9019 ( 
.A1(n_7940),
.A2(n_816),
.B(n_815),
.Y(n_9019)
);

AND2x2_ASAP7_75t_L g9020 ( 
.A(n_8186),
.B(n_816),
.Y(n_9020)
);

HB1xp67_ASAP7_75t_L g9021 ( 
.A(n_8117),
.Y(n_9021)
);

HB1xp67_ASAP7_75t_L g9022 ( 
.A(n_8117),
.Y(n_9022)
);

NOR2xp33_ASAP7_75t_L g9023 ( 
.A(n_7926),
.B(n_817),
.Y(n_9023)
);

AOI21xp5_ASAP7_75t_L g9024 ( 
.A1(n_7940),
.A2(n_818),
.B(n_817),
.Y(n_9024)
);

NOR3xp33_ASAP7_75t_SL g9025 ( 
.A(n_7990),
.B(n_344),
.C(n_345),
.Y(n_9025)
);

AOI21xp5_ASAP7_75t_L g9026 ( 
.A1(n_7940),
.A2(n_819),
.B(n_818),
.Y(n_9026)
);

AOI21xp5_ASAP7_75t_L g9027 ( 
.A1(n_7940),
.A2(n_821),
.B(n_820),
.Y(n_9027)
);

BUFx6f_ASAP7_75t_L g9028 ( 
.A(n_8693),
.Y(n_9028)
);

OAI22xp5_ASAP7_75t_L g9029 ( 
.A1(n_8474),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_9029)
);

BUFx3_ASAP7_75t_L g9030 ( 
.A(n_8649),
.Y(n_9030)
);

BUFx12f_ASAP7_75t_L g9031 ( 
.A(n_8522),
.Y(n_9031)
);

NAND2x1p5_ASAP7_75t_L g9032 ( 
.A(n_8810),
.B(n_820),
.Y(n_9032)
);

AOI222xp33_ASAP7_75t_L g9033 ( 
.A1(n_8580),
.A2(n_348),
.B1(n_350),
.B2(n_346),
.C1(n_347),
.C2(n_349),
.Y(n_9033)
);

OAI22xp5_ASAP7_75t_L g9034 ( 
.A1(n_9025),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_9034)
);

BUFx6f_ASAP7_75t_L g9035 ( 
.A(n_8693),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_8481),
.Y(n_9036)
);

OR2x2_ASAP7_75t_L g9037 ( 
.A(n_8925),
.B(n_821),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_8490),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8494),
.Y(n_9039)
);

NAND2xp33_ASAP7_75t_L g9040 ( 
.A(n_8518),
.B(n_347),
.Y(n_9040)
);

NOR2xp33_ASAP7_75t_L g9041 ( 
.A(n_8517),
.B(n_822),
.Y(n_9041)
);

BUFx3_ASAP7_75t_L g9042 ( 
.A(n_8649),
.Y(n_9042)
);

NAND2xp5_ASAP7_75t_L g9043 ( 
.A(n_8485),
.B(n_823),
.Y(n_9043)
);

AND2x6_ASAP7_75t_L g9044 ( 
.A(n_8500),
.B(n_823),
.Y(n_9044)
);

INVx3_ASAP7_75t_L g9045 ( 
.A(n_8606),
.Y(n_9045)
);

INVx2_ASAP7_75t_L g9046 ( 
.A(n_8664),
.Y(n_9046)
);

BUFx6f_ASAP7_75t_L g9047 ( 
.A(n_8661),
.Y(n_9047)
);

A2O1A1Ixp33_ASAP7_75t_L g9048 ( 
.A1(n_8471),
.A2(n_825),
.B(n_826),
.C(n_824),
.Y(n_9048)
);

NOR3xp33_ASAP7_75t_L g9049 ( 
.A(n_9016),
.B(n_349),
.C(n_350),
.Y(n_9049)
);

INVxp67_ASAP7_75t_SL g9050 ( 
.A(n_8534),
.Y(n_9050)
);

INVx1_ASAP7_75t_SL g9051 ( 
.A(n_8773),
.Y(n_9051)
);

HB1xp67_ASAP7_75t_L g9052 ( 
.A(n_8480),
.Y(n_9052)
);

BUFx3_ASAP7_75t_L g9053 ( 
.A(n_8661),
.Y(n_9053)
);

CKINVDCx20_ASAP7_75t_R g9054 ( 
.A(n_8493),
.Y(n_9054)
);

INVx1_ASAP7_75t_L g9055 ( 
.A(n_8499),
.Y(n_9055)
);

OAI22xp5_ASAP7_75t_L g9056 ( 
.A1(n_8624),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_9056)
);

BUFx4f_ASAP7_75t_SL g9057 ( 
.A(n_8653),
.Y(n_9057)
);

BUFx3_ASAP7_75t_L g9058 ( 
.A(n_8639),
.Y(n_9058)
);

NOR2xp33_ASAP7_75t_L g9059 ( 
.A(n_8861),
.B(n_825),
.Y(n_9059)
);

INVx2_ASAP7_75t_L g9060 ( 
.A(n_8680),
.Y(n_9060)
);

NAND2xp5_ASAP7_75t_L g9061 ( 
.A(n_8987),
.B(n_826),
.Y(n_9061)
);

O2A1O1Ixp33_ASAP7_75t_SL g9062 ( 
.A1(n_8864),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_L g9063 ( 
.A(n_8996),
.B(n_827),
.Y(n_9063)
);

AOI22xp33_ASAP7_75t_L g9064 ( 
.A1(n_8531),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_9064)
);

INVx3_ASAP7_75t_L g9065 ( 
.A(n_8606),
.Y(n_9065)
);

INVx1_ASAP7_75t_L g9066 ( 
.A(n_8505),
.Y(n_9066)
);

OR2x2_ASAP7_75t_L g9067 ( 
.A(n_8928),
.B(n_828),
.Y(n_9067)
);

INVxp67_ASAP7_75t_SL g9068 ( 
.A(n_8712),
.Y(n_9068)
);

OR2x2_ASAP7_75t_L g9069 ( 
.A(n_8927),
.B(n_828),
.Y(n_9069)
);

AND2x2_ASAP7_75t_L g9070 ( 
.A(n_8619),
.B(n_829),
.Y(n_9070)
);

NOR2xp33_ASAP7_75t_L g9071 ( 
.A(n_8571),
.B(n_830),
.Y(n_9071)
);

BUFx6f_ASAP7_75t_L g9072 ( 
.A(n_8479),
.Y(n_9072)
);

CKINVDCx11_ASAP7_75t_R g9073 ( 
.A(n_8983),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8507),
.Y(n_9074)
);

OAI22xp5_ASAP7_75t_L g9075 ( 
.A1(n_8656),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8520),
.Y(n_9076)
);

INVx2_ASAP7_75t_SL g9077 ( 
.A(n_8639),
.Y(n_9077)
);

INVx1_ASAP7_75t_L g9078 ( 
.A(n_8524),
.Y(n_9078)
);

OR2x2_ASAP7_75t_L g9079 ( 
.A(n_8910),
.B(n_830),
.Y(n_9079)
);

BUFx6f_ASAP7_75t_L g9080 ( 
.A(n_8479),
.Y(n_9080)
);

OR2x2_ASAP7_75t_L g9081 ( 
.A(n_8932),
.B(n_831),
.Y(n_9081)
);

INVx2_ASAP7_75t_L g9082 ( 
.A(n_8745),
.Y(n_9082)
);

HB1xp67_ASAP7_75t_L g9083 ( 
.A(n_9021),
.Y(n_9083)
);

INVx2_ASAP7_75t_L g9084 ( 
.A(n_8688),
.Y(n_9084)
);

INVx3_ASAP7_75t_L g9085 ( 
.A(n_8488),
.Y(n_9085)
);

AND2x4_ASAP7_75t_L g9086 ( 
.A(n_8978),
.B(n_831),
.Y(n_9086)
);

INVx2_ASAP7_75t_SL g9087 ( 
.A(n_8488),
.Y(n_9087)
);

BUFx3_ASAP7_75t_L g9088 ( 
.A(n_8589),
.Y(n_9088)
);

NAND2xp5_ASAP7_75t_L g9089 ( 
.A(n_9022),
.B(n_832),
.Y(n_9089)
);

NAND2xp5_ASAP7_75t_L g9090 ( 
.A(n_8732),
.B(n_832),
.Y(n_9090)
);

NAND2xp5_ASAP7_75t_SL g9091 ( 
.A(n_8810),
.B(n_833),
.Y(n_9091)
);

INVx3_ASAP7_75t_L g9092 ( 
.A(n_8551),
.Y(n_9092)
);

INVx2_ASAP7_75t_SL g9093 ( 
.A(n_8551),
.Y(n_9093)
);

INVx2_ASAP7_75t_SL g9094 ( 
.A(n_8578),
.Y(n_9094)
);

INVx4_ASAP7_75t_L g9095 ( 
.A(n_8823),
.Y(n_9095)
);

AOI22xp33_ASAP7_75t_L g9096 ( 
.A1(n_8629),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_9096)
);

BUFx8_ASAP7_75t_L g9097 ( 
.A(n_8707),
.Y(n_9097)
);

NOR2xp33_ASAP7_75t_L g9098 ( 
.A(n_8875),
.B(n_833),
.Y(n_9098)
);

NAND2xp5_ASAP7_75t_L g9099 ( 
.A(n_8743),
.B(n_834),
.Y(n_9099)
);

HB1xp67_ASAP7_75t_L g9100 ( 
.A(n_8755),
.Y(n_9100)
);

AND2x2_ASAP7_75t_SL g9101 ( 
.A(n_8626),
.B(n_354),
.Y(n_9101)
);

INVx1_ASAP7_75t_L g9102 ( 
.A(n_8526),
.Y(n_9102)
);

BUFx6f_ASAP7_75t_L g9103 ( 
.A(n_8578),
.Y(n_9103)
);

AO22x1_ASAP7_75t_L g9104 ( 
.A1(n_8810),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_9104)
);

AND2x4_ASAP7_75t_L g9105 ( 
.A(n_8994),
.B(n_8609),
.Y(n_9105)
);

INVx1_ASAP7_75t_L g9106 ( 
.A(n_8536),
.Y(n_9106)
);

NAND2x1p5_ASAP7_75t_L g9107 ( 
.A(n_8869),
.B(n_834),
.Y(n_9107)
);

BUFx2_ASAP7_75t_L g9108 ( 
.A(n_8563),
.Y(n_9108)
);

CKINVDCx20_ASAP7_75t_R g9109 ( 
.A(n_8989),
.Y(n_9109)
);

INVx5_ASAP7_75t_L g9110 ( 
.A(n_8696),
.Y(n_9110)
);

INVx4_ASAP7_75t_L g9111 ( 
.A(n_8832),
.Y(n_9111)
);

INVx2_ASAP7_75t_L g9112 ( 
.A(n_8691),
.Y(n_9112)
);

NAND2x1p5_ASAP7_75t_L g9113 ( 
.A(n_8869),
.B(n_835),
.Y(n_9113)
);

INVx2_ASAP7_75t_L g9114 ( 
.A(n_8720),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_8538),
.Y(n_9115)
);

NOR2xp33_ASAP7_75t_L g9116 ( 
.A(n_8937),
.B(n_835),
.Y(n_9116)
);

INVx2_ASAP7_75t_SL g9117 ( 
.A(n_8985),
.Y(n_9117)
);

OAI22xp5_ASAP7_75t_L g9118 ( 
.A1(n_8621),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_9118)
);

NAND2xp5_ASAP7_75t_L g9119 ( 
.A(n_8831),
.B(n_836),
.Y(n_9119)
);

INVx2_ASAP7_75t_L g9120 ( 
.A(n_8703),
.Y(n_9120)
);

NAND2xp5_ASAP7_75t_L g9121 ( 
.A(n_8748),
.B(n_837),
.Y(n_9121)
);

NOR2x1_ASAP7_75t_SL g9122 ( 
.A(n_8869),
.B(n_837),
.Y(n_9122)
);

HB1xp67_ASAP7_75t_L g9123 ( 
.A(n_8756),
.Y(n_9123)
);

A2O1A1Ixp33_ASAP7_75t_L g9124 ( 
.A1(n_8573),
.A2(n_839),
.B(n_840),
.C(n_838),
.Y(n_9124)
);

INVx4_ASAP7_75t_L g9125 ( 
.A(n_8985),
.Y(n_9125)
);

INVx2_ASAP7_75t_L g9126 ( 
.A(n_8541),
.Y(n_9126)
);

NOR2x1_ASAP7_75t_L g9127 ( 
.A(n_8473),
.B(n_838),
.Y(n_9127)
);

AND2x2_ASAP7_75t_L g9128 ( 
.A(n_8918),
.B(n_839),
.Y(n_9128)
);

NOR2xp33_ASAP7_75t_SL g9129 ( 
.A(n_8803),
.B(n_357),
.Y(n_9129)
);

NAND3xp33_ASAP7_75t_L g9130 ( 
.A(n_8616),
.B(n_358),
.C(n_359),
.Y(n_9130)
);

INVx1_ASAP7_75t_L g9131 ( 
.A(n_8567),
.Y(n_9131)
);

INVx1_ASAP7_75t_L g9132 ( 
.A(n_8574),
.Y(n_9132)
);

INVx2_ASAP7_75t_L g9133 ( 
.A(n_8586),
.Y(n_9133)
);

INVx5_ASAP7_75t_L g9134 ( 
.A(n_8807),
.Y(n_9134)
);

AOI22xp33_ASAP7_75t_L g9135 ( 
.A1(n_8508),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_9135)
);

INVx2_ASAP7_75t_L g9136 ( 
.A(n_8599),
.Y(n_9136)
);

BUFx6f_ASAP7_75t_L g9137 ( 
.A(n_9014),
.Y(n_9137)
);

INVx3_ASAP7_75t_L g9138 ( 
.A(n_9014),
.Y(n_9138)
);

BUFx3_ASAP7_75t_L g9139 ( 
.A(n_8568),
.Y(n_9139)
);

BUFx3_ASAP7_75t_L g9140 ( 
.A(n_8759),
.Y(n_9140)
);

AO32x1_ASAP7_75t_L g9141 ( 
.A1(n_8770),
.A2(n_362),
.A3(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_9141)
);

HB1xp67_ASAP7_75t_L g9142 ( 
.A(n_8794),
.Y(n_9142)
);

INVx2_ASAP7_75t_L g9143 ( 
.A(n_8622),
.Y(n_9143)
);

BUFx6f_ASAP7_75t_L g9144 ( 
.A(n_8730),
.Y(n_9144)
);

NOR2xp33_ASAP7_75t_L g9145 ( 
.A(n_8711),
.B(n_8893),
.Y(n_9145)
);

BUFx2_ASAP7_75t_L g9146 ( 
.A(n_8613),
.Y(n_9146)
);

AOI21xp5_ASAP7_75t_L g9147 ( 
.A1(n_8549),
.A2(n_361),
.B(n_362),
.Y(n_9147)
);

A2O1A1Ixp33_ASAP7_75t_L g9148 ( 
.A1(n_8628),
.A2(n_841),
.B(n_842),
.C(n_840),
.Y(n_9148)
);

OR2x6_ASAP7_75t_L g9149 ( 
.A(n_8733),
.B(n_841),
.Y(n_9149)
);

NAND2xp5_ASAP7_75t_L g9150 ( 
.A(n_8849),
.B(n_842),
.Y(n_9150)
);

BUFx2_ASAP7_75t_L g9151 ( 
.A(n_8805),
.Y(n_9151)
);

AOI22xp33_ASAP7_75t_SL g9152 ( 
.A1(n_8620),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_9152)
);

INVx1_ASAP7_75t_L g9153 ( 
.A(n_8636),
.Y(n_9153)
);

AND2x2_ASAP7_75t_L g9154 ( 
.A(n_8919),
.B(n_843),
.Y(n_9154)
);

BUFx6f_ASAP7_75t_L g9155 ( 
.A(n_8730),
.Y(n_9155)
);

INVx2_ASAP7_75t_SL g9156 ( 
.A(n_8557),
.Y(n_9156)
);

INVx3_ASAP7_75t_L g9157 ( 
.A(n_8516),
.Y(n_9157)
);

INVx2_ASAP7_75t_L g9158 ( 
.A(n_8648),
.Y(n_9158)
);

AND2x2_ASAP7_75t_SL g9159 ( 
.A(n_8941),
.B(n_363),
.Y(n_9159)
);

OAI22xp5_ASAP7_75t_L g9160 ( 
.A1(n_8638),
.A2(n_367),
.B1(n_364),
.B2(n_366),
.Y(n_9160)
);

CKINVDCx20_ASAP7_75t_R g9161 ( 
.A(n_9015),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8654),
.Y(n_9162)
);

OAI21xp33_ASAP7_75t_L g9163 ( 
.A1(n_8509),
.A2(n_364),
.B(n_366),
.Y(n_9163)
);

BUFx3_ASAP7_75t_L g9164 ( 
.A(n_8789),
.Y(n_9164)
);

INVx2_ASAP7_75t_L g9165 ( 
.A(n_8689),
.Y(n_9165)
);

CKINVDCx6p67_ASAP7_75t_R g9166 ( 
.A(n_8726),
.Y(n_9166)
);

BUFx2_ASAP7_75t_L g9167 ( 
.A(n_8566),
.Y(n_9167)
);

INVx4_ASAP7_75t_L g9168 ( 
.A(n_8768),
.Y(n_9168)
);

NAND2xp5_ASAP7_75t_L g9169 ( 
.A(n_8855),
.B(n_844),
.Y(n_9169)
);

INVx1_ASAP7_75t_L g9170 ( 
.A(n_8698),
.Y(n_9170)
);

BUFx3_ASAP7_75t_L g9171 ( 
.A(n_8771),
.Y(n_9171)
);

BUFx3_ASAP7_75t_L g9172 ( 
.A(n_8811),
.Y(n_9172)
);

NAND2xp5_ASAP7_75t_L g9173 ( 
.A(n_8858),
.B(n_844),
.Y(n_9173)
);

OAI21xp33_ASAP7_75t_L g9174 ( 
.A1(n_8973),
.A2(n_366),
.B(n_367),
.Y(n_9174)
);

AOI22xp33_ASAP7_75t_L g9175 ( 
.A1(n_8496),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_9175)
);

AOI22xp5_ASAP7_75t_L g9176 ( 
.A1(n_8477),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_9176)
);

INVx1_ASAP7_75t_L g9177 ( 
.A(n_8700),
.Y(n_9177)
);

INVx5_ASAP7_75t_L g9178 ( 
.A(n_8795),
.Y(n_9178)
);

INVx1_ASAP7_75t_L g9179 ( 
.A(n_8977),
.Y(n_9179)
);

HB1xp67_ASAP7_75t_L g9180 ( 
.A(n_8728),
.Y(n_9180)
);

AOI22xp33_ASAP7_75t_SL g9181 ( 
.A1(n_8663),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_9181)
);

BUFx12f_ASAP7_75t_L g9182 ( 
.A(n_8795),
.Y(n_9182)
);

INVx3_ASAP7_75t_L g9183 ( 
.A(n_8572),
.Y(n_9183)
);

INVx1_ASAP7_75t_L g9184 ( 
.A(n_8992),
.Y(n_9184)
);

CKINVDCx5p33_ASAP7_75t_R g9185 ( 
.A(n_8658),
.Y(n_9185)
);

INVx2_ASAP7_75t_SL g9186 ( 
.A(n_8816),
.Y(n_9186)
);

AOI22xp33_ASAP7_75t_L g9187 ( 
.A1(n_8595),
.A2(n_8637),
.B1(n_8603),
.B2(n_8677),
.Y(n_9187)
);

AOI22xp33_ASAP7_75t_L g9188 ( 
.A1(n_8590),
.A2(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_9188)
);

HB1xp67_ASAP7_75t_L g9189 ( 
.A(n_8740),
.Y(n_9189)
);

AND3x2_ASAP7_75t_L g9190 ( 
.A(n_8540),
.B(n_372),
.C(n_373),
.Y(n_9190)
);

INVx1_ASAP7_75t_L g9191 ( 
.A(n_8995),
.Y(n_9191)
);

OAI21xp5_ASAP7_75t_L g9192 ( 
.A1(n_8824),
.A2(n_372),
.B(n_373),
.Y(n_9192)
);

INVxp67_ASAP7_75t_SL g9193 ( 
.A(n_8800),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_9004),
.Y(n_9194)
);

AOI22xp5_ASAP7_75t_L g9195 ( 
.A1(n_8585),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_9195)
);

AOI21xp5_ASAP7_75t_L g9196 ( 
.A1(n_8587),
.A2(n_374),
.B(n_375),
.Y(n_9196)
);

INVxp67_ASAP7_75t_L g9197 ( 
.A(n_8697),
.Y(n_9197)
);

INVx1_ASAP7_75t_SL g9198 ( 
.A(n_8822),
.Y(n_9198)
);

INVx2_ASAP7_75t_L g9199 ( 
.A(n_9006),
.Y(n_9199)
);

INVx1_ASAP7_75t_SL g9200 ( 
.A(n_8836),
.Y(n_9200)
);

BUFx6f_ASAP7_75t_SL g9201 ( 
.A(n_8655),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_9017),
.Y(n_9202)
);

HB1xp67_ASAP7_75t_L g9203 ( 
.A(n_8934),
.Y(n_9203)
);

BUFx6f_ASAP7_75t_L g9204 ( 
.A(n_9011),
.Y(n_9204)
);

AOI22xp33_ASAP7_75t_L g9205 ( 
.A1(n_8647),
.A2(n_8594),
.B1(n_8705),
.B2(n_8652),
.Y(n_9205)
);

NAND2xp5_ASAP7_75t_L g9206 ( 
.A(n_8881),
.B(n_845),
.Y(n_9206)
);

BUFx2_ASAP7_75t_R g9207 ( 
.A(n_8887),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_9018),
.Y(n_9208)
);

BUFx12f_ASAP7_75t_L g9209 ( 
.A(n_8655),
.Y(n_9209)
);

AND2x4_ASAP7_75t_L g9210 ( 
.A(n_8754),
.B(n_845),
.Y(n_9210)
);

NAND2xp5_ASAP7_75t_L g9211 ( 
.A(n_8884),
.B(n_846),
.Y(n_9211)
);

BUFx12f_ASAP7_75t_L g9212 ( 
.A(n_8716),
.Y(n_9212)
);

CKINVDCx20_ASAP7_75t_R g9213 ( 
.A(n_8848),
.Y(n_9213)
);

INVx3_ASAP7_75t_L g9214 ( 
.A(n_9005),
.Y(n_9214)
);

BUFx6f_ASAP7_75t_L g9215 ( 
.A(n_8891),
.Y(n_9215)
);

BUFx2_ASAP7_75t_L g9216 ( 
.A(n_8758),
.Y(n_9216)
);

AOI222xp33_ASAP7_75t_L g9217 ( 
.A1(n_8731),
.A2(n_376),
.B1(n_378),
.B2(n_374),
.C1(n_375),
.C2(n_377),
.Y(n_9217)
);

AOI22xp5_ASAP7_75t_L g9218 ( 
.A1(n_8874),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_9218)
);

BUFx3_ASAP7_75t_L g9219 ( 
.A(n_8513),
.Y(n_9219)
);

CKINVDCx20_ASAP7_75t_R g9220 ( 
.A(n_8879),
.Y(n_9220)
);

INVx1_ASAP7_75t_L g9221 ( 
.A(n_8719),
.Y(n_9221)
);

BUFx3_ASAP7_75t_L g9222 ( 
.A(n_9010),
.Y(n_9222)
);

INVx3_ASAP7_75t_L g9223 ( 
.A(n_8704),
.Y(n_9223)
);

BUFx3_ASAP7_75t_L g9224 ( 
.A(n_8762),
.Y(n_9224)
);

OAI22xp5_ASAP7_75t_L g9225 ( 
.A1(n_8544),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_9225)
);

INVx1_ASAP7_75t_L g9226 ( 
.A(n_8809),
.Y(n_9226)
);

INVx1_ASAP7_75t_L g9227 ( 
.A(n_8657),
.Y(n_9227)
);

BUFx6f_ASAP7_75t_L g9228 ( 
.A(n_8777),
.Y(n_9228)
);

NAND2x2_ASAP7_75t_L g9229 ( 
.A(n_8949),
.B(n_8623),
.Y(n_9229)
);

AND2x4_ASAP7_75t_L g9230 ( 
.A(n_8894),
.B(n_846),
.Y(n_9230)
);

AOI22xp5_ASAP7_75t_L g9231 ( 
.A1(n_8723),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_9231)
);

INVx1_ASAP7_75t_SL g9232 ( 
.A(n_8898),
.Y(n_9232)
);

INVx4_ASAP7_75t_L g9233 ( 
.A(n_8877),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8833),
.Y(n_9234)
);

BUFx2_ASAP7_75t_L g9235 ( 
.A(n_8929),
.Y(n_9235)
);

CKINVDCx6p67_ASAP7_75t_R g9236 ( 
.A(n_8837),
.Y(n_9236)
);

AND2x4_ASAP7_75t_L g9237 ( 
.A(n_8906),
.B(n_847),
.Y(n_9237)
);

BUFx6f_ASAP7_75t_L g9238 ( 
.A(n_8632),
.Y(n_9238)
);

INVx2_ASAP7_75t_L g9239 ( 
.A(n_8472),
.Y(n_9239)
);

INVx3_ASAP7_75t_L g9240 ( 
.A(n_8497),
.Y(n_9240)
);

INVx1_ASAP7_75t_L g9241 ( 
.A(n_8751),
.Y(n_9241)
);

NAND2xp5_ASAP7_75t_SL g9242 ( 
.A(n_8671),
.B(n_848),
.Y(n_9242)
);

INVx4_ASAP7_75t_L g9243 ( 
.A(n_8582),
.Y(n_9243)
);

INVx6_ASAP7_75t_L g9244 ( 
.A(n_8873),
.Y(n_9244)
);

INVx4_ASAP7_75t_L g9245 ( 
.A(n_8617),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_8482),
.Y(n_9246)
);

INVx2_ASAP7_75t_SL g9247 ( 
.A(n_8532),
.Y(n_9247)
);

BUFx4f_ASAP7_75t_L g9248 ( 
.A(n_8716),
.Y(n_9248)
);

NOR3xp33_ASAP7_75t_L g9249 ( 
.A(n_8690),
.B(n_379),
.C(n_380),
.Y(n_9249)
);

AOI22xp33_ASAP7_75t_L g9250 ( 
.A1(n_8615),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_8487),
.Y(n_9251)
);

INVx1_ASAP7_75t_SL g9252 ( 
.A(n_8909),
.Y(n_9252)
);

AOI22xp33_ASAP7_75t_L g9253 ( 
.A1(n_8476),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_9253)
);

AOI22xp33_ASAP7_75t_L g9254 ( 
.A1(n_8752),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_9254)
);

AOI21xp5_ASAP7_75t_L g9255 ( 
.A1(n_8896),
.A2(n_383),
.B(n_384),
.Y(n_9255)
);

NAND2xp5_ASAP7_75t_L g9256 ( 
.A(n_8814),
.B(n_848),
.Y(n_9256)
);

BUFx2_ASAP7_75t_L g9257 ( 
.A(n_8929),
.Y(n_9257)
);

AOI21xp5_ASAP7_75t_L g9258 ( 
.A1(n_8886),
.A2(n_384),
.B(n_385),
.Y(n_9258)
);

NOR2xp67_ASAP7_75t_L g9259 ( 
.A(n_8781),
.B(n_385),
.Y(n_9259)
);

BUFx4f_ASAP7_75t_L g9260 ( 
.A(n_8676),
.Y(n_9260)
);

AND2x6_ASAP7_75t_L g9261 ( 
.A(n_8971),
.B(n_8959),
.Y(n_9261)
);

BUFx3_ASAP7_75t_L g9262 ( 
.A(n_8642),
.Y(n_9262)
);

INVx4_ASAP7_75t_L g9263 ( 
.A(n_8521),
.Y(n_9263)
);

BUFx2_ASAP7_75t_L g9264 ( 
.A(n_8845),
.Y(n_9264)
);

BUFx2_ASAP7_75t_L g9265 ( 
.A(n_8907),
.Y(n_9265)
);

INVx4_ASAP7_75t_L g9266 ( 
.A(n_8981),
.Y(n_9266)
);

INVx2_ASAP7_75t_SL g9267 ( 
.A(n_8529),
.Y(n_9267)
);

A2O1A1Ixp33_ASAP7_75t_L g9268 ( 
.A1(n_8979),
.A2(n_851),
.B(n_852),
.C(n_849),
.Y(n_9268)
);

AOI22xp33_ASAP7_75t_L g9269 ( 
.A1(n_8746),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_8815),
.B(n_851),
.Y(n_9270)
);

INVx3_ASAP7_75t_SL g9271 ( 
.A(n_8844),
.Y(n_9271)
);

AND2x2_ASAP7_75t_L g9272 ( 
.A(n_8506),
.B(n_8483),
.Y(n_9272)
);

INVx1_ASAP7_75t_L g9273 ( 
.A(n_8501),
.Y(n_9273)
);

AOI22xp5_ASAP7_75t_L g9274 ( 
.A1(n_9002),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8510),
.Y(n_9275)
);

AND2x4_ASAP7_75t_L g9276 ( 
.A(n_8523),
.B(n_852),
.Y(n_9276)
);

AND2x2_ASAP7_75t_L g9277 ( 
.A(n_8788),
.B(n_853),
.Y(n_9277)
);

AND2x6_ASAP7_75t_L g9278 ( 
.A(n_8948),
.B(n_853),
.Y(n_9278)
);

OR2x6_ASAP7_75t_L g9279 ( 
.A(n_8868),
.B(n_854),
.Y(n_9279)
);

INVx1_ASAP7_75t_SL g9280 ( 
.A(n_8546),
.Y(n_9280)
);

BUFx2_ASAP7_75t_L g9281 ( 
.A(n_8542),
.Y(n_9281)
);

AND2x4_ASAP7_75t_L g9282 ( 
.A(n_8604),
.B(n_854),
.Y(n_9282)
);

BUFx3_ASAP7_75t_L g9283 ( 
.A(n_8687),
.Y(n_9283)
);

BUFx6f_ASAP7_75t_L g9284 ( 
.A(n_8634),
.Y(n_9284)
);

AOI22xp5_ASAP7_75t_L g9285 ( 
.A1(n_9007),
.A2(n_9023),
.B1(n_8605),
.B2(n_8668),
.Y(n_9285)
);

AOI21x1_ASAP7_75t_L g9286 ( 
.A1(n_9000),
.A2(n_386),
.B(n_387),
.Y(n_9286)
);

OR2x6_ASAP7_75t_L g9287 ( 
.A(n_8820),
.B(n_855),
.Y(n_9287)
);

INVx3_ASAP7_75t_L g9288 ( 
.A(n_8635),
.Y(n_9288)
);

AND2x4_ASAP7_75t_L g9289 ( 
.A(n_8660),
.B(n_855),
.Y(n_9289)
);

BUFx2_ASAP7_75t_L g9290 ( 
.A(n_8982),
.Y(n_9290)
);

OAI22xp33_ASAP7_75t_L g9291 ( 
.A1(n_8812),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_9291)
);

CKINVDCx6p67_ASAP7_75t_R g9292 ( 
.A(n_8591),
.Y(n_9292)
);

OR2x2_ASAP7_75t_L g9293 ( 
.A(n_8778),
.B(n_858),
.Y(n_9293)
);

BUFx3_ASAP7_75t_L g9294 ( 
.A(n_8905),
.Y(n_9294)
);

INVx1_ASAP7_75t_L g9295 ( 
.A(n_8999),
.Y(n_9295)
);

AND2x4_ASAP7_75t_L g9296 ( 
.A(n_9001),
.B(n_858),
.Y(n_9296)
);

BUFx3_ASAP7_75t_L g9297 ( 
.A(n_8535),
.Y(n_9297)
);

INVx2_ASAP7_75t_L g9298 ( 
.A(n_8684),
.Y(n_9298)
);

AND2x2_ASAP7_75t_L g9299 ( 
.A(n_8779),
.B(n_8786),
.Y(n_9299)
);

NAND2xp5_ASAP7_75t_L g9300 ( 
.A(n_8847),
.B(n_859),
.Y(n_9300)
);

BUFx2_ASAP7_75t_L g9301 ( 
.A(n_8859),
.Y(n_9301)
);

INVx1_ASAP7_75t_SL g9302 ( 
.A(n_8911),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_8685),
.Y(n_9303)
);

AOI22xp33_ASAP7_75t_SL g9304 ( 
.A1(n_8511),
.A2(n_8577),
.B1(n_8502),
.B2(n_8997),
.Y(n_9304)
);

INVx2_ASAP7_75t_L g9305 ( 
.A(n_8729),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_8738),
.Y(n_9306)
);

INVxp67_ASAP7_75t_SL g9307 ( 
.A(n_8776),
.Y(n_9307)
);

BUFx6f_ASAP7_75t_L g9308 ( 
.A(n_8819),
.Y(n_9308)
);

AOI21xp5_ASAP7_75t_L g9309 ( 
.A1(n_8784),
.A2(n_389),
.B(n_390),
.Y(n_9309)
);

INVx5_ASAP7_75t_L g9310 ( 
.A(n_8820),
.Y(n_9310)
);

OR2x6_ASAP7_75t_L g9311 ( 
.A(n_8744),
.B(n_859),
.Y(n_9311)
);

INVx1_ASAP7_75t_L g9312 ( 
.A(n_8897),
.Y(n_9312)
);

BUFx6f_ASAP7_75t_L g9313 ( 
.A(n_8643),
.Y(n_9313)
);

NAND2xp5_ASAP7_75t_L g9314 ( 
.A(n_8852),
.B(n_860),
.Y(n_9314)
);

O2A1O1Ixp33_ASAP7_75t_L g9315 ( 
.A1(n_8675),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_9315)
);

BUFx2_ASAP7_75t_L g9316 ( 
.A(n_8802),
.Y(n_9316)
);

INVx2_ASAP7_75t_SL g9317 ( 
.A(n_8673),
.Y(n_9317)
);

INVx1_ASAP7_75t_L g9318 ( 
.A(n_8659),
.Y(n_9318)
);

INVx3_ASAP7_75t_L g9319 ( 
.A(n_8926),
.Y(n_9319)
);

AND2x2_ASAP7_75t_SL g9320 ( 
.A(n_8939),
.B(n_391),
.Y(n_9320)
);

BUFx6f_ASAP7_75t_L g9321 ( 
.A(n_8724),
.Y(n_9321)
);

NAND2xp5_ASAP7_75t_L g9322 ( 
.A(n_8857),
.B(n_8792),
.Y(n_9322)
);

INVx4_ASAP7_75t_L g9323 ( 
.A(n_8930),
.Y(n_9323)
);

NOR2xp33_ASAP7_75t_SL g9324 ( 
.A(n_8627),
.B(n_392),
.Y(n_9324)
);

NOR2xp33_ASAP7_75t_L g9325 ( 
.A(n_8581),
.B(n_861),
.Y(n_9325)
);

INVx6_ASAP7_75t_L g9326 ( 
.A(n_8527),
.Y(n_9326)
);

NAND2xp5_ASAP7_75t_SL g9327 ( 
.A(n_8562),
.B(n_862),
.Y(n_9327)
);

NAND2xp5_ASAP7_75t_L g9328 ( 
.A(n_8798),
.B(n_862),
.Y(n_9328)
);

AOI22xp5_ASAP7_75t_L g9329 ( 
.A1(n_8646),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_9329)
);

AND2x2_ASAP7_75t_L g9330 ( 
.A(n_8625),
.B(n_863),
.Y(n_9330)
);

NOR2xp67_ASAP7_75t_L g9331 ( 
.A(n_8512),
.B(n_393),
.Y(n_9331)
);

INVx4_ASAP7_75t_L g9332 ( 
.A(n_8976),
.Y(n_9332)
);

INVx2_ASAP7_75t_SL g9333 ( 
.A(n_8757),
.Y(n_9333)
);

NAND2x1_ASAP7_75t_SL g9334 ( 
.A(n_8963),
.B(n_863),
.Y(n_9334)
);

INVx2_ASAP7_75t_L g9335 ( 
.A(n_8774),
.Y(n_9335)
);

BUFx2_ASAP7_75t_L g9336 ( 
.A(n_8961),
.Y(n_9336)
);

INVx3_ASAP7_75t_L g9337 ( 
.A(n_8842),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8674),
.Y(n_9338)
);

AND2x2_ASAP7_75t_L g9339 ( 
.A(n_8630),
.B(n_864),
.Y(n_9339)
);

AND2x2_ASAP7_75t_L g9340 ( 
.A(n_8640),
.B(n_865),
.Y(n_9340)
);

BUFx2_ASAP7_75t_L g9341 ( 
.A(n_8964),
.Y(n_9341)
);

AOI22xp33_ASAP7_75t_L g9342 ( 
.A1(n_8960),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_9342)
);

INVx3_ASAP7_75t_L g9343 ( 
.A(n_8950),
.Y(n_9343)
);

INVx1_ASAP7_75t_L g9344 ( 
.A(n_8686),
.Y(n_9344)
);

BUFx2_ASAP7_75t_SL g9345 ( 
.A(n_8491),
.Y(n_9345)
);

HB1xp67_ASAP7_75t_L g9346 ( 
.A(n_8965),
.Y(n_9346)
);

BUFx12f_ASAP7_75t_L g9347 ( 
.A(n_8880),
.Y(n_9347)
);

AOI33xp33_ASAP7_75t_L g9348 ( 
.A1(n_8901),
.A2(n_396),
.A3(n_398),
.B1(n_394),
.B2(n_395),
.B3(n_397),
.Y(n_9348)
);

INVxp67_ASAP7_75t_L g9349 ( 
.A(n_8569),
.Y(n_9349)
);

INVxp67_ASAP7_75t_SL g9350 ( 
.A(n_8954),
.Y(n_9350)
);

AND2x4_ASAP7_75t_L g9351 ( 
.A(n_8958),
.B(n_865),
.Y(n_9351)
);

AOI22xp33_ASAP7_75t_SL g9352 ( 
.A1(n_8651),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_9352)
);

INVx1_ASAP7_75t_L g9353 ( 
.A(n_8699),
.Y(n_9353)
);

INVx1_ASAP7_75t_L g9354 ( 
.A(n_8706),
.Y(n_9354)
);

NAND2xp5_ASAP7_75t_L g9355 ( 
.A(n_8470),
.B(n_867),
.Y(n_9355)
);

INVx2_ASAP7_75t_SL g9356 ( 
.A(n_8990),
.Y(n_9356)
);

INVx1_ASAP7_75t_SL g9357 ( 
.A(n_8753),
.Y(n_9357)
);

INVx3_ASAP7_75t_L g9358 ( 
.A(n_8734),
.Y(n_9358)
);

INVx2_ASAP7_75t_L g9359 ( 
.A(n_8988),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_8558),
.Y(n_9360)
);

NAND2xp5_ASAP7_75t_L g9361 ( 
.A(n_8991),
.B(n_867),
.Y(n_9361)
);

AOI22xp5_ASAP7_75t_L g9362 ( 
.A1(n_8714),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_9362)
);

O2A1O1Ixp33_ASAP7_75t_L g9363 ( 
.A1(n_8498),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_9363)
);

INVx1_ASAP7_75t_L g9364 ( 
.A(n_8679),
.Y(n_9364)
);

HB1xp67_ASAP7_75t_L g9365 ( 
.A(n_8972),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_8559),
.Y(n_9366)
);

BUFx6f_ASAP7_75t_L g9367 ( 
.A(n_8519),
.Y(n_9367)
);

BUFx3_ASAP7_75t_L g9368 ( 
.A(n_8561),
.Y(n_9368)
);

OAI22xp5_ASAP7_75t_L g9369 ( 
.A1(n_8564),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_9369)
);

INVx2_ASAP7_75t_L g9370 ( 
.A(n_8588),
.Y(n_9370)
);

AND2x4_ASAP7_75t_L g9371 ( 
.A(n_8749),
.B(n_868),
.Y(n_9371)
);

AND2x6_ASAP7_75t_L g9372 ( 
.A(n_8955),
.B(n_868),
.Y(n_9372)
);

INVx1_ASAP7_75t_L g9373 ( 
.A(n_8763),
.Y(n_9373)
);

BUFx3_ASAP7_75t_L g9374 ( 
.A(n_8545),
.Y(n_9374)
);

OAI22xp33_ASAP7_75t_L g9375 ( 
.A1(n_8860),
.A2(n_8611),
.B1(n_8956),
.B2(n_8854),
.Y(n_9375)
);

INVx2_ASAP7_75t_SL g9376 ( 
.A(n_9020),
.Y(n_9376)
);

INVx1_ASAP7_75t_SL g9377 ( 
.A(n_8888),
.Y(n_9377)
);

AOI21xp5_ASAP7_75t_L g9378 ( 
.A1(n_8975),
.A2(n_403),
.B(n_404),
.Y(n_9378)
);

AND2x2_ASAP7_75t_L g9379 ( 
.A(n_8683),
.B(n_869),
.Y(n_9379)
);

NAND2xp5_ASAP7_75t_SL g9380 ( 
.A(n_8736),
.B(n_870),
.Y(n_9380)
);

BUFx2_ASAP7_75t_L g9381 ( 
.A(n_8495),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8853),
.Y(n_9382)
);

A2O1A1Ixp33_ASAP7_75t_L g9383 ( 
.A1(n_8993),
.A2(n_871),
.B(n_872),
.C(n_870),
.Y(n_9383)
);

AND2x4_ASAP7_75t_L g9384 ( 
.A(n_8944),
.B(n_873),
.Y(n_9384)
);

BUFx2_ASAP7_75t_L g9385 ( 
.A(n_8998),
.Y(n_9385)
);

INVx8_ASAP7_75t_L g9386 ( 
.A(n_8892),
.Y(n_9386)
);

BUFx2_ASAP7_75t_L g9387 ( 
.A(n_9008),
.Y(n_9387)
);

BUFx2_ASAP7_75t_L g9388 ( 
.A(n_9012),
.Y(n_9388)
);

NAND2xp5_ASAP7_75t_L g9389 ( 
.A(n_8537),
.B(n_873),
.Y(n_9389)
);

INVx2_ASAP7_75t_L g9390 ( 
.A(n_8853),
.Y(n_9390)
);

INVx3_ASAP7_75t_L g9391 ( 
.A(n_8902),
.Y(n_9391)
);

INVx1_ASAP7_75t_L g9392 ( 
.A(n_8935),
.Y(n_9392)
);

BUFx2_ASAP7_75t_L g9393 ( 
.A(n_8612),
.Y(n_9393)
);

INVx3_ASAP7_75t_L g9394 ( 
.A(n_8593),
.Y(n_9394)
);

BUFx2_ASAP7_75t_L g9395 ( 
.A(n_8550),
.Y(n_9395)
);

CKINVDCx11_ASAP7_75t_R g9396 ( 
.A(n_8592),
.Y(n_9396)
);

OAI21x1_ASAP7_75t_SL g9397 ( 
.A1(n_8631),
.A2(n_403),
.B(n_404),
.Y(n_9397)
);

OAI22x1_ASAP7_75t_L g9398 ( 
.A1(n_8584),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_9398)
);

INVx2_ASAP7_75t_SL g9399 ( 
.A(n_8694),
.Y(n_9399)
);

INVx1_ASAP7_75t_L g9400 ( 
.A(n_8936),
.Y(n_9400)
);

INVx2_ASAP7_75t_SL g9401 ( 
.A(n_8871),
.Y(n_9401)
);

NAND2xp5_ASAP7_75t_L g9402 ( 
.A(n_8923),
.B(n_874),
.Y(n_9402)
);

AOI21xp33_ASAP7_75t_L g9403 ( 
.A1(n_9003),
.A2(n_405),
.B(n_406),
.Y(n_9403)
);

NOR2x1_ASAP7_75t_L g9404 ( 
.A(n_8920),
.B(n_875),
.Y(n_9404)
);

AND2x4_ASAP7_75t_L g9405 ( 
.A(n_8515),
.B(n_875),
.Y(n_9405)
);

OR2x2_ASAP7_75t_L g9406 ( 
.A(n_8760),
.B(n_876),
.Y(n_9406)
);

OR2x6_ASAP7_75t_L g9407 ( 
.A(n_8601),
.B(n_876),
.Y(n_9407)
);

AOI222xp33_ASAP7_75t_L g9408 ( 
.A1(n_8618),
.A2(n_407),
.B1(n_409),
.B2(n_405),
.C1(n_406),
.C2(n_408),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_8908),
.Y(n_9409)
);

AND2x4_ASAP7_75t_L g9410 ( 
.A(n_8943),
.B(n_877),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_8945),
.Y(n_9411)
);

INVx1_ASAP7_75t_L g9412 ( 
.A(n_8913),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8914),
.Y(n_9413)
);

CKINVDCx5p33_ASAP7_75t_R g9414 ( 
.A(n_9013),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8924),
.Y(n_9415)
);

BUFx3_ASAP7_75t_L g9416 ( 
.A(n_8560),
.Y(n_9416)
);

AND2x2_ASAP7_75t_L g9417 ( 
.A(n_8737),
.B(n_877),
.Y(n_9417)
);

OR2x2_ASAP7_75t_L g9418 ( 
.A(n_8701),
.B(n_878),
.Y(n_9418)
);

BUFx3_ASAP7_75t_L g9419 ( 
.A(n_8775),
.Y(n_9419)
);

INVx4_ASAP7_75t_L g9420 ( 
.A(n_8957),
.Y(n_9420)
);

INVx3_ASAP7_75t_L g9421 ( 
.A(n_8840),
.Y(n_9421)
);

INVx1_ASAP7_75t_SL g9422 ( 
.A(n_8555),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8917),
.Y(n_9423)
);

INVx2_ASAP7_75t_L g9424 ( 
.A(n_8782),
.Y(n_9424)
);

AOI22xp5_ASAP7_75t_L g9425 ( 
.A1(n_8797),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_9425)
);

NAND2xp5_ASAP7_75t_L g9426 ( 
.A(n_8899),
.B(n_879),
.Y(n_9426)
);

INVx2_ASAP7_75t_L g9427 ( 
.A(n_8912),
.Y(n_9427)
);

INVx2_ASAP7_75t_SL g9428 ( 
.A(n_8838),
.Y(n_9428)
);

AOI21xp5_ASAP7_75t_L g9429 ( 
.A1(n_8984),
.A2(n_9019),
.B(n_9009),
.Y(n_9429)
);

OAI22xp5_ASAP7_75t_L g9430 ( 
.A1(n_8670),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_9430)
);

CKINVDCx8_ASAP7_75t_R g9431 ( 
.A(n_8829),
.Y(n_9431)
);

OAI22xp5_ASAP7_75t_SL g9432 ( 
.A1(n_8727),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_9432)
);

OR2x6_ASAP7_75t_SL g9433 ( 
.A(n_8922),
.B(n_410),
.Y(n_9433)
);

BUFx6f_ASAP7_75t_L g9434 ( 
.A(n_8556),
.Y(n_9434)
);

BUFx2_ASAP7_75t_SL g9435 ( 
.A(n_8839),
.Y(n_9435)
);

NOR3xp33_ASAP7_75t_L g9436 ( 
.A(n_8682),
.B(n_411),
.C(n_412),
.Y(n_9436)
);

OAI22xp5_ASAP7_75t_L g9437 ( 
.A1(n_8717),
.A2(n_411),
.B1(n_412),
.B2(n_881),
.Y(n_9437)
);

AND2x2_ASAP7_75t_L g9438 ( 
.A(n_8915),
.B(n_882),
.Y(n_9438)
);

AOI22xp5_ASAP7_75t_L g9439 ( 
.A1(n_8846),
.A2(n_884),
.B1(n_882),
.B2(n_883),
.Y(n_9439)
);

OR2x2_ASAP7_75t_L g9440 ( 
.A(n_8841),
.B(n_883),
.Y(n_9440)
);

HB1xp67_ASAP7_75t_L g9441 ( 
.A(n_8947),
.Y(n_9441)
);

AND2x4_ASAP7_75t_L g9442 ( 
.A(n_8878),
.B(n_886),
.Y(n_9442)
);

INVx2_ASAP7_75t_L g9443 ( 
.A(n_8862),
.Y(n_9443)
);

AOI22xp33_ASAP7_75t_L g9444 ( 
.A1(n_8785),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.Y(n_9444)
);

INVx1_ASAP7_75t_L g9445 ( 
.A(n_8721),
.Y(n_9445)
);

NOR2xp33_ASAP7_75t_SL g9446 ( 
.A(n_8739),
.B(n_887),
.Y(n_9446)
);

AOI22xp33_ASAP7_75t_L g9447 ( 
.A1(n_8780),
.A2(n_890),
.B1(n_888),
.B2(n_889),
.Y(n_9447)
);

INVx3_ASAP7_75t_L g9448 ( 
.A(n_8575),
.Y(n_9448)
);

NAND3x1_ASAP7_75t_L g9449 ( 
.A(n_8806),
.B(n_8825),
.C(n_8850),
.Y(n_9449)
);

BUFx6f_ASAP7_75t_L g9450 ( 
.A(n_8596),
.Y(n_9450)
);

BUFx3_ASAP7_75t_L g9451 ( 
.A(n_8876),
.Y(n_9451)
);

AOI22xp33_ASAP7_75t_SL g9452 ( 
.A1(n_8765),
.A2(n_892),
.B1(n_889),
.B2(n_891),
.Y(n_9452)
);

OR2x2_ASAP7_75t_L g9453 ( 
.A(n_8890),
.B(n_891),
.Y(n_9453)
);

INVx6_ASAP7_75t_SL g9454 ( 
.A(n_8830),
.Y(n_9454)
);

INVx4_ASAP7_75t_L g9455 ( 
.A(n_8952),
.Y(n_9455)
);

BUFx12f_ASAP7_75t_L g9456 ( 
.A(n_8813),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_L g9457 ( 
.A(n_8863),
.B(n_893),
.Y(n_9457)
);

BUFx3_ASAP7_75t_L g9458 ( 
.A(n_8597),
.Y(n_9458)
);

NAND2x1p5_ASAP7_75t_L g9459 ( 
.A(n_8966),
.B(n_893),
.Y(n_9459)
);

BUFx3_ASAP7_75t_L g9460 ( 
.A(n_8598),
.Y(n_9460)
);

NAND2xp5_ASAP7_75t_L g9461 ( 
.A(n_8867),
.B(n_894),
.Y(n_9461)
);

AND2x2_ASAP7_75t_L g9462 ( 
.A(n_8796),
.B(n_894),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_8528),
.Y(n_9463)
);

AOI21xp33_ASAP7_75t_L g9464 ( 
.A1(n_8986),
.A2(n_895),
.B(n_896),
.Y(n_9464)
);

NOR2xp33_ASAP7_75t_L g9465 ( 
.A(n_8708),
.B(n_898),
.Y(n_9465)
);

AOI21xp5_ASAP7_75t_L g9466 ( 
.A1(n_9024),
.A2(n_898),
.B(n_899),
.Y(n_9466)
);

AOI22xp5_ASAP7_75t_L g9467 ( 
.A1(n_8772),
.A2(n_903),
.B1(n_901),
.B2(n_902),
.Y(n_9467)
);

INVx5_ASAP7_75t_L g9468 ( 
.A(n_8821),
.Y(n_9468)
);

CKINVDCx20_ASAP7_75t_R g9469 ( 
.A(n_8783),
.Y(n_9469)
);

NOR2xp67_ASAP7_75t_L g9470 ( 
.A(n_8484),
.B(n_902),
.Y(n_9470)
);

INVx1_ASAP7_75t_L g9471 ( 
.A(n_8644),
.Y(n_9471)
);

INVx2_ASAP7_75t_SL g9472 ( 
.A(n_8903),
.Y(n_9472)
);

INVx3_ASAP7_75t_L g9473 ( 
.A(n_8790),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_8722),
.Y(n_9474)
);

AOI21xp5_ASAP7_75t_L g9475 ( 
.A1(n_9026),
.A2(n_903),
.B(n_904),
.Y(n_9475)
);

NAND2xp5_ASAP7_75t_L g9476 ( 
.A(n_8791),
.B(n_904),
.Y(n_9476)
);

OAI22xp5_ASAP7_75t_L g9477 ( 
.A1(n_8543),
.A2(n_907),
.B1(n_905),
.B2(n_906),
.Y(n_9477)
);

INVx1_ASAP7_75t_L g9478 ( 
.A(n_8916),
.Y(n_9478)
);

AND2x4_ASAP7_75t_SL g9479 ( 
.A(n_8870),
.B(n_8672),
.Y(n_9479)
);

AND2x4_ASAP7_75t_L g9480 ( 
.A(n_8530),
.B(n_905),
.Y(n_9480)
);

AND2x4_ASAP7_75t_L g9481 ( 
.A(n_8968),
.B(n_906),
.Y(n_9481)
);

BUFx12f_ASAP7_75t_L g9482 ( 
.A(n_8769),
.Y(n_9482)
);

INVx1_ASAP7_75t_L g9483 ( 
.A(n_8650),
.Y(n_9483)
);

INVx4_ASAP7_75t_L g9484 ( 
.A(n_8662),
.Y(n_9484)
);

HB1xp67_ASAP7_75t_L g9485 ( 
.A(n_8969),
.Y(n_9485)
);

AND2x2_ASAP7_75t_L g9486 ( 
.A(n_8799),
.B(n_908),
.Y(n_9486)
);

INVx1_ASAP7_75t_L g9487 ( 
.A(n_8946),
.Y(n_9487)
);

NAND2xp5_ASAP7_75t_L g9488 ( 
.A(n_8801),
.B(n_909),
.Y(n_9488)
);

NAND2xp5_ASAP7_75t_SL g9489 ( 
.A(n_9027),
.B(n_909),
.Y(n_9489)
);

AOI22xp33_ASAP7_75t_L g9490 ( 
.A1(n_8608),
.A2(n_912),
.B1(n_910),
.B2(n_911),
.Y(n_9490)
);

NAND2xp5_ASAP7_75t_L g9491 ( 
.A(n_8804),
.B(n_910),
.Y(n_9491)
);

HB1xp67_ASAP7_75t_L g9492 ( 
.A(n_8645),
.Y(n_9492)
);

INVx2_ASAP7_75t_SL g9493 ( 
.A(n_8962),
.Y(n_9493)
);

BUFx6f_ASAP7_75t_L g9494 ( 
.A(n_8940),
.Y(n_9494)
);

AND2x4_ASAP7_75t_L g9495 ( 
.A(n_8750),
.B(n_911),
.Y(n_9495)
);

BUFx2_ASAP7_75t_L g9496 ( 
.A(n_8885),
.Y(n_9496)
);

AND2x4_ASAP7_75t_L g9497 ( 
.A(n_9108),
.B(n_8475),
.Y(n_9497)
);

BUFx3_ASAP7_75t_L g9498 ( 
.A(n_9031),
.Y(n_9498)
);

INVx1_ASAP7_75t_L g9499 ( 
.A(n_9100),
.Y(n_9499)
);

AOI21xp5_ASAP7_75t_L g9500 ( 
.A1(n_9429),
.A2(n_8514),
.B(n_8503),
.Y(n_9500)
);

AOI21xp5_ASAP7_75t_L g9501 ( 
.A1(n_9040),
.A2(n_8552),
.B(n_8547),
.Y(n_9501)
);

AO21x1_ASAP7_75t_L g9502 ( 
.A1(n_9249),
.A2(n_8761),
.B(n_8702),
.Y(n_9502)
);

NAND2xp5_ASAP7_75t_L g9503 ( 
.A(n_9365),
.B(n_8602),
.Y(n_9503)
);

AND2x2_ASAP7_75t_L g9504 ( 
.A(n_9052),
.B(n_8766),
.Y(n_9504)
);

BUFx3_ASAP7_75t_L g9505 ( 
.A(n_9144),
.Y(n_9505)
);

CKINVDCx20_ASAP7_75t_R g9506 ( 
.A(n_9054),
.Y(n_9506)
);

AO21x1_ASAP7_75t_L g9507 ( 
.A1(n_9192),
.A2(n_8713),
.B(n_8933),
.Y(n_9507)
);

AOI21xp5_ASAP7_75t_L g9508 ( 
.A1(n_9350),
.A2(n_8565),
.B(n_8554),
.Y(n_9508)
);

INVx5_ASAP7_75t_L g9509 ( 
.A(n_9110),
.Y(n_9509)
);

NAND2xp5_ASAP7_75t_L g9510 ( 
.A(n_9265),
.B(n_8492),
.Y(n_9510)
);

INVx1_ASAP7_75t_L g9511 ( 
.A(n_9123),
.Y(n_9511)
);

BUFx3_ASAP7_75t_L g9512 ( 
.A(n_9144),
.Y(n_9512)
);

AOI22xp33_ASAP7_75t_L g9513 ( 
.A1(n_9049),
.A2(n_8548),
.B1(n_8865),
.B2(n_8793),
.Y(n_9513)
);

NOR2xp33_ASAP7_75t_L g9514 ( 
.A(n_9294),
.B(n_8504),
.Y(n_9514)
);

INVx1_ASAP7_75t_L g9515 ( 
.A(n_9180),
.Y(n_9515)
);

BUFx3_ASAP7_75t_L g9516 ( 
.A(n_9155),
.Y(n_9516)
);

AND2x2_ASAP7_75t_L g9517 ( 
.A(n_9083),
.B(n_9264),
.Y(n_9517)
);

AND2x4_ASAP7_75t_L g9518 ( 
.A(n_9167),
.B(n_8741),
.Y(n_9518)
);

INVx2_ASAP7_75t_SL g9519 ( 
.A(n_9178),
.Y(n_9519)
);

AND2x4_ASAP7_75t_L g9520 ( 
.A(n_9216),
.B(n_8610),
.Y(n_9520)
);

INVx2_ASAP7_75t_L g9521 ( 
.A(n_9126),
.Y(n_9521)
);

AND2x2_ASAP7_75t_L g9522 ( 
.A(n_9050),
.B(n_8681),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_9189),
.Y(n_9523)
);

BUFx2_ASAP7_75t_L g9524 ( 
.A(n_9301),
.Y(n_9524)
);

INVx2_ASAP7_75t_L g9525 ( 
.A(n_9133),
.Y(n_9525)
);

NAND2xp5_ASAP7_75t_L g9526 ( 
.A(n_9280),
.B(n_8633),
.Y(n_9526)
);

NAND2xp5_ASAP7_75t_SL g9527 ( 
.A(n_9332),
.B(n_8883),
.Y(n_9527)
);

AOI21xp5_ASAP7_75t_L g9528 ( 
.A1(n_9163),
.A2(n_8576),
.B(n_8570),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_9151),
.B(n_8951),
.Y(n_9529)
);

BUFx4_ASAP7_75t_SL g9530 ( 
.A(n_9109),
.Y(n_9530)
);

INVxp67_ASAP7_75t_L g9531 ( 
.A(n_9316),
.Y(n_9531)
);

INVx2_ASAP7_75t_L g9532 ( 
.A(n_9136),
.Y(n_9532)
);

NAND2xp5_ASAP7_75t_L g9533 ( 
.A(n_9227),
.B(n_8808),
.Y(n_9533)
);

OR2x6_ASAP7_75t_L g9534 ( 
.A(n_9336),
.B(n_8579),
.Y(n_9534)
);

AND2x4_ASAP7_75t_L g9535 ( 
.A(n_9139),
.B(n_8818),
.Y(n_9535)
);

NAND3xp33_ASAP7_75t_L g9536 ( 
.A(n_9130),
.B(n_9187),
.C(n_9258),
.Y(n_9536)
);

AND2x4_ASAP7_75t_L g9537 ( 
.A(n_9105),
.B(n_8834),
.Y(n_9537)
);

INVx1_ASAP7_75t_SL g9538 ( 
.A(n_9232),
.Y(n_9538)
);

INVx2_ASAP7_75t_L g9539 ( 
.A(n_9143),
.Y(n_9539)
);

INVx2_ASAP7_75t_L g9540 ( 
.A(n_9158),
.Y(n_9540)
);

INVx2_ASAP7_75t_SL g9541 ( 
.A(n_9178),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_9036),
.Y(n_9542)
);

AOI21xp5_ASAP7_75t_L g9543 ( 
.A1(n_9489),
.A2(n_8486),
.B(n_8678),
.Y(n_9543)
);

INVx2_ASAP7_75t_L g9544 ( 
.A(n_9165),
.Y(n_9544)
);

OAI21x1_ASAP7_75t_L g9545 ( 
.A1(n_9378),
.A2(n_8669),
.B(n_8665),
.Y(n_9545)
);

BUFx6f_ASAP7_75t_L g9546 ( 
.A(n_9047),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_9038),
.Y(n_9547)
);

INVx5_ASAP7_75t_L g9548 ( 
.A(n_9110),
.Y(n_9548)
);

AND2x4_ASAP7_75t_L g9549 ( 
.A(n_9068),
.B(n_8835),
.Y(n_9549)
);

AND2x2_ASAP7_75t_L g9550 ( 
.A(n_9235),
.B(n_8895),
.Y(n_9550)
);

NAND2xp5_ASAP7_75t_L g9551 ( 
.A(n_9221),
.B(n_8921),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9039),
.Y(n_9552)
);

INVx1_ASAP7_75t_SL g9553 ( 
.A(n_9252),
.Y(n_9553)
);

INVx2_ASAP7_75t_L g9554 ( 
.A(n_9194),
.Y(n_9554)
);

INVx1_ASAP7_75t_L g9555 ( 
.A(n_9055),
.Y(n_9555)
);

OAI21x1_ASAP7_75t_L g9556 ( 
.A1(n_9409),
.A2(n_8767),
.B(n_8764),
.Y(n_9556)
);

INVx2_ASAP7_75t_L g9557 ( 
.A(n_9199),
.Y(n_9557)
);

HB1xp67_ASAP7_75t_L g9558 ( 
.A(n_9142),
.Y(n_9558)
);

INVx3_ASAP7_75t_L g9559 ( 
.A(n_9171),
.Y(n_9559)
);

INVx2_ASAP7_75t_SL g9560 ( 
.A(n_9172),
.Y(n_9560)
);

INVx3_ASAP7_75t_L g9561 ( 
.A(n_9204),
.Y(n_9561)
);

BUFx6f_ASAP7_75t_L g9562 ( 
.A(n_9047),
.Y(n_9562)
);

INVx1_ASAP7_75t_L g9563 ( 
.A(n_9066),
.Y(n_9563)
);

BUFx3_ASAP7_75t_L g9564 ( 
.A(n_9155),
.Y(n_9564)
);

BUFx6f_ASAP7_75t_L g9565 ( 
.A(n_9028),
.Y(n_9565)
);

AND2x4_ASAP7_75t_L g9566 ( 
.A(n_9197),
.B(n_8817),
.Y(n_9566)
);

CKINVDCx5p33_ASAP7_75t_R g9567 ( 
.A(n_9185),
.Y(n_9567)
);

NAND2xp5_ASAP7_75t_L g9568 ( 
.A(n_9341),
.B(n_8942),
.Y(n_9568)
);

AOI22xp33_ASAP7_75t_L g9569 ( 
.A1(n_9496),
.A2(n_8667),
.B1(n_8826),
.B2(n_8900),
.Y(n_9569)
);

INVxp67_ASAP7_75t_L g9570 ( 
.A(n_9257),
.Y(n_9570)
);

INVx4_ASAP7_75t_L g9571 ( 
.A(n_9134),
.Y(n_9571)
);

AOI21xp5_ASAP7_75t_L g9572 ( 
.A1(n_9309),
.A2(n_8489),
.B(n_8539),
.Y(n_9572)
);

OAI22xp5_ASAP7_75t_L g9573 ( 
.A1(n_9304),
.A2(n_8827),
.B1(n_8735),
.B2(n_8725),
.Y(n_9573)
);

NOR2xp33_ASAP7_75t_L g9574 ( 
.A(n_9349),
.B(n_8533),
.Y(n_9574)
);

AND2x2_ASAP7_75t_L g9575 ( 
.A(n_9051),
.B(n_8931),
.Y(n_9575)
);

CKINVDCx5p33_ASAP7_75t_R g9576 ( 
.A(n_9161),
.Y(n_9576)
);

INVx1_ASAP7_75t_L g9577 ( 
.A(n_9074),
.Y(n_9577)
);

BUFx2_ASAP7_75t_L g9578 ( 
.A(n_9261),
.Y(n_9578)
);

INVx3_ASAP7_75t_L g9579 ( 
.A(n_9204),
.Y(n_9579)
);

INVx1_ASAP7_75t_L g9580 ( 
.A(n_9076),
.Y(n_9580)
);

INVx3_ASAP7_75t_L g9581 ( 
.A(n_9125),
.Y(n_9581)
);

INVx2_ASAP7_75t_L g9582 ( 
.A(n_9208),
.Y(n_9582)
);

NAND2xp5_ASAP7_75t_L g9583 ( 
.A(n_9385),
.B(n_8967),
.Y(n_9583)
);

INVx2_ASAP7_75t_SL g9584 ( 
.A(n_9164),
.Y(n_9584)
);

INVx2_ASAP7_75t_L g9585 ( 
.A(n_9082),
.Y(n_9585)
);

INVx2_ASAP7_75t_SL g9586 ( 
.A(n_9224),
.Y(n_9586)
);

HB1xp67_ASAP7_75t_L g9587 ( 
.A(n_9281),
.Y(n_9587)
);

INVx2_ASAP7_75t_L g9588 ( 
.A(n_9120),
.Y(n_9588)
);

INVx3_ASAP7_75t_L g9589 ( 
.A(n_9228),
.Y(n_9589)
);

BUFx6f_ASAP7_75t_L g9590 ( 
.A(n_9028),
.Y(n_9590)
);

NAND2xp5_ASAP7_75t_L g9591 ( 
.A(n_9387),
.B(n_8692),
.Y(n_9591)
);

AND2x4_ASAP7_75t_L g9592 ( 
.A(n_9290),
.B(n_8851),
.Y(n_9592)
);

NAND2xp5_ASAP7_75t_L g9593 ( 
.A(n_9388),
.B(n_9441),
.Y(n_9593)
);

AND2x2_ASAP7_75t_L g9594 ( 
.A(n_9146),
.B(n_8974),
.Y(n_9594)
);

OA21x2_ASAP7_75t_L g9595 ( 
.A1(n_9312),
.A2(n_8980),
.B(n_8889),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_9078),
.Y(n_9596)
);

NAND2xp5_ASAP7_75t_L g9597 ( 
.A(n_9427),
.B(n_8695),
.Y(n_9597)
);

AND2x2_ASAP7_75t_L g9598 ( 
.A(n_9337),
.B(n_8553),
.Y(n_9598)
);

INVx1_ASAP7_75t_L g9599 ( 
.A(n_9102),
.Y(n_9599)
);

BUFx2_ASAP7_75t_L g9600 ( 
.A(n_9261),
.Y(n_9600)
);

INVx3_ASAP7_75t_L g9601 ( 
.A(n_9228),
.Y(n_9601)
);

NAND2xp5_ASAP7_75t_L g9602 ( 
.A(n_9392),
.B(n_8583),
.Y(n_9602)
);

BUFx6f_ASAP7_75t_L g9603 ( 
.A(n_9035),
.Y(n_9603)
);

BUFx6f_ASAP7_75t_L g9604 ( 
.A(n_9035),
.Y(n_9604)
);

INVx2_ASAP7_75t_L g9605 ( 
.A(n_9106),
.Y(n_9605)
);

AOI21xp5_ASAP7_75t_L g9606 ( 
.A1(n_9147),
.A2(n_8866),
.B(n_8525),
.Y(n_9606)
);

NAND2xp5_ASAP7_75t_L g9607 ( 
.A(n_9400),
.B(n_9411),
.Y(n_9607)
);

INVx1_ASAP7_75t_L g9608 ( 
.A(n_9115),
.Y(n_9608)
);

BUFx8_ASAP7_75t_SL g9609 ( 
.A(n_9213),
.Y(n_9609)
);

AND2x4_ASAP7_75t_L g9610 ( 
.A(n_9046),
.B(n_8747),
.Y(n_9610)
);

AND2x4_ASAP7_75t_L g9611 ( 
.A(n_9060),
.B(n_912),
.Y(n_9611)
);

CKINVDCx5p33_ASAP7_75t_R g9612 ( 
.A(n_9396),
.Y(n_9612)
);

CKINVDCx20_ASAP7_75t_R g9613 ( 
.A(n_9220),
.Y(n_9613)
);

NAND2xp5_ASAP7_75t_L g9614 ( 
.A(n_9412),
.B(n_8478),
.Y(n_9614)
);

BUFx3_ASAP7_75t_L g9615 ( 
.A(n_9030),
.Y(n_9615)
);

BUFx6f_ASAP7_75t_L g9616 ( 
.A(n_9072),
.Y(n_9616)
);

INVx1_ASAP7_75t_L g9617 ( 
.A(n_9131),
.Y(n_9617)
);

OAI21xp5_ASAP7_75t_L g9618 ( 
.A1(n_9255),
.A2(n_8666),
.B(n_8843),
.Y(n_9618)
);

O2A1O1Ixp5_ASAP7_75t_SL g9619 ( 
.A1(n_9445),
.A2(n_8970),
.B(n_8742),
.C(n_8882),
.Y(n_9619)
);

AOI21xp5_ASAP7_75t_L g9620 ( 
.A1(n_9196),
.A2(n_8715),
.B(n_8710),
.Y(n_9620)
);

AOI21xp5_ASAP7_75t_L g9621 ( 
.A1(n_9205),
.A2(n_8709),
.B(n_8718),
.Y(n_9621)
);

AOI21xp5_ASAP7_75t_L g9622 ( 
.A1(n_9363),
.A2(n_8787),
.B(n_8856),
.Y(n_9622)
);

NAND2xp5_ASAP7_75t_L g9623 ( 
.A(n_9413),
.B(n_8872),
.Y(n_9623)
);

BUFx3_ASAP7_75t_L g9624 ( 
.A(n_9042),
.Y(n_9624)
);

BUFx12f_ASAP7_75t_L g9625 ( 
.A(n_9073),
.Y(n_9625)
);

AND2x4_ASAP7_75t_L g9626 ( 
.A(n_9084),
.B(n_913),
.Y(n_9626)
);

A2O1A1Ixp33_ASAP7_75t_L g9627 ( 
.A1(n_9315),
.A2(n_8607),
.B(n_8614),
.C(n_8641),
.Y(n_9627)
);

OR2x2_ASAP7_75t_L g9628 ( 
.A(n_9307),
.B(n_8600),
.Y(n_9628)
);

INVx3_ASAP7_75t_L g9629 ( 
.A(n_9072),
.Y(n_9629)
);

AOI21xp5_ASAP7_75t_L g9630 ( 
.A1(n_9403),
.A2(n_8904),
.B(n_8828),
.Y(n_9630)
);

AOI21xp5_ASAP7_75t_L g9631 ( 
.A1(n_9203),
.A2(n_8953),
.B(n_8938),
.Y(n_9631)
);

BUFx2_ASAP7_75t_L g9632 ( 
.A(n_9261),
.Y(n_9632)
);

INVx3_ASAP7_75t_L g9633 ( 
.A(n_9080),
.Y(n_9633)
);

CKINVDCx20_ASAP7_75t_R g9634 ( 
.A(n_9097),
.Y(n_9634)
);

INVx5_ASAP7_75t_L g9635 ( 
.A(n_9278),
.Y(n_9635)
);

NAND2xp5_ASAP7_75t_L g9636 ( 
.A(n_9415),
.B(n_9423),
.Y(n_9636)
);

INVx1_ASAP7_75t_L g9637 ( 
.A(n_9132),
.Y(n_9637)
);

AND2x2_ASAP7_75t_L g9638 ( 
.A(n_9421),
.B(n_914),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_9153),
.Y(n_9639)
);

INVx2_ASAP7_75t_L g9640 ( 
.A(n_9162),
.Y(n_9640)
);

BUFx10_ASAP7_75t_L g9641 ( 
.A(n_9201),
.Y(n_9641)
);

BUFx2_ASAP7_75t_SL g9642 ( 
.A(n_9134),
.Y(n_9642)
);

OAI22xp5_ASAP7_75t_L g9643 ( 
.A1(n_9285),
.A2(n_916),
.B1(n_914),
.B2(n_915),
.Y(n_9643)
);

INVx3_ASAP7_75t_L g9644 ( 
.A(n_9080),
.Y(n_9644)
);

AOI21xp5_ASAP7_75t_L g9645 ( 
.A1(n_9346),
.A2(n_915),
.B(n_917),
.Y(n_9645)
);

A2O1A1Ixp33_ASAP7_75t_L g9646 ( 
.A1(n_9174),
.A2(n_919),
.B(n_917),
.C(n_918),
.Y(n_9646)
);

AND2x2_ASAP7_75t_L g9647 ( 
.A(n_9333),
.B(n_918),
.Y(n_9647)
);

NAND2xp5_ASAP7_75t_SL g9648 ( 
.A(n_9310),
.B(n_919),
.Y(n_9648)
);

INVx1_ASAP7_75t_L g9649 ( 
.A(n_9170),
.Y(n_9649)
);

INVx2_ASAP7_75t_L g9650 ( 
.A(n_9177),
.Y(n_9650)
);

AOI221x1_ASAP7_75t_L g9651 ( 
.A1(n_9436),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.C(n_923),
.Y(n_9651)
);

INVx2_ASAP7_75t_L g9652 ( 
.A(n_9179),
.Y(n_9652)
);

INVx2_ASAP7_75t_SL g9653 ( 
.A(n_9215),
.Y(n_9653)
);

BUFx12f_ASAP7_75t_L g9654 ( 
.A(n_9182),
.Y(n_9654)
);

INVx1_ASAP7_75t_L g9655 ( 
.A(n_9184),
.Y(n_9655)
);

BUFx2_ASAP7_75t_L g9656 ( 
.A(n_9313),
.Y(n_9656)
);

OAI22xp5_ASAP7_75t_L g9657 ( 
.A1(n_9181),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.Y(n_9657)
);

INVx1_ASAP7_75t_L g9658 ( 
.A(n_9191),
.Y(n_9658)
);

AND2x2_ASAP7_75t_L g9659 ( 
.A(n_9393),
.B(n_924),
.Y(n_9659)
);

AOI21xp5_ASAP7_75t_L g9660 ( 
.A1(n_9466),
.A2(n_925),
.B(n_926),
.Y(n_9660)
);

AND2x4_ASAP7_75t_L g9661 ( 
.A(n_9112),
.B(n_926),
.Y(n_9661)
);

NAND2xp33_ASAP7_75t_L g9662 ( 
.A(n_9044),
.B(n_927),
.Y(n_9662)
);

AOI22xp33_ASAP7_75t_L g9663 ( 
.A1(n_9217),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.Y(n_9663)
);

INVx3_ASAP7_75t_L g9664 ( 
.A(n_9103),
.Y(n_9664)
);

OAI22xp5_ASAP7_75t_L g9665 ( 
.A1(n_9064),
.A2(n_932),
.B1(n_929),
.B2(n_930),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_9202),
.Y(n_9666)
);

OAI21xp5_ASAP7_75t_L g9667 ( 
.A1(n_9475),
.A2(n_930),
.B(n_932),
.Y(n_9667)
);

INVx1_ASAP7_75t_L g9668 ( 
.A(n_9226),
.Y(n_9668)
);

INVxp67_ASAP7_75t_SL g9669 ( 
.A(n_9193),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_L g9670 ( 
.A(n_9395),
.B(n_933),
.Y(n_9670)
);

OR2x2_ASAP7_75t_L g9671 ( 
.A(n_9234),
.B(n_934),
.Y(n_9671)
);

AO32x1_ASAP7_75t_L g9672 ( 
.A1(n_9034),
.A2(n_936),
.A3(n_934),
.B1(n_935),
.B2(n_937),
.Y(n_9672)
);

AOI21x1_ASAP7_75t_L g9673 ( 
.A1(n_9242),
.A2(n_935),
.B(n_936),
.Y(n_9673)
);

AOI21xp5_ASAP7_75t_L g9674 ( 
.A1(n_9268),
.A2(n_937),
.B(n_938),
.Y(n_9674)
);

AND2x4_ASAP7_75t_L g9675 ( 
.A(n_9114),
.B(n_938),
.Y(n_9675)
);

AND2x4_ASAP7_75t_L g9676 ( 
.A(n_9246),
.B(n_9251),
.Y(n_9676)
);

INVx5_ASAP7_75t_L g9677 ( 
.A(n_9278),
.Y(n_9677)
);

NAND2xp5_ASAP7_75t_L g9678 ( 
.A(n_9422),
.B(n_939),
.Y(n_9678)
);

AO21x1_ASAP7_75t_L g9679 ( 
.A1(n_9371),
.A2(n_939),
.B(n_940),
.Y(n_9679)
);

NAND2xp5_ASAP7_75t_L g9680 ( 
.A(n_9318),
.B(n_940),
.Y(n_9680)
);

INVx2_ASAP7_75t_SL g9681 ( 
.A(n_9215),
.Y(n_9681)
);

NAND2x1p5_ASAP7_75t_L g9682 ( 
.A(n_9310),
.B(n_941),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_9241),
.Y(n_9683)
);

NAND2x1p5_ASAP7_75t_L g9684 ( 
.A(n_9420),
.B(n_941),
.Y(n_9684)
);

AND2x2_ASAP7_75t_L g9685 ( 
.A(n_9317),
.B(n_942),
.Y(n_9685)
);

INVx2_ASAP7_75t_SL g9686 ( 
.A(n_9186),
.Y(n_9686)
);

NAND2xp5_ASAP7_75t_L g9687 ( 
.A(n_9338),
.B(n_942),
.Y(n_9687)
);

CKINVDCx5p33_ASAP7_75t_R g9688 ( 
.A(n_9414),
.Y(n_9688)
);

INVx1_ASAP7_75t_L g9689 ( 
.A(n_9273),
.Y(n_9689)
);

OR2x2_ASAP7_75t_L g9690 ( 
.A(n_9267),
.B(n_943),
.Y(n_9690)
);

AND2x2_ASAP7_75t_L g9691 ( 
.A(n_9394),
.B(n_943),
.Y(n_9691)
);

INVx1_ASAP7_75t_L g9692 ( 
.A(n_9275),
.Y(n_9692)
);

O2A1O1Ixp5_ASAP7_75t_L g9693 ( 
.A1(n_9104),
.A2(n_946),
.B(n_944),
.C(n_945),
.Y(n_9693)
);

AOI21xp5_ASAP7_75t_L g9694 ( 
.A1(n_9383),
.A2(n_944),
.B(n_945),
.Y(n_9694)
);

AND2x4_ASAP7_75t_L g9695 ( 
.A(n_9295),
.B(n_947),
.Y(n_9695)
);

AND2x4_ASAP7_75t_L g9696 ( 
.A(n_9303),
.B(n_947),
.Y(n_9696)
);

NAND2xp5_ASAP7_75t_L g9697 ( 
.A(n_9344),
.B(n_948),
.Y(n_9697)
);

NAND2xp5_ASAP7_75t_L g9698 ( 
.A(n_9353),
.B(n_9354),
.Y(n_9698)
);

INVx2_ASAP7_75t_L g9699 ( 
.A(n_9306),
.Y(n_9699)
);

BUFx6f_ASAP7_75t_L g9700 ( 
.A(n_9103),
.Y(n_9700)
);

OR2x2_ASAP7_75t_L g9701 ( 
.A(n_9428),
.B(n_948),
.Y(n_9701)
);

OAI22xp5_ASAP7_75t_SL g9702 ( 
.A1(n_9381),
.A2(n_951),
.B1(n_949),
.B2(n_950),
.Y(n_9702)
);

INVx1_ASAP7_75t_L g9703 ( 
.A(n_9239),
.Y(n_9703)
);

OAI22xp33_ASAP7_75t_L g9704 ( 
.A1(n_9176),
.A2(n_951),
.B1(n_949),
.B2(n_950),
.Y(n_9704)
);

AND2x2_ASAP7_75t_L g9705 ( 
.A(n_9391),
.B(n_952),
.Y(n_9705)
);

NAND2xp5_ASAP7_75t_L g9706 ( 
.A(n_9424),
.B(n_953),
.Y(n_9706)
);

NAND2xp5_ASAP7_75t_L g9707 ( 
.A(n_9358),
.B(n_953),
.Y(n_9707)
);

BUFx2_ASAP7_75t_L g9708 ( 
.A(n_9313),
.Y(n_9708)
);

NAND2xp5_ASAP7_75t_L g9709 ( 
.A(n_9448),
.B(n_954),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_9298),
.Y(n_9710)
);

BUFx2_ASAP7_75t_L g9711 ( 
.A(n_9321),
.Y(n_9711)
);

AOI22xp33_ASAP7_75t_SL g9712 ( 
.A1(n_9320),
.A2(n_958),
.B1(n_955),
.B2(n_956),
.Y(n_9712)
);

NOR3xp33_ASAP7_75t_L g9713 ( 
.A(n_9484),
.B(n_955),
.C(n_956),
.Y(n_9713)
);

AND2x2_ASAP7_75t_L g9714 ( 
.A(n_9399),
.B(n_959),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_9305),
.Y(n_9715)
);

INVx1_ASAP7_75t_L g9716 ( 
.A(n_9390),
.Y(n_9716)
);

AND2x2_ASAP7_75t_L g9717 ( 
.A(n_9272),
.B(n_960),
.Y(n_9717)
);

INVx5_ASAP7_75t_L g9718 ( 
.A(n_9278),
.Y(n_9718)
);

NAND2xp5_ASAP7_75t_L g9719 ( 
.A(n_9483),
.B(n_961),
.Y(n_9719)
);

O2A1O1Ixp33_ASAP7_75t_L g9720 ( 
.A1(n_9124),
.A2(n_964),
.B(n_962),
.C(n_963),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9382),
.Y(n_9721)
);

OAI22xp5_ASAP7_75t_L g9722 ( 
.A1(n_9269),
.A2(n_964),
.B1(n_962),
.B2(n_963),
.Y(n_9722)
);

CKINVDCx8_ASAP7_75t_R g9723 ( 
.A(n_9435),
.Y(n_9723)
);

INVx5_ASAP7_75t_L g9724 ( 
.A(n_9372),
.Y(n_9724)
);

AOI22xp33_ASAP7_75t_L g9725 ( 
.A1(n_9482),
.A2(n_967),
.B1(n_965),
.B2(n_966),
.Y(n_9725)
);

O2A1O1Ixp5_ASAP7_75t_SL g9726 ( 
.A1(n_9360),
.A2(n_968),
.B(n_965),
.C(n_966),
.Y(n_9726)
);

NAND2xp5_ASAP7_75t_L g9727 ( 
.A(n_9299),
.B(n_968),
.Y(n_9727)
);

NAND2xp5_ASAP7_75t_L g9728 ( 
.A(n_9443),
.B(n_969),
.Y(n_9728)
);

INVx1_ASAP7_75t_L g9729 ( 
.A(n_9335),
.Y(n_9729)
);

HB1xp67_ASAP7_75t_L g9730 ( 
.A(n_9288),
.Y(n_9730)
);

INVxp67_ASAP7_75t_SL g9731 ( 
.A(n_9284),
.Y(n_9731)
);

BUFx3_ASAP7_75t_L g9732 ( 
.A(n_9053),
.Y(n_9732)
);

BUFx6f_ASAP7_75t_L g9733 ( 
.A(n_9137),
.Y(n_9733)
);

OAI22xp5_ASAP7_75t_L g9734 ( 
.A1(n_9253),
.A2(n_972),
.B1(n_970),
.B2(n_971),
.Y(n_9734)
);

INVxp67_ASAP7_75t_L g9735 ( 
.A(n_9434),
.Y(n_9735)
);

BUFx12f_ASAP7_75t_L g9736 ( 
.A(n_9168),
.Y(n_9736)
);

OR2x2_ASAP7_75t_L g9737 ( 
.A(n_9037),
.B(n_970),
.Y(n_9737)
);

INVx1_ASAP7_75t_L g9738 ( 
.A(n_9364),
.Y(n_9738)
);

INVx3_ASAP7_75t_L g9739 ( 
.A(n_9137),
.Y(n_9739)
);

NOR2xp33_ASAP7_75t_L g9740 ( 
.A(n_9473),
.B(n_971),
.Y(n_9740)
);

A2O1A1Ixp33_ASAP7_75t_SL g9741 ( 
.A1(n_9471),
.A2(n_974),
.B(n_972),
.C(n_973),
.Y(n_9741)
);

NAND2xp5_ASAP7_75t_L g9742 ( 
.A(n_9487),
.B(n_9322),
.Y(n_9742)
);

NAND2xp5_ASAP7_75t_L g9743 ( 
.A(n_9367),
.B(n_974),
.Y(n_9743)
);

INVx2_ASAP7_75t_L g9744 ( 
.A(n_9284),
.Y(n_9744)
);

OR2x2_ASAP7_75t_L g9745 ( 
.A(n_9067),
.B(n_976),
.Y(n_9745)
);

INVx3_ASAP7_75t_L g9746 ( 
.A(n_9223),
.Y(n_9746)
);

AND2x2_ASAP7_75t_L g9747 ( 
.A(n_9198),
.B(n_977),
.Y(n_9747)
);

OAI22xp5_ASAP7_75t_L g9748 ( 
.A1(n_9135),
.A2(n_980),
.B1(n_978),
.B2(n_979),
.Y(n_9748)
);

INVx4_ASAP7_75t_L g9749 ( 
.A(n_9057),
.Y(n_9749)
);

AOI21xp5_ASAP7_75t_L g9750 ( 
.A1(n_9148),
.A2(n_978),
.B(n_979),
.Y(n_9750)
);

AOI21xp5_ASAP7_75t_L g9751 ( 
.A1(n_9470),
.A2(n_981),
.B(n_983),
.Y(n_9751)
);

NAND2xp5_ASAP7_75t_L g9752 ( 
.A(n_9367),
.B(n_983),
.Y(n_9752)
);

INVx2_ASAP7_75t_L g9753 ( 
.A(n_9366),
.Y(n_9753)
);

CKINVDCx5p33_ASAP7_75t_R g9754 ( 
.A(n_9166),
.Y(n_9754)
);

A2O1A1Ixp33_ASAP7_75t_L g9755 ( 
.A1(n_9348),
.A2(n_986),
.B(n_984),
.C(n_985),
.Y(n_9755)
);

INVx1_ASAP7_75t_L g9756 ( 
.A(n_9373),
.Y(n_9756)
);

AOI22xp33_ASAP7_75t_L g9757 ( 
.A1(n_9432),
.A2(n_987),
.B1(n_985),
.B2(n_986),
.Y(n_9757)
);

INVx2_ASAP7_75t_L g9758 ( 
.A(n_9359),
.Y(n_9758)
);

BUFx3_ASAP7_75t_L g9759 ( 
.A(n_9058),
.Y(n_9759)
);

INVx1_ASAP7_75t_L g9760 ( 
.A(n_9370),
.Y(n_9760)
);

NAND2xp5_ASAP7_75t_L g9761 ( 
.A(n_9463),
.B(n_987),
.Y(n_9761)
);

AND2x2_ASAP7_75t_L g9762 ( 
.A(n_9200),
.B(n_988),
.Y(n_9762)
);

AND2x2_ASAP7_75t_SL g9763 ( 
.A(n_9248),
.B(n_989),
.Y(n_9763)
);

NAND2xp5_ASAP7_75t_L g9764 ( 
.A(n_9321),
.B(n_990),
.Y(n_9764)
);

AND2x4_ASAP7_75t_L g9765 ( 
.A(n_9233),
.B(n_990),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9374),
.B(n_991),
.Y(n_9766)
);

AOI22xp33_ASAP7_75t_L g9767 ( 
.A1(n_9033),
.A2(n_993),
.B1(n_991),
.B2(n_992),
.Y(n_9767)
);

INVx2_ASAP7_75t_L g9768 ( 
.A(n_9455),
.Y(n_9768)
);

BUFx3_ASAP7_75t_L g9769 ( 
.A(n_9088),
.Y(n_9769)
);

OR2x6_ASAP7_75t_L g9770 ( 
.A(n_9345),
.B(n_992),
.Y(n_9770)
);

HB1xp67_ASAP7_75t_L g9771 ( 
.A(n_9485),
.Y(n_9771)
);

A2O1A1Ixp33_ASAP7_75t_SL g9772 ( 
.A1(n_9474),
.A2(n_995),
.B(n_993),
.C(n_994),
.Y(n_9772)
);

AOI22xp33_ASAP7_75t_L g9773 ( 
.A1(n_9495),
.A2(n_997),
.B1(n_994),
.B2(n_996),
.Y(n_9773)
);

INVx3_ASAP7_75t_L g9774 ( 
.A(n_9308),
.Y(n_9774)
);

A2O1A1Ixp33_ASAP7_75t_L g9775 ( 
.A1(n_9048),
.A2(n_999),
.B(n_997),
.C(n_998),
.Y(n_9775)
);

OA21x2_ASAP7_75t_L g9776 ( 
.A1(n_9478),
.A2(n_998),
.B(n_999),
.Y(n_9776)
);

OR2x2_ASAP7_75t_L g9777 ( 
.A(n_9458),
.B(n_1000),
.Y(n_9777)
);

AND2x2_ASAP7_75t_L g9778 ( 
.A(n_9434),
.B(n_1000),
.Y(n_9778)
);

BUFx12f_ASAP7_75t_L g9779 ( 
.A(n_9209),
.Y(n_9779)
);

AND2x4_ASAP7_75t_L g9780 ( 
.A(n_9323),
.B(n_1001),
.Y(n_9780)
);

HB1xp67_ASAP7_75t_L g9781 ( 
.A(n_9492),
.Y(n_9781)
);

BUFx2_ASAP7_75t_L g9782 ( 
.A(n_9308),
.Y(n_9782)
);

AOI21x1_ASAP7_75t_L g9783 ( 
.A1(n_9327),
.A2(n_1001),
.B(n_1002),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9090),
.Y(n_9784)
);

NAND2xp5_ASAP7_75t_L g9785 ( 
.A(n_9460),
.B(n_1002),
.Y(n_9785)
);

INVx1_ASAP7_75t_L g9786 ( 
.A(n_9293),
.Y(n_9786)
);

AND2x4_ASAP7_75t_L g9787 ( 
.A(n_9156),
.B(n_1003),
.Y(n_9787)
);

INVx2_ASAP7_75t_SL g9788 ( 
.A(n_9244),
.Y(n_9788)
);

AOI21xp5_ASAP7_75t_L g9789 ( 
.A1(n_9141),
.A2(n_1004),
.B(n_1005),
.Y(n_9789)
);

OAI22xp5_ASAP7_75t_SL g9790 ( 
.A1(n_9159),
.A2(n_1006),
.B1(n_1004),
.B2(n_1005),
.Y(n_9790)
);

AND2x2_ASAP7_75t_L g9791 ( 
.A(n_9450),
.B(n_1006),
.Y(n_9791)
);

INVx2_ASAP7_75t_L g9792 ( 
.A(n_9450),
.Y(n_9792)
);

AND2x4_ASAP7_75t_L g9793 ( 
.A(n_9157),
.B(n_1007),
.Y(n_9793)
);

CKINVDCx5p33_ASAP7_75t_R g9794 ( 
.A(n_9236),
.Y(n_9794)
);

INVx1_ASAP7_75t_L g9795 ( 
.A(n_9099),
.Y(n_9795)
);

AOI21xp5_ASAP7_75t_L g9796 ( 
.A1(n_9141),
.A2(n_1007),
.B(n_1009),
.Y(n_9796)
);

BUFx2_ASAP7_75t_L g9797 ( 
.A(n_9183),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_9061),
.Y(n_9798)
);

INVx2_ASAP7_75t_L g9799 ( 
.A(n_9069),
.Y(n_9799)
);

INVx3_ASAP7_75t_L g9800 ( 
.A(n_9085),
.Y(n_9800)
);

AOI21xp33_ASAP7_75t_SL g9801 ( 
.A1(n_9101),
.A2(n_1009),
.B(n_1010),
.Y(n_9801)
);

OAI21xp33_ASAP7_75t_L g9802 ( 
.A1(n_9467),
.A2(n_1011),
.B(n_1012),
.Y(n_9802)
);

INVx2_ASAP7_75t_L g9803 ( 
.A(n_9081),
.Y(n_9803)
);

INVx4_ASAP7_75t_L g9804 ( 
.A(n_9140),
.Y(n_9804)
);

INVx1_ASAP7_75t_L g9805 ( 
.A(n_9063),
.Y(n_9805)
);

BUFx3_ASAP7_75t_L g9806 ( 
.A(n_9219),
.Y(n_9806)
);

INVx1_ASAP7_75t_L g9807 ( 
.A(n_9089),
.Y(n_9807)
);

INVxp67_ASAP7_75t_L g9808 ( 
.A(n_9419),
.Y(n_9808)
);

HAxp5_ASAP7_75t_L g9809 ( 
.A(n_9449),
.B(n_1011),
.CON(n_9809),
.SN(n_9809)
);

INVx2_ASAP7_75t_L g9810 ( 
.A(n_9121),
.Y(n_9810)
);

AOI22xp33_ASAP7_75t_L g9811 ( 
.A1(n_9465),
.A2(n_1014),
.B1(n_1012),
.B2(n_1013),
.Y(n_9811)
);

AND2x2_ASAP7_75t_L g9812 ( 
.A(n_9356),
.B(n_9376),
.Y(n_9812)
);

BUFx2_ASAP7_75t_L g9813 ( 
.A(n_9214),
.Y(n_9813)
);

AND2x2_ASAP7_75t_L g9814 ( 
.A(n_9451),
.B(n_1014),
.Y(n_9814)
);

OAI22xp5_ASAP7_75t_L g9815 ( 
.A1(n_9218),
.A2(n_1018),
.B1(n_1016),
.B2(n_1017),
.Y(n_9815)
);

AOI21xp5_ASAP7_75t_L g9816 ( 
.A1(n_9375),
.A2(n_1016),
.B(n_1017),
.Y(n_9816)
);

INVx1_ASAP7_75t_SL g9817 ( 
.A(n_9222),
.Y(n_9817)
);

NAND2xp5_ASAP7_75t_L g9818 ( 
.A(n_9472),
.B(n_1019),
.Y(n_9818)
);

NAND2xp5_ASAP7_75t_L g9819 ( 
.A(n_9154),
.B(n_1019),
.Y(n_9819)
);

INVx1_ASAP7_75t_L g9820 ( 
.A(n_9119),
.Y(n_9820)
);

BUFx2_ASAP7_75t_L g9821 ( 
.A(n_9095),
.Y(n_9821)
);

AOI21xp5_ASAP7_75t_L g9822 ( 
.A1(n_9062),
.A2(n_1020),
.B(n_1021),
.Y(n_9822)
);

NAND2xp5_ASAP7_75t_L g9823 ( 
.A(n_9325),
.B(n_1020),
.Y(n_9823)
);

AND2x2_ASAP7_75t_L g9824 ( 
.A(n_9145),
.B(n_1021),
.Y(n_9824)
);

NAND2x1p5_ASAP7_75t_L g9825 ( 
.A(n_9343),
.B(n_1022),
.Y(n_9825)
);

NAND2xp5_ASAP7_75t_L g9826 ( 
.A(n_9071),
.B(n_1022),
.Y(n_9826)
);

INVx2_ASAP7_75t_L g9827 ( 
.A(n_9087),
.Y(n_9827)
);

INVxp67_ASAP7_75t_L g9828 ( 
.A(n_9416),
.Y(n_9828)
);

A2O1A1Ixp33_ASAP7_75t_L g9829 ( 
.A1(n_9231),
.A2(n_9404),
.B(n_9425),
.C(n_9362),
.Y(n_9829)
);

A2O1A1Ixp33_ASAP7_75t_SL g9830 ( 
.A1(n_9250),
.A2(n_1025),
.B(n_1023),
.C(n_1024),
.Y(n_9830)
);

INVx1_ASAP7_75t_L g9831 ( 
.A(n_9150),
.Y(n_9831)
);

INVx3_ASAP7_75t_L g9832 ( 
.A(n_9092),
.Y(n_9832)
);

INVx3_ASAP7_75t_L g9833 ( 
.A(n_9138),
.Y(n_9833)
);

INVx2_ASAP7_75t_L g9834 ( 
.A(n_9093),
.Y(n_9834)
);

BUFx5_ASAP7_75t_L g9835 ( 
.A(n_9372),
.Y(n_9835)
);

BUFx3_ASAP7_75t_L g9836 ( 
.A(n_9045),
.Y(n_9836)
);

AOI21xp5_ASAP7_75t_L g9837 ( 
.A1(n_9160),
.A2(n_1024),
.B(n_1025),
.Y(n_9837)
);

OR2x2_ASAP7_75t_L g9838 ( 
.A(n_9079),
.B(n_1026),
.Y(n_9838)
);

AOI222xp33_ASAP7_75t_L g9839 ( 
.A1(n_9225),
.A2(n_1028),
.B1(n_1030),
.B2(n_1026),
.C1(n_1027),
.C2(n_1029),
.Y(n_9839)
);

NOR2xp67_ASAP7_75t_SL g9840 ( 
.A(n_9212),
.B(n_1027),
.Y(n_9840)
);

INVx2_ASAP7_75t_L g9841 ( 
.A(n_9094),
.Y(n_9841)
);

NAND2xp5_ASAP7_75t_L g9842 ( 
.A(n_9043),
.B(n_1030),
.Y(n_9842)
);

AND2x4_ASAP7_75t_L g9843 ( 
.A(n_9117),
.B(n_1031),
.Y(n_9843)
);

INVx3_ASAP7_75t_L g9844 ( 
.A(n_9065),
.Y(n_9844)
);

INVx1_ASAP7_75t_L g9845 ( 
.A(n_9169),
.Y(n_9845)
);

INVx3_ASAP7_75t_SL g9846 ( 
.A(n_9271),
.Y(n_9846)
);

AOI21xp33_ASAP7_75t_L g9847 ( 
.A1(n_9127),
.A2(n_1031),
.B(n_1032),
.Y(n_9847)
);

BUFx3_ASAP7_75t_L g9848 ( 
.A(n_9077),
.Y(n_9848)
);

INVx5_ASAP7_75t_L g9849 ( 
.A(n_9372),
.Y(n_9849)
);

BUFx6f_ASAP7_75t_L g9850 ( 
.A(n_9238),
.Y(n_9850)
);

AND2x4_ASAP7_75t_L g9851 ( 
.A(n_9262),
.B(n_1033),
.Y(n_9851)
);

NAND2xp5_ASAP7_75t_L g9852 ( 
.A(n_9128),
.B(n_1033),
.Y(n_9852)
);

INVx1_ASAP7_75t_L g9853 ( 
.A(n_9173),
.Y(n_9853)
);

BUFx3_ASAP7_75t_L g9854 ( 
.A(n_9238),
.Y(n_9854)
);

AOI21xp5_ASAP7_75t_L g9855 ( 
.A1(n_9369),
.A2(n_1034),
.B(n_1035),
.Y(n_9855)
);

HB1xp67_ASAP7_75t_L g9856 ( 
.A(n_9493),
.Y(n_9856)
);

INVx2_ASAP7_75t_L g9857 ( 
.A(n_9276),
.Y(n_9857)
);

INVx3_ASAP7_75t_L g9858 ( 
.A(n_9243),
.Y(n_9858)
);

INVx3_ASAP7_75t_L g9859 ( 
.A(n_9245),
.Y(n_9859)
);

AOI21xp5_ASAP7_75t_L g9860 ( 
.A1(n_9437),
.A2(n_1034),
.B(n_1035),
.Y(n_9860)
);

AND2x2_ASAP7_75t_SL g9861 ( 
.A(n_9324),
.B(n_1036),
.Y(n_9861)
);

INVx1_ASAP7_75t_L g9862 ( 
.A(n_9206),
.Y(n_9862)
);

NAND2xp5_ASAP7_75t_L g9863 ( 
.A(n_9098),
.B(n_1036),
.Y(n_9863)
);

INVx2_ASAP7_75t_L g9864 ( 
.A(n_9282),
.Y(n_9864)
);

O2A1O1Ixp33_ASAP7_75t_SL g9865 ( 
.A1(n_9380),
.A2(n_1039),
.B(n_1037),
.C(n_1038),
.Y(n_9865)
);

AOI21xp5_ASAP7_75t_L g9866 ( 
.A1(n_9477),
.A2(n_1038),
.B(n_1039),
.Y(n_9866)
);

O2A1O1Ixp33_ASAP7_75t_L g9867 ( 
.A1(n_9056),
.A2(n_1042),
.B(n_1040),
.C(n_1041),
.Y(n_9867)
);

BUFx2_ASAP7_75t_L g9868 ( 
.A(n_9283),
.Y(n_9868)
);

BUFx6f_ASAP7_75t_L g9869 ( 
.A(n_9111),
.Y(n_9869)
);

OR2x6_ASAP7_75t_L g9870 ( 
.A(n_9032),
.B(n_1040),
.Y(n_9870)
);

INVx1_ASAP7_75t_L g9871 ( 
.A(n_9211),
.Y(n_9871)
);

AOI22xp5_ASAP7_75t_L g9872 ( 
.A1(n_9044),
.A2(n_1044),
.B1(n_1042),
.B2(n_1043),
.Y(n_9872)
);

AO22x2_ASAP7_75t_L g9873 ( 
.A1(n_9091),
.A2(n_1045),
.B1(n_1043),
.B2(n_1044),
.Y(n_9873)
);

NOR2xp33_ASAP7_75t_L g9874 ( 
.A(n_9431),
.B(n_1045),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_9738),
.Y(n_9875)
);

OAI22xp5_ASAP7_75t_L g9876 ( 
.A1(n_9569),
.A2(n_9188),
.B1(n_9096),
.B2(n_9452),
.Y(n_9876)
);

AOI22xp33_ASAP7_75t_L g9877 ( 
.A1(n_9536),
.A2(n_9292),
.B1(n_9494),
.B2(n_9044),
.Y(n_9877)
);

INVx4_ASAP7_75t_L g9878 ( 
.A(n_9509),
.Y(n_9878)
);

INVx2_ASAP7_75t_L g9879 ( 
.A(n_9524),
.Y(n_9879)
);

AOI22xp33_ASAP7_75t_L g9880 ( 
.A1(n_9507),
.A2(n_9494),
.B1(n_9479),
.B2(n_9408),
.Y(n_9880)
);

AOI22xp33_ASAP7_75t_SL g9881 ( 
.A1(n_9662),
.A2(n_9129),
.B1(n_9468),
.B2(n_9397),
.Y(n_9881)
);

OAI22xp5_ASAP7_75t_L g9882 ( 
.A1(n_9513),
.A2(n_9274),
.B1(n_9447),
.B2(n_9329),
.Y(n_9882)
);

CKINVDCx6p67_ASAP7_75t_R g9883 ( 
.A(n_9509),
.Y(n_9883)
);

OAI22xp5_ASAP7_75t_SL g9884 ( 
.A1(n_9790),
.A2(n_9548),
.B1(n_9702),
.B2(n_9763),
.Y(n_9884)
);

AOI22xp33_ASAP7_75t_SL g9885 ( 
.A1(n_9573),
.A2(n_9468),
.B1(n_9122),
.B2(n_9446),
.Y(n_9885)
);

BUFx3_ASAP7_75t_L g9886 ( 
.A(n_9634),
.Y(n_9886)
);

AOI22xp33_ASAP7_75t_L g9887 ( 
.A1(n_9502),
.A2(n_9152),
.B1(n_9456),
.B2(n_9407),
.Y(n_9887)
);

INVx1_ASAP7_75t_SL g9888 ( 
.A(n_9530),
.Y(n_9888)
);

OAI22xp33_ASAP7_75t_SL g9889 ( 
.A1(n_9724),
.A2(n_9433),
.B1(n_9229),
.B2(n_9476),
.Y(n_9889)
);

INVx1_ASAP7_75t_L g9890 ( 
.A(n_9756),
.Y(n_9890)
);

INVx2_ASAP7_75t_SL g9891 ( 
.A(n_9548),
.Y(n_9891)
);

INVx2_ASAP7_75t_L g9892 ( 
.A(n_9605),
.Y(n_9892)
);

INVx3_ASAP7_75t_L g9893 ( 
.A(n_9806),
.Y(n_9893)
);

OAI21xp5_ASAP7_75t_SL g9894 ( 
.A1(n_9621),
.A2(n_9190),
.B(n_9352),
.Y(n_9894)
);

AOI22xp33_ASAP7_75t_SL g9895 ( 
.A1(n_9724),
.A2(n_9118),
.B1(n_9459),
.B2(n_9384),
.Y(n_9895)
);

BUFx12f_ASAP7_75t_L g9896 ( 
.A(n_9612),
.Y(n_9896)
);

INVx2_ASAP7_75t_L g9897 ( 
.A(n_9640),
.Y(n_9897)
);

INVx1_ASAP7_75t_L g9898 ( 
.A(n_9668),
.Y(n_9898)
);

INVx2_ASAP7_75t_L g9899 ( 
.A(n_9650),
.Y(n_9899)
);

INVx1_ASAP7_75t_L g9900 ( 
.A(n_9683),
.Y(n_9900)
);

NAND2xp5_ASAP7_75t_L g9901 ( 
.A(n_9771),
.B(n_9041),
.Y(n_9901)
);

INVx6_ASAP7_75t_L g9902 ( 
.A(n_9625),
.Y(n_9902)
);

INVx1_ASAP7_75t_L g9903 ( 
.A(n_9542),
.Y(n_9903)
);

INVx2_ASAP7_75t_L g9904 ( 
.A(n_9652),
.Y(n_9904)
);

OAI22xp5_ASAP7_75t_L g9905 ( 
.A1(n_9663),
.A2(n_9254),
.B1(n_9195),
.B2(n_9490),
.Y(n_9905)
);

BUFx12f_ASAP7_75t_L g9906 ( 
.A(n_9794),
.Y(n_9906)
);

OAI22xp5_ASAP7_75t_L g9907 ( 
.A1(n_9849),
.A2(n_9175),
.B1(n_9444),
.B2(n_9439),
.Y(n_9907)
);

NAND2x1p5_ASAP7_75t_L g9908 ( 
.A(n_9635),
.B(n_9677),
.Y(n_9908)
);

CKINVDCx20_ASAP7_75t_R g9909 ( 
.A(n_9506),
.Y(n_9909)
);

BUFx2_ASAP7_75t_L g9910 ( 
.A(n_9578),
.Y(n_9910)
);

INVx1_ASAP7_75t_L g9911 ( 
.A(n_9547),
.Y(n_9911)
);

BUFx3_ASAP7_75t_L g9912 ( 
.A(n_9609),
.Y(n_9912)
);

OAI22xp5_ASAP7_75t_L g9913 ( 
.A1(n_9849),
.A2(n_9287),
.B1(n_9107),
.B2(n_9113),
.Y(n_9913)
);

INVx3_ASAP7_75t_L g9914 ( 
.A(n_9571),
.Y(n_9914)
);

AND2x2_ASAP7_75t_L g9915 ( 
.A(n_9517),
.B(n_9368),
.Y(n_9915)
);

INVx6_ASAP7_75t_L g9916 ( 
.A(n_9641),
.Y(n_9916)
);

INVxp67_ASAP7_75t_SL g9917 ( 
.A(n_9558),
.Y(n_9917)
);

OAI22xp5_ASAP7_75t_L g9918 ( 
.A1(n_9767),
.A2(n_9342),
.B1(n_9291),
.B2(n_9297),
.Y(n_9918)
);

BUFx2_ASAP7_75t_SL g9919 ( 
.A(n_9723),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_9552),
.Y(n_9920)
);

BUFx12f_ASAP7_75t_L g9921 ( 
.A(n_9688),
.Y(n_9921)
);

OAI22xp33_ASAP7_75t_L g9922 ( 
.A1(n_9635),
.A2(n_9398),
.B1(n_9311),
.B2(n_9029),
.Y(n_9922)
);

BUFx6f_ASAP7_75t_L g9923 ( 
.A(n_9616),
.Y(n_9923)
);

INVx2_ASAP7_75t_L g9924 ( 
.A(n_9555),
.Y(n_9924)
);

AOI22xp33_ASAP7_75t_L g9925 ( 
.A1(n_9713),
.A2(n_9430),
.B1(n_9075),
.B2(n_9454),
.Y(n_9925)
);

INVx6_ASAP7_75t_L g9926 ( 
.A(n_9654),
.Y(n_9926)
);

INVx1_ASAP7_75t_SL g9927 ( 
.A(n_9817),
.Y(n_9927)
);

AOI22xp33_ASAP7_75t_L g9928 ( 
.A1(n_9802),
.A2(n_9464),
.B1(n_9402),
.B2(n_9426),
.Y(n_9928)
);

BUFx10_ASAP7_75t_L g9929 ( 
.A(n_9754),
.Y(n_9929)
);

NAND2xp5_ASAP7_75t_L g9930 ( 
.A(n_9781),
.B(n_9331),
.Y(n_9930)
);

INVx2_ASAP7_75t_SL g9931 ( 
.A(n_9769),
.Y(n_9931)
);

NAND2xp5_ASAP7_75t_L g9932 ( 
.A(n_9593),
.B(n_9486),
.Y(n_9932)
);

BUFx12f_ASAP7_75t_L g9933 ( 
.A(n_9749),
.Y(n_9933)
);

BUFx8_ASAP7_75t_L g9934 ( 
.A(n_9498),
.Y(n_9934)
);

INVx6_ASAP7_75t_L g9935 ( 
.A(n_9736),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_9563),
.Y(n_9936)
);

OAI22xp5_ASAP7_75t_L g9937 ( 
.A1(n_9755),
.A2(n_9260),
.B1(n_9461),
.B2(n_9457),
.Y(n_9937)
);

AOI22xp33_ASAP7_75t_L g9938 ( 
.A1(n_9618),
.A2(n_9572),
.B1(n_9620),
.B2(n_9622),
.Y(n_9938)
);

INVx2_ASAP7_75t_L g9939 ( 
.A(n_9577),
.Y(n_9939)
);

NAND2xp5_ASAP7_75t_L g9940 ( 
.A(n_9742),
.B(n_9438),
.Y(n_9940)
);

INVx3_ASAP7_75t_L g9941 ( 
.A(n_9836),
.Y(n_9941)
);

CKINVDCx20_ASAP7_75t_R g9942 ( 
.A(n_9613),
.Y(n_9942)
);

INVxp67_ASAP7_75t_SL g9943 ( 
.A(n_9587),
.Y(n_9943)
);

CKINVDCx11_ASAP7_75t_R g9944 ( 
.A(n_9846),
.Y(n_9944)
);

AOI22xp33_ASAP7_75t_SL g9945 ( 
.A1(n_9677),
.A2(n_9481),
.B1(n_9405),
.B2(n_9469),
.Y(n_9945)
);

INVx2_ASAP7_75t_L g9946 ( 
.A(n_9580),
.Y(n_9946)
);

AOI22xp33_ASAP7_75t_L g9947 ( 
.A1(n_9816),
.A2(n_9401),
.B1(n_9319),
.B2(n_9462),
.Y(n_9947)
);

AOI22xp33_ASAP7_75t_L g9948 ( 
.A1(n_9667),
.A2(n_9059),
.B1(n_9347),
.B2(n_9480),
.Y(n_9948)
);

INVx1_ASAP7_75t_L g9949 ( 
.A(n_9596),
.Y(n_9949)
);

INVx1_ASAP7_75t_L g9950 ( 
.A(n_9599),
.Y(n_9950)
);

INVx2_ASAP7_75t_L g9951 ( 
.A(n_9608),
.Y(n_9951)
);

AOI22xp33_ASAP7_75t_L g9952 ( 
.A1(n_9501),
.A2(n_9326),
.B1(n_9442),
.B2(n_9386),
.Y(n_9952)
);

NAND2x1p5_ASAP7_75t_L g9953 ( 
.A(n_9718),
.B(n_9263),
.Y(n_9953)
);

INVx11_ASAP7_75t_L g9954 ( 
.A(n_9779),
.Y(n_9954)
);

OAI22xp33_ASAP7_75t_L g9955 ( 
.A1(n_9718),
.A2(n_9418),
.B1(n_9377),
.B2(n_9149),
.Y(n_9955)
);

INVx2_ASAP7_75t_L g9956 ( 
.A(n_9617),
.Y(n_9956)
);

BUFx8_ASAP7_75t_L g9957 ( 
.A(n_9766),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_9637),
.Y(n_9958)
);

BUFx6f_ASAP7_75t_L g9959 ( 
.A(n_9616),
.Y(n_9959)
);

AOI22xp33_ASAP7_75t_L g9960 ( 
.A1(n_9606),
.A2(n_9386),
.B1(n_9351),
.B2(n_9116),
.Y(n_9960)
);

OAI22xp5_ASAP7_75t_L g9961 ( 
.A1(n_9775),
.A2(n_9207),
.B1(n_9259),
.B2(n_9240),
.Y(n_9961)
);

OAI22xp5_ASAP7_75t_L g9962 ( 
.A1(n_9872),
.A2(n_9355),
.B1(n_9361),
.B2(n_9410),
.Y(n_9962)
);

INVx1_ASAP7_75t_L g9963 ( 
.A(n_9639),
.Y(n_9963)
);

INVx2_ASAP7_75t_L g9964 ( 
.A(n_9649),
.Y(n_9964)
);

AOI22xp5_ASAP7_75t_L g9965 ( 
.A1(n_9527),
.A2(n_9070),
.B1(n_9237),
.B2(n_9230),
.Y(n_9965)
);

INVx2_ASAP7_75t_L g9966 ( 
.A(n_9655),
.Y(n_9966)
);

AOI22xp33_ASAP7_75t_L g9967 ( 
.A1(n_9528),
.A2(n_9247),
.B1(n_9277),
.B2(n_9302),
.Y(n_9967)
);

HB1xp67_ASAP7_75t_L g9968 ( 
.A(n_9499),
.Y(n_9968)
);

AOI22xp33_ASAP7_75t_L g9969 ( 
.A1(n_9750),
.A2(n_9488),
.B1(n_9491),
.B2(n_9266),
.Y(n_9969)
);

INVx2_ASAP7_75t_L g9970 ( 
.A(n_9658),
.Y(n_9970)
);

INVx1_ASAP7_75t_L g9971 ( 
.A(n_9666),
.Y(n_9971)
);

NAND2x1p5_ASAP7_75t_L g9972 ( 
.A(n_9600),
.B(n_9289),
.Y(n_9972)
);

CKINVDCx6p67_ASAP7_75t_R g9973 ( 
.A(n_9770),
.Y(n_9973)
);

AOI22xp5_ASAP7_75t_L g9974 ( 
.A1(n_9835),
.A2(n_9210),
.B1(n_9296),
.B2(n_9389),
.Y(n_9974)
);

OAI22xp5_ASAP7_75t_L g9975 ( 
.A1(n_9829),
.A2(n_9256),
.B1(n_9270),
.B2(n_9300),
.Y(n_9975)
);

INVx4_ASAP7_75t_L g9976 ( 
.A(n_9576),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_9721),
.Y(n_9977)
);

AOI22xp33_ASAP7_75t_L g9978 ( 
.A1(n_9674),
.A2(n_9339),
.B1(n_9340),
.B2(n_9330),
.Y(n_9978)
);

AOI22xp33_ASAP7_75t_L g9979 ( 
.A1(n_9694),
.A2(n_9417),
.B1(n_9379),
.B2(n_9279),
.Y(n_9979)
);

INVx1_ASAP7_75t_L g9980 ( 
.A(n_9760),
.Y(n_9980)
);

BUFx8_ASAP7_75t_L g9981 ( 
.A(n_9778),
.Y(n_9981)
);

BUFx12f_ASAP7_75t_L g9982 ( 
.A(n_9567),
.Y(n_9982)
);

BUFx2_ASAP7_75t_L g9983 ( 
.A(n_9632),
.Y(n_9983)
);

CKINVDCx11_ASAP7_75t_R g9984 ( 
.A(n_9565),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9511),
.Y(n_9985)
);

INVx1_ASAP7_75t_SL g9986 ( 
.A(n_9821),
.Y(n_9986)
);

BUFx2_ASAP7_75t_L g9987 ( 
.A(n_9797),
.Y(n_9987)
);

INVx6_ASAP7_75t_L g9988 ( 
.A(n_9804),
.Y(n_9988)
);

AOI22xp33_ASAP7_75t_L g9989 ( 
.A1(n_9537),
.A2(n_9406),
.B1(n_9453),
.B2(n_9440),
.Y(n_9989)
);

INVx1_ASAP7_75t_L g9990 ( 
.A(n_9515),
.Y(n_9990)
);

AOI22xp33_ASAP7_75t_L g9991 ( 
.A1(n_9861),
.A2(n_9086),
.B1(n_9357),
.B2(n_9328),
.Y(n_9991)
);

CKINVDCx11_ASAP7_75t_R g9992 ( 
.A(n_9565),
.Y(n_9992)
);

CKINVDCx20_ASAP7_75t_R g9993 ( 
.A(n_9759),
.Y(n_9993)
);

OAI22xp5_ASAP7_75t_L g9994 ( 
.A1(n_9627),
.A2(n_9314),
.B1(n_9286),
.B2(n_9334),
.Y(n_9994)
);

INVx3_ASAP7_75t_SL g9995 ( 
.A(n_9770),
.Y(n_9995)
);

INVx1_ASAP7_75t_L g9996 ( 
.A(n_9523),
.Y(n_9996)
);

OAI22xp5_ASAP7_75t_L g9997 ( 
.A1(n_9757),
.A2(n_1048),
.B1(n_1046),
.B2(n_1047),
.Y(n_9997)
);

BUFx12f_ASAP7_75t_L g9998 ( 
.A(n_9788),
.Y(n_9998)
);

INVx1_ASAP7_75t_L g9999 ( 
.A(n_9689),
.Y(n_9999)
);

AOI22xp5_ASAP7_75t_L g10000 ( 
.A1(n_9835),
.A2(n_1048),
.B1(n_1046),
.B2(n_1047),
.Y(n_10000)
);

AOI22xp33_ASAP7_75t_L g10001 ( 
.A1(n_9712),
.A2(n_1051),
.B1(n_1049),
.B2(n_1050),
.Y(n_10001)
);

NAND2xp5_ASAP7_75t_L g10002 ( 
.A(n_9607),
.B(n_9636),
.Y(n_10002)
);

INVx6_ASAP7_75t_L g10003 ( 
.A(n_9590),
.Y(n_10003)
);

CKINVDCx6p67_ASAP7_75t_R g10004 ( 
.A(n_9642),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_9692),
.Y(n_10005)
);

CKINVDCx11_ASAP7_75t_R g10006 ( 
.A(n_9590),
.Y(n_10006)
);

INVx6_ASAP7_75t_L g10007 ( 
.A(n_9603),
.Y(n_10007)
);

INVx1_ASAP7_75t_L g10008 ( 
.A(n_9699),
.Y(n_10008)
);

INVx6_ASAP7_75t_L g10009 ( 
.A(n_9603),
.Y(n_10009)
);

INVx1_ASAP7_75t_L g10010 ( 
.A(n_9521),
.Y(n_10010)
);

BUFx3_ASAP7_75t_L g10011 ( 
.A(n_9615),
.Y(n_10011)
);

INVx2_ASAP7_75t_L g10012 ( 
.A(n_9676),
.Y(n_10012)
);

AOI22xp33_ASAP7_75t_L g10013 ( 
.A1(n_9679),
.A2(n_1055),
.B1(n_1052),
.B2(n_1054),
.Y(n_10013)
);

INVx2_ASAP7_75t_L g10014 ( 
.A(n_9525),
.Y(n_10014)
);

INVx1_ASAP7_75t_L g10015 ( 
.A(n_9532),
.Y(n_10015)
);

INVx2_ASAP7_75t_SL g10016 ( 
.A(n_9624),
.Y(n_10016)
);

HB1xp67_ASAP7_75t_L g10017 ( 
.A(n_9531),
.Y(n_10017)
);

AOI22xp5_ASAP7_75t_SL g10018 ( 
.A1(n_9856),
.A2(n_1055),
.B1(n_1052),
.B2(n_1054),
.Y(n_10018)
);

OAI22xp5_ASAP7_75t_L g10019 ( 
.A1(n_9646),
.A2(n_1058),
.B1(n_1056),
.B2(n_1057),
.Y(n_10019)
);

INVx11_ASAP7_75t_L g10020 ( 
.A(n_9560),
.Y(n_10020)
);

AOI22xp33_ASAP7_75t_SL g10021 ( 
.A1(n_9835),
.A2(n_1058),
.B1(n_1056),
.B2(n_1057),
.Y(n_10021)
);

CKINVDCx20_ASAP7_75t_R g10022 ( 
.A(n_9732),
.Y(n_10022)
);

INVx1_ASAP7_75t_SL g10023 ( 
.A(n_9538),
.Y(n_10023)
);

CKINVDCx11_ASAP7_75t_R g10024 ( 
.A(n_9604),
.Y(n_10024)
);

AND2x2_ASAP7_75t_L g10025 ( 
.A(n_9656),
.B(n_1059),
.Y(n_10025)
);

INVx1_ASAP7_75t_L g10026 ( 
.A(n_9539),
.Y(n_10026)
);

AOI22xp33_ASAP7_75t_L g10027 ( 
.A1(n_9866),
.A2(n_1061),
.B1(n_1059),
.B2(n_1060),
.Y(n_10027)
);

AOI22xp5_ASAP7_75t_L g10028 ( 
.A1(n_9643),
.A2(n_1062),
.B1(n_1060),
.B2(n_1061),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_9540),
.Y(n_10029)
);

AOI22xp33_ASAP7_75t_SL g10030 ( 
.A1(n_9594),
.A2(n_9543),
.B1(n_9657),
.B2(n_9815),
.Y(n_10030)
);

AOI22xp33_ASAP7_75t_SL g10031 ( 
.A1(n_9514),
.A2(n_9500),
.B1(n_9623),
.B2(n_9873),
.Y(n_10031)
);

AND2x2_ASAP7_75t_L g10032 ( 
.A(n_9708),
.B(n_1062),
.Y(n_10032)
);

OAI22xp33_ASAP7_75t_L g10033 ( 
.A1(n_9651),
.A2(n_1065),
.B1(n_1063),
.B2(n_1064),
.Y(n_10033)
);

INVx2_ASAP7_75t_L g10034 ( 
.A(n_9544),
.Y(n_10034)
);

INVx2_ASAP7_75t_SL g10035 ( 
.A(n_9559),
.Y(n_10035)
);

INVx1_ASAP7_75t_L g10036 ( 
.A(n_9554),
.Y(n_10036)
);

OAI21xp5_ASAP7_75t_SL g10037 ( 
.A1(n_9811),
.A2(n_1063),
.B(n_1064),
.Y(n_10037)
);

INVx6_ASAP7_75t_L g10038 ( 
.A(n_9604),
.Y(n_10038)
);

INVx3_ASAP7_75t_L g10039 ( 
.A(n_9505),
.Y(n_10039)
);

OAI22xp5_ASAP7_75t_L g10040 ( 
.A1(n_9720),
.A2(n_1067),
.B1(n_1065),
.B2(n_1066),
.Y(n_10040)
);

NAND2xp5_ASAP7_75t_L g10041 ( 
.A(n_9799),
.B(n_1066),
.Y(n_10041)
);

INVx1_ASAP7_75t_L g10042 ( 
.A(n_9557),
.Y(n_10042)
);

OAI22xp33_ASAP7_75t_L g10043 ( 
.A1(n_9822),
.A2(n_1069),
.B1(n_1067),
.B2(n_1068),
.Y(n_10043)
);

CKINVDCx5p33_ASAP7_75t_R g10044 ( 
.A(n_9546),
.Y(n_10044)
);

BUFx10_ASAP7_75t_L g10045 ( 
.A(n_9874),
.Y(n_10045)
);

INVx4_ASAP7_75t_L g10046 ( 
.A(n_9700),
.Y(n_10046)
);

INVx2_ASAP7_75t_L g10047 ( 
.A(n_9582),
.Y(n_10047)
);

INVx1_ASAP7_75t_L g10048 ( 
.A(n_9588),
.Y(n_10048)
);

INVx1_ASAP7_75t_L g10049 ( 
.A(n_9585),
.Y(n_10049)
);

CKINVDCx20_ASAP7_75t_R g10050 ( 
.A(n_9854),
.Y(n_10050)
);

INVx1_ASAP7_75t_SL g10051 ( 
.A(n_9553),
.Y(n_10051)
);

BUFx2_ASAP7_75t_L g10052 ( 
.A(n_9813),
.Y(n_10052)
);

INVx2_ASAP7_75t_L g10053 ( 
.A(n_9703),
.Y(n_10053)
);

BUFx8_ASAP7_75t_L g10054 ( 
.A(n_9791),
.Y(n_10054)
);

BUFx4_ASAP7_75t_R g10055 ( 
.A(n_9848),
.Y(n_10055)
);

INVx2_ASAP7_75t_L g10056 ( 
.A(n_9710),
.Y(n_10056)
);

BUFx2_ASAP7_75t_L g10057 ( 
.A(n_9731),
.Y(n_10057)
);

INVx1_ASAP7_75t_SL g10058 ( 
.A(n_9711),
.Y(n_10058)
);

INVx3_ASAP7_75t_L g10059 ( 
.A(n_9512),
.Y(n_10059)
);

AND2x2_ASAP7_75t_L g10060 ( 
.A(n_9570),
.B(n_1070),
.Y(n_10060)
);

OAI22xp33_ASAP7_75t_L g10061 ( 
.A1(n_9630),
.A2(n_1073),
.B1(n_1071),
.B2(n_1072),
.Y(n_10061)
);

CKINVDCx6p67_ASAP7_75t_R g10062 ( 
.A(n_9870),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_9715),
.Y(n_10063)
);

INVx3_ASAP7_75t_L g10064 ( 
.A(n_9516),
.Y(n_10064)
);

INVx1_ASAP7_75t_L g10065 ( 
.A(n_9669),
.Y(n_10065)
);

INVx3_ASAP7_75t_L g10066 ( 
.A(n_9564),
.Y(n_10066)
);

BUFx2_ASAP7_75t_L g10067 ( 
.A(n_9868),
.Y(n_10067)
);

INVx2_ASAP7_75t_SL g10068 ( 
.A(n_9519),
.Y(n_10068)
);

INVx6_ASAP7_75t_L g10069 ( 
.A(n_9546),
.Y(n_10069)
);

CKINVDCx11_ASAP7_75t_R g10070 ( 
.A(n_9850),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_9803),
.Y(n_10071)
);

CKINVDCx20_ASAP7_75t_R g10072 ( 
.A(n_9782),
.Y(n_10072)
);

AOI22xp33_ASAP7_75t_L g10073 ( 
.A1(n_9860),
.A2(n_9566),
.B1(n_9837),
.B2(n_9839),
.Y(n_10073)
);

AOI22xp33_ASAP7_75t_L g10074 ( 
.A1(n_9497),
.A2(n_1075),
.B1(n_1071),
.B2(n_1072),
.Y(n_10074)
);

OAI22xp5_ASAP7_75t_L g10075 ( 
.A1(n_9773),
.A2(n_1077),
.B1(n_1075),
.B2(n_1076),
.Y(n_10075)
);

AOI22xp33_ASAP7_75t_L g10076 ( 
.A1(n_9535),
.A2(n_1079),
.B1(n_1076),
.B2(n_1078),
.Y(n_10076)
);

OAI22xp33_ASAP7_75t_L g10077 ( 
.A1(n_9568),
.A2(n_1080),
.B1(n_1078),
.B2(n_1079),
.Y(n_10077)
);

OAI22xp5_ASAP7_75t_L g10078 ( 
.A1(n_9855),
.A2(n_1082),
.B1(n_1080),
.B2(n_1081),
.Y(n_10078)
);

CKINVDCx6p67_ASAP7_75t_R g10079 ( 
.A(n_9870),
.Y(n_10079)
);

BUFx3_ASAP7_75t_L g10080 ( 
.A(n_9850),
.Y(n_10080)
);

INVx1_ASAP7_75t_L g10081 ( 
.A(n_9729),
.Y(n_10081)
);

BUFx8_ASAP7_75t_L g10082 ( 
.A(n_9824),
.Y(n_10082)
);

INVx5_ASAP7_75t_L g10083 ( 
.A(n_9869),
.Y(n_10083)
);

CKINVDCx5p33_ASAP7_75t_R g10084 ( 
.A(n_9562),
.Y(n_10084)
);

OAI22xp33_ASAP7_75t_L g10085 ( 
.A1(n_9534),
.A2(n_1084),
.B1(n_1081),
.B2(n_1083),
.Y(n_10085)
);

CKINVDCx5p33_ASAP7_75t_R g10086 ( 
.A(n_9562),
.Y(n_10086)
);

INVx6_ASAP7_75t_L g10087 ( 
.A(n_9700),
.Y(n_10087)
);

INVx1_ASAP7_75t_L g10088 ( 
.A(n_9716),
.Y(n_10088)
);

INVx1_ASAP7_75t_L g10089 ( 
.A(n_9730),
.Y(n_10089)
);

BUFx2_ASAP7_75t_L g10090 ( 
.A(n_9768),
.Y(n_10090)
);

AOI22xp33_ASAP7_75t_L g10091 ( 
.A1(n_9660),
.A2(n_1085),
.B1(n_1083),
.B2(n_1084),
.Y(n_10091)
);

AOI22xp33_ASAP7_75t_L g10092 ( 
.A1(n_9704),
.A2(n_1088),
.B1(n_1086),
.B2(n_1087),
.Y(n_10092)
);

CKINVDCx11_ASAP7_75t_R g10093 ( 
.A(n_9869),
.Y(n_10093)
);

AOI22xp33_ASAP7_75t_L g10094 ( 
.A1(n_9549),
.A2(n_1091),
.B1(n_1086),
.B2(n_1088),
.Y(n_10094)
);

BUFx8_ASAP7_75t_SL g10095 ( 
.A(n_9589),
.Y(n_10095)
);

INVx1_ASAP7_75t_L g10096 ( 
.A(n_9758),
.Y(n_10096)
);

OAI22xp33_ASAP7_75t_L g10097 ( 
.A1(n_9534),
.A2(n_1093),
.B1(n_1091),
.B2(n_1092),
.Y(n_10097)
);

CKINVDCx11_ASAP7_75t_R g10098 ( 
.A(n_9733),
.Y(n_10098)
);

BUFx3_ASAP7_75t_L g10099 ( 
.A(n_9653),
.Y(n_10099)
);

INVx1_ASAP7_75t_L g10100 ( 
.A(n_9698),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_9786),
.Y(n_10101)
);

AOI22xp5_ASAP7_75t_L g10102 ( 
.A1(n_9503),
.A2(n_1095),
.B1(n_1092),
.B2(n_1094),
.Y(n_10102)
);

INVx1_ASAP7_75t_L g10103 ( 
.A(n_9753),
.Y(n_10103)
);

CKINVDCx11_ASAP7_75t_R g10104 ( 
.A(n_9733),
.Y(n_10104)
);

INVx1_ASAP7_75t_L g10105 ( 
.A(n_9784),
.Y(n_10105)
);

BUFx4f_ASAP7_75t_L g10106 ( 
.A(n_9682),
.Y(n_10106)
);

INVx1_ASAP7_75t_L g10107 ( 
.A(n_9820),
.Y(n_10107)
);

BUFx10_ASAP7_75t_L g10108 ( 
.A(n_9780),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_9831),
.Y(n_10109)
);

NAND2xp5_ASAP7_75t_L g10110 ( 
.A(n_9798),
.B(n_1094),
.Y(n_10110)
);

BUFx3_ASAP7_75t_L g10111 ( 
.A(n_9681),
.Y(n_10111)
);

OAI22xp5_ASAP7_75t_L g10112 ( 
.A1(n_9725),
.A2(n_1100),
.B1(n_1097),
.B2(n_1098),
.Y(n_10112)
);

BUFx8_ASAP7_75t_SL g10113 ( 
.A(n_9601),
.Y(n_10113)
);

BUFx12f_ASAP7_75t_L g10114 ( 
.A(n_9851),
.Y(n_10114)
);

AO22x1_ASAP7_75t_L g10115 ( 
.A1(n_9541),
.A2(n_9586),
.B1(n_9659),
.B2(n_9808),
.Y(n_10115)
);

AOI22xp33_ASAP7_75t_L g10116 ( 
.A1(n_9518),
.A2(n_1102),
.B1(n_1100),
.B2(n_1101),
.Y(n_10116)
);

BUFx4f_ASAP7_75t_SL g10117 ( 
.A(n_9561),
.Y(n_10117)
);

AOI22xp5_ASAP7_75t_L g10118 ( 
.A1(n_9520),
.A2(n_1103),
.B1(n_1101),
.B2(n_1102),
.Y(n_10118)
);

AOI22xp33_ASAP7_75t_SL g10119 ( 
.A1(n_9665),
.A2(n_1105),
.B1(n_1103),
.B2(n_1104),
.Y(n_10119)
);

INVx2_ASAP7_75t_SL g10120 ( 
.A(n_9792),
.Y(n_10120)
);

INVx6_ASAP7_75t_L g10121 ( 
.A(n_9793),
.Y(n_10121)
);

BUFx12f_ASAP7_75t_L g10122 ( 
.A(n_9765),
.Y(n_10122)
);

AOI22xp33_ASAP7_75t_L g10123 ( 
.A1(n_9592),
.A2(n_9574),
.B1(n_9734),
.B2(n_9748),
.Y(n_10123)
);

AOI22xp33_ASAP7_75t_SL g10124 ( 
.A1(n_9504),
.A2(n_1106),
.B1(n_1104),
.B2(n_1105),
.Y(n_10124)
);

CKINVDCx5p33_ASAP7_75t_R g10125 ( 
.A(n_9629),
.Y(n_10125)
);

OAI22xp33_ASAP7_75t_L g10126 ( 
.A1(n_9631),
.A2(n_1108),
.B1(n_1106),
.B2(n_1107),
.Y(n_10126)
);

BUFx6f_ASAP7_75t_L g10127 ( 
.A(n_9633),
.Y(n_10127)
);

AOI22xp33_ASAP7_75t_L g10128 ( 
.A1(n_9722),
.A2(n_1109),
.B1(n_1107),
.B2(n_1108),
.Y(n_10128)
);

AOI22xp5_ASAP7_75t_SL g10129 ( 
.A1(n_9828),
.A2(n_1111),
.B1(n_1109),
.B2(n_1110),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_9845),
.Y(n_10130)
);

INVx1_ASAP7_75t_L g10131 ( 
.A(n_9853),
.Y(n_10131)
);

INVx6_ASAP7_75t_L g10132 ( 
.A(n_9787),
.Y(n_10132)
);

AOI22xp33_ASAP7_75t_L g10133 ( 
.A1(n_9598),
.A2(n_1113),
.B1(n_1110),
.B2(n_1112),
.Y(n_10133)
);

OAI22xp5_ASAP7_75t_L g10134 ( 
.A1(n_9867),
.A2(n_1115),
.B1(n_1113),
.B2(n_1114),
.Y(n_10134)
);

INVx1_ASAP7_75t_L g10135 ( 
.A(n_9862),
.Y(n_10135)
);

INVx1_ASAP7_75t_L g10136 ( 
.A(n_9871),
.Y(n_10136)
);

INVx1_ASAP7_75t_L g10137 ( 
.A(n_9510),
.Y(n_10137)
);

BUFx3_ASAP7_75t_L g10138 ( 
.A(n_9774),
.Y(n_10138)
);

NAND2xp5_ASAP7_75t_L g10139 ( 
.A(n_9805),
.B(n_1114),
.Y(n_10139)
);

AOI22xp5_ASAP7_75t_L g10140 ( 
.A1(n_9550),
.A2(n_1117),
.B1(n_1115),
.B2(n_1116),
.Y(n_10140)
);

CKINVDCx11_ASAP7_75t_R g10141 ( 
.A(n_9843),
.Y(n_10141)
);

INVx2_ASAP7_75t_L g10142 ( 
.A(n_9744),
.Y(n_10142)
);

AOI22xp33_ASAP7_75t_L g10143 ( 
.A1(n_9823),
.A2(n_1119),
.B1(n_1116),
.B2(n_1118),
.Y(n_10143)
);

INVx6_ASAP7_75t_L g10144 ( 
.A(n_9695),
.Y(n_10144)
);

BUFx6f_ASAP7_75t_L g10145 ( 
.A(n_9644),
.Y(n_10145)
);

AOI22xp33_ASAP7_75t_L g10146 ( 
.A1(n_9847),
.A2(n_1120),
.B1(n_1118),
.B2(n_1119),
.Y(n_10146)
);

BUFx3_ASAP7_75t_L g10147 ( 
.A(n_9579),
.Y(n_10147)
);

INVx1_ASAP7_75t_L g10148 ( 
.A(n_9533),
.Y(n_10148)
);

AOI22xp33_ASAP7_75t_L g10149 ( 
.A1(n_9583),
.A2(n_1123),
.B1(n_1121),
.B2(n_1122),
.Y(n_10149)
);

INVx2_ASAP7_75t_L g10150 ( 
.A(n_9827),
.Y(n_10150)
);

OAI22xp33_ASAP7_75t_SL g10151 ( 
.A1(n_9648),
.A2(n_1123),
.B1(n_1121),
.B2(n_1122),
.Y(n_10151)
);

OAI22xp33_ASAP7_75t_L g10152 ( 
.A1(n_9645),
.A2(n_1126),
.B1(n_1124),
.B2(n_1125),
.Y(n_10152)
);

NAND2xp5_ASAP7_75t_L g10153 ( 
.A(n_9807),
.B(n_1125),
.Y(n_10153)
);

INVx1_ASAP7_75t_L g10154 ( 
.A(n_9551),
.Y(n_10154)
);

BUFx4f_ASAP7_75t_SL g10155 ( 
.A(n_9664),
.Y(n_10155)
);

INVx1_ASAP7_75t_SL g10156 ( 
.A(n_9746),
.Y(n_10156)
);

INVx2_ASAP7_75t_SL g10157 ( 
.A(n_9686),
.Y(n_10157)
);

AND2x2_ASAP7_75t_L g10158 ( 
.A(n_9584),
.B(n_1126),
.Y(n_10158)
);

BUFx2_ASAP7_75t_L g10159 ( 
.A(n_9735),
.Y(n_10159)
);

AOI22xp33_ASAP7_75t_SL g10160 ( 
.A1(n_9595),
.A2(n_1129),
.B1(n_1127),
.B2(n_1128),
.Y(n_10160)
);

INVx1_ASAP7_75t_L g10161 ( 
.A(n_9671),
.Y(n_10161)
);

CKINVDCx6p67_ASAP7_75t_R g10162 ( 
.A(n_9785),
.Y(n_10162)
);

INVx2_ASAP7_75t_L g10163 ( 
.A(n_9834),
.Y(n_10163)
);

INVx1_ASAP7_75t_SL g10164 ( 
.A(n_9858),
.Y(n_10164)
);

BUFx6f_ASAP7_75t_SL g10165 ( 
.A(n_9696),
.Y(n_10165)
);

OAI22xp33_ASAP7_75t_L g10166 ( 
.A1(n_9526),
.A2(n_1129),
.B1(n_1127),
.B2(n_1128),
.Y(n_10166)
);

CKINVDCx16_ASAP7_75t_R g10167 ( 
.A(n_9812),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_9529),
.Y(n_10168)
);

AOI22xp33_ASAP7_75t_SL g10169 ( 
.A1(n_9575),
.A2(n_1132),
.B1(n_1130),
.B2(n_1131),
.Y(n_10169)
);

INVx2_ASAP7_75t_SL g10170 ( 
.A(n_9859),
.Y(n_10170)
);

BUFx12f_ASAP7_75t_L g10171 ( 
.A(n_9777),
.Y(n_10171)
);

OAI22xp5_ASAP7_75t_L g10172 ( 
.A1(n_9591),
.A2(n_1132),
.B1(n_1130),
.B2(n_1131),
.Y(n_10172)
);

INVx1_ASAP7_75t_L g10173 ( 
.A(n_9597),
.Y(n_10173)
);

BUFx3_ASAP7_75t_L g10174 ( 
.A(n_9739),
.Y(n_10174)
);

BUFx6f_ASAP7_75t_L g10175 ( 
.A(n_9581),
.Y(n_10175)
);

AOI22xp33_ASAP7_75t_L g10176 ( 
.A1(n_9610),
.A2(n_1136),
.B1(n_1133),
.B2(n_1134),
.Y(n_10176)
);

CKINVDCx20_ASAP7_75t_R g10177 ( 
.A(n_9717),
.Y(n_10177)
);

INVx4_ASAP7_75t_L g10178 ( 
.A(n_9844),
.Y(n_10178)
);

INVx1_ASAP7_75t_L g10179 ( 
.A(n_9795),
.Y(n_10179)
);

INVx1_ASAP7_75t_SL g10180 ( 
.A(n_9841),
.Y(n_10180)
);

AOI22xp33_ASAP7_75t_L g10181 ( 
.A1(n_9508),
.A2(n_1137),
.B1(n_1134),
.B2(n_1136),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_9977),
.Y(n_10182)
);

INVx1_ASAP7_75t_L g10183 ( 
.A(n_9875),
.Y(n_10183)
);

BUFx2_ASAP7_75t_R g10184 ( 
.A(n_9919),
.Y(n_10184)
);

INVx2_ASAP7_75t_L g10185 ( 
.A(n_9890),
.Y(n_10185)
);

OAI22xp5_ASAP7_75t_L g10186 ( 
.A1(n_9938),
.A2(n_9628),
.B1(n_9796),
.B2(n_9789),
.Y(n_10186)
);

HB1xp67_ASAP7_75t_L g10187 ( 
.A(n_9968),
.Y(n_10187)
);

BUFx2_ASAP7_75t_L g10188 ( 
.A(n_9908),
.Y(n_10188)
);

INVx2_ASAP7_75t_L g10189 ( 
.A(n_9924),
.Y(n_10189)
);

HB1xp67_ASAP7_75t_L g10190 ( 
.A(n_10173),
.Y(n_10190)
);

AND2x2_ASAP7_75t_L g10191 ( 
.A(n_10167),
.B(n_9810),
.Y(n_10191)
);

AOI21x1_ASAP7_75t_L g10192 ( 
.A1(n_10115),
.A2(n_9670),
.B(n_9719),
.Y(n_10192)
);

BUFx3_ASAP7_75t_L g10193 ( 
.A(n_9934),
.Y(n_10193)
);

BUFx2_ASAP7_75t_L g10194 ( 
.A(n_10004),
.Y(n_10194)
);

AND2x2_ASAP7_75t_L g10195 ( 
.A(n_10067),
.B(n_9800),
.Y(n_10195)
);

INVxp67_ASAP7_75t_L g10196 ( 
.A(n_10137),
.Y(n_10196)
);

INVx2_ASAP7_75t_L g10197 ( 
.A(n_9939),
.Y(n_10197)
);

OAI21x1_ASAP7_75t_L g10198 ( 
.A1(n_10088),
.A2(n_9556),
.B(n_9545),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_L g10199 ( 
.A(n_10148),
.B(n_9522),
.Y(n_10199)
);

INVx1_ASAP7_75t_L g10200 ( 
.A(n_9980),
.Y(n_10200)
);

OAI21x1_ASAP7_75t_L g10201 ( 
.A1(n_10154),
.A2(n_9602),
.B(n_9761),
.Y(n_10201)
);

AO21x1_ASAP7_75t_SL g10202 ( 
.A1(n_9877),
.A2(n_9614),
.B(n_9707),
.Y(n_10202)
);

INVx1_ASAP7_75t_L g10203 ( 
.A(n_9898),
.Y(n_10203)
);

HB1xp67_ASAP7_75t_L g10204 ( 
.A(n_9943),
.Y(n_10204)
);

INVx1_ASAP7_75t_SL g10205 ( 
.A(n_10055),
.Y(n_10205)
);

HB1xp67_ASAP7_75t_L g10206 ( 
.A(n_9917),
.Y(n_10206)
);

AOI21x1_ASAP7_75t_L g10207 ( 
.A1(n_9891),
.A2(n_9687),
.B(n_9680),
.Y(n_10207)
);

INVx2_ASAP7_75t_L g10208 ( 
.A(n_9946),
.Y(n_10208)
);

INVx2_ASAP7_75t_L g10209 ( 
.A(n_9951),
.Y(n_10209)
);

INVx2_ASAP7_75t_L g10210 ( 
.A(n_9956),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_9958),
.Y(n_10211)
);

BUFx2_ASAP7_75t_SL g10212 ( 
.A(n_10022),
.Y(n_10212)
);

INVx2_ASAP7_75t_L g10213 ( 
.A(n_9964),
.Y(n_10213)
);

INVx6_ASAP7_75t_L g10214 ( 
.A(n_9896),
.Y(n_10214)
);

INVx2_ASAP7_75t_L g10215 ( 
.A(n_9966),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9900),
.Y(n_10216)
);

BUFx6f_ASAP7_75t_L g10217 ( 
.A(n_10093),
.Y(n_10217)
);

HB1xp67_ASAP7_75t_L g10218 ( 
.A(n_10065),
.Y(n_10218)
);

OA21x2_ASAP7_75t_L g10219 ( 
.A1(n_9910),
.A2(n_9697),
.B(n_9706),
.Y(n_10219)
);

AND2x2_ASAP7_75t_L g10220 ( 
.A(n_9987),
.B(n_9832),
.Y(n_10220)
);

AOI21x1_ASAP7_75t_L g10221 ( 
.A1(n_10110),
.A2(n_10153),
.B(n_10139),
.Y(n_10221)
);

INVx11_ASAP7_75t_L g10222 ( 
.A(n_9982),
.Y(n_10222)
);

INVx2_ASAP7_75t_SL g10223 ( 
.A(n_9988),
.Y(n_10223)
);

AND2x2_ASAP7_75t_L g10224 ( 
.A(n_10052),
.B(n_9983),
.Y(n_10224)
);

INVx1_ASAP7_75t_L g10225 ( 
.A(n_9903),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_9911),
.Y(n_10226)
);

OR2x2_ASAP7_75t_L g10227 ( 
.A(n_10168),
.B(n_9857),
.Y(n_10227)
);

BUFx2_ASAP7_75t_L g10228 ( 
.A(n_9878),
.Y(n_10228)
);

INVx2_ASAP7_75t_L g10229 ( 
.A(n_9970),
.Y(n_10229)
);

OAI21xp5_ASAP7_75t_L g10230 ( 
.A1(n_10031),
.A2(n_9619),
.B(n_9693),
.Y(n_10230)
);

INVx1_ASAP7_75t_L g10231 ( 
.A(n_9920),
.Y(n_10231)
);

AOI22xp33_ASAP7_75t_SL g10232 ( 
.A1(n_9884),
.A2(n_9776),
.B1(n_9684),
.B2(n_9740),
.Y(n_10232)
);

AOI22xp33_ASAP7_75t_L g10233 ( 
.A1(n_10030),
.A2(n_9882),
.B1(n_9876),
.B2(n_10033),
.Y(n_10233)
);

BUFx2_ASAP7_75t_L g10234 ( 
.A(n_9953),
.Y(n_10234)
);

AND2x4_ASAP7_75t_L g10235 ( 
.A(n_9914),
.B(n_9833),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9936),
.Y(n_10236)
);

INVx1_ASAP7_75t_L g10237 ( 
.A(n_9949),
.Y(n_10237)
);

INVx2_ASAP7_75t_L g10238 ( 
.A(n_10057),
.Y(n_10238)
);

INVx2_ASAP7_75t_L g10239 ( 
.A(n_10053),
.Y(n_10239)
);

INVx1_ASAP7_75t_L g10240 ( 
.A(n_9950),
.Y(n_10240)
);

INVx2_ASAP7_75t_L g10241 ( 
.A(n_10056),
.Y(n_10241)
);

BUFx3_ASAP7_75t_L g10242 ( 
.A(n_10095),
.Y(n_10242)
);

OA21x2_ASAP7_75t_L g10243 ( 
.A1(n_9930),
.A2(n_9678),
.B(n_9728),
.Y(n_10243)
);

CKINVDCx11_ASAP7_75t_R g10244 ( 
.A(n_9944),
.Y(n_10244)
);

HB1xp67_ASAP7_75t_L g10245 ( 
.A(n_10017),
.Y(n_10245)
);

CKINVDCx6p67_ASAP7_75t_R g10246 ( 
.A(n_10083),
.Y(n_10246)
);

INVx1_ASAP7_75t_L g10247 ( 
.A(n_9963),
.Y(n_10247)
);

INVx2_ASAP7_75t_L g10248 ( 
.A(n_10096),
.Y(n_10248)
);

INVx2_ASAP7_75t_L g10249 ( 
.A(n_10103),
.Y(n_10249)
);

INVx1_ASAP7_75t_L g10250 ( 
.A(n_9971),
.Y(n_10250)
);

OA21x2_ASAP7_75t_L g10251 ( 
.A1(n_10063),
.A2(n_9709),
.B(n_9727),
.Y(n_10251)
);

INVx1_ASAP7_75t_L g10252 ( 
.A(n_9999),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_10005),
.Y(n_10253)
);

INVx2_ASAP7_75t_L g10254 ( 
.A(n_9892),
.Y(n_10254)
);

INVx2_ASAP7_75t_L g10255 ( 
.A(n_9897),
.Y(n_10255)
);

INVx2_ASAP7_75t_L g10256 ( 
.A(n_9899),
.Y(n_10256)
);

INVx2_ASAP7_75t_SL g10257 ( 
.A(n_9988),
.Y(n_10257)
);

AO21x2_ASAP7_75t_L g10258 ( 
.A1(n_9901),
.A2(n_9772),
.B(n_9741),
.Y(n_10258)
);

INVx3_ASAP7_75t_L g10259 ( 
.A(n_9916),
.Y(n_10259)
);

INVx3_ASAP7_75t_L g10260 ( 
.A(n_9916),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_10081),
.Y(n_10261)
);

INVx2_ASAP7_75t_L g10262 ( 
.A(n_9904),
.Y(n_10262)
);

AND2x2_ASAP7_75t_L g10263 ( 
.A(n_10058),
.B(n_9864),
.Y(n_10263)
);

INVx2_ASAP7_75t_L g10264 ( 
.A(n_10014),
.Y(n_10264)
);

BUFx2_ASAP7_75t_R g10265 ( 
.A(n_9912),
.Y(n_10265)
);

BUFx3_ASAP7_75t_L g10266 ( 
.A(n_10113),
.Y(n_10266)
);

INVx1_ASAP7_75t_L g10267 ( 
.A(n_10008),
.Y(n_10267)
);

INVx3_ASAP7_75t_L g10268 ( 
.A(n_9883),
.Y(n_10268)
);

INVx2_ASAP7_75t_L g10269 ( 
.A(n_10034),
.Y(n_10269)
);

INVx2_ASAP7_75t_SL g10270 ( 
.A(n_10020),
.Y(n_10270)
);

NAND2xp5_ASAP7_75t_SL g10271 ( 
.A(n_9889),
.B(n_10023),
.Y(n_10271)
);

AOI22xp33_ASAP7_75t_L g10272 ( 
.A1(n_9905),
.A2(n_9840),
.B1(n_9751),
.B2(n_9826),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_10107),
.Y(n_10273)
);

AOI221xp5_ASAP7_75t_L g10274 ( 
.A1(n_9894),
.A2(n_10061),
.B1(n_10126),
.B2(n_10077),
.C(n_10166),
.Y(n_10274)
);

INVxp67_ASAP7_75t_SL g10275 ( 
.A(n_10002),
.Y(n_10275)
);

AO21x2_ASAP7_75t_L g10276 ( 
.A1(n_10041),
.A2(n_9801),
.B(n_9818),
.Y(n_10276)
);

INVx1_ASAP7_75t_L g10277 ( 
.A(n_10109),
.Y(n_10277)
);

AND2x2_ASAP7_75t_L g10278 ( 
.A(n_10159),
.B(n_9814),
.Y(n_10278)
);

INVx2_ASAP7_75t_L g10279 ( 
.A(n_10047),
.Y(n_10279)
);

AND2x2_ASAP7_75t_L g10280 ( 
.A(n_9986),
.B(n_9747),
.Y(n_10280)
);

OAI21x1_ASAP7_75t_L g10281 ( 
.A1(n_10130),
.A2(n_9783),
.B(n_9726),
.Y(n_10281)
);

INVx1_ASAP7_75t_L g10282 ( 
.A(n_10131),
.Y(n_10282)
);

INVx2_ASAP7_75t_L g10283 ( 
.A(n_10135),
.Y(n_10283)
);

INVx2_ASAP7_75t_L g10284 ( 
.A(n_10136),
.Y(n_10284)
);

INVx2_ASAP7_75t_L g10285 ( 
.A(n_10090),
.Y(n_10285)
);

AND2x2_ASAP7_75t_L g10286 ( 
.A(n_9879),
.B(n_9762),
.Y(n_10286)
);

OAI21x1_ASAP7_75t_L g10287 ( 
.A1(n_10105),
.A2(n_9673),
.B(n_9764),
.Y(n_10287)
);

INVx2_ASAP7_75t_L g10288 ( 
.A(n_10179),
.Y(n_10288)
);

INVx2_ASAP7_75t_L g10289 ( 
.A(n_10010),
.Y(n_10289)
);

OR2x2_ASAP7_75t_L g10290 ( 
.A(n_10089),
.B(n_9737),
.Y(n_10290)
);

INVx2_ASAP7_75t_L g10291 ( 
.A(n_10015),
.Y(n_10291)
);

INVx4_ASAP7_75t_L g10292 ( 
.A(n_9906),
.Y(n_10292)
);

INVx3_ASAP7_75t_L g10293 ( 
.A(n_10178),
.Y(n_10293)
);

OAI22xp5_ASAP7_75t_L g10294 ( 
.A1(n_9887),
.A2(n_9863),
.B1(n_9690),
.B2(n_9701),
.Y(n_10294)
);

INVx2_ASAP7_75t_L g10295 ( 
.A(n_10026),
.Y(n_10295)
);

AOI22xp33_ASAP7_75t_L g10296 ( 
.A1(n_9885),
.A2(n_9842),
.B1(n_9819),
.B2(n_9626),
.Y(n_10296)
);

INVx1_ASAP7_75t_L g10297 ( 
.A(n_9985),
.Y(n_10297)
);

INVx1_ASAP7_75t_L g10298 ( 
.A(n_9990),
.Y(n_10298)
);

INVx1_ASAP7_75t_L g10299 ( 
.A(n_9996),
.Y(n_10299)
);

NAND2x1_ASAP7_75t_L g10300 ( 
.A(n_10100),
.B(n_9611),
.Y(n_10300)
);

INVx1_ASAP7_75t_L g10301 ( 
.A(n_10029),
.Y(n_10301)
);

INVx1_ASAP7_75t_L g10302 ( 
.A(n_10036),
.Y(n_10302)
);

AOI22xp33_ASAP7_75t_L g10303 ( 
.A1(n_10073),
.A2(n_9661),
.B1(n_9675),
.B2(n_9825),
.Y(n_10303)
);

BUFx6f_ASAP7_75t_L g10304 ( 
.A(n_9984),
.Y(n_10304)
);

BUFx6f_ASAP7_75t_L g10305 ( 
.A(n_9992),
.Y(n_10305)
);

INVx2_ASAP7_75t_L g10306 ( 
.A(n_10042),
.Y(n_10306)
);

INVx2_ASAP7_75t_SL g10307 ( 
.A(n_9902),
.Y(n_10307)
);

INVx2_ASAP7_75t_SL g10308 ( 
.A(n_9902),
.Y(n_10308)
);

INVx2_ASAP7_75t_L g10309 ( 
.A(n_10048),
.Y(n_10309)
);

INVx1_ASAP7_75t_L g10310 ( 
.A(n_10049),
.Y(n_10310)
);

INVx3_ASAP7_75t_L g10311 ( 
.A(n_9935),
.Y(n_10311)
);

INVx2_ASAP7_75t_L g10312 ( 
.A(n_10012),
.Y(n_10312)
);

INVx1_ASAP7_75t_SL g10313 ( 
.A(n_9993),
.Y(n_10313)
);

BUFx2_ASAP7_75t_L g10314 ( 
.A(n_10072),
.Y(n_10314)
);

INVx2_ASAP7_75t_SL g10315 ( 
.A(n_9935),
.Y(n_10315)
);

INVx3_ASAP7_75t_L g10316 ( 
.A(n_10175),
.Y(n_10316)
);

INVx3_ASAP7_75t_L g10317 ( 
.A(n_10175),
.Y(n_10317)
);

INVx1_ASAP7_75t_L g10318 ( 
.A(n_10101),
.Y(n_10318)
);

AND2x2_ASAP7_75t_L g10319 ( 
.A(n_9915),
.B(n_9685),
.Y(n_10319)
);

INVx1_ASAP7_75t_L g10320 ( 
.A(n_10071),
.Y(n_10320)
);

INVx1_ASAP7_75t_L g10321 ( 
.A(n_10161),
.Y(n_10321)
);

INVx4_ASAP7_75t_L g10322 ( 
.A(n_9954),
.Y(n_10322)
);

BUFx3_ASAP7_75t_L g10323 ( 
.A(n_9921),
.Y(n_10323)
);

CKINVDCx5p33_ASAP7_75t_R g10324 ( 
.A(n_9909),
.Y(n_10324)
);

AOI21x1_ASAP7_75t_L g10325 ( 
.A1(n_9975),
.A2(n_9994),
.B(n_10025),
.Y(n_10325)
);

INVx2_ASAP7_75t_L g10326 ( 
.A(n_10150),
.Y(n_10326)
);

INVx3_ASAP7_75t_L g10327 ( 
.A(n_10046),
.Y(n_10327)
);

INVx2_ASAP7_75t_L g10328 ( 
.A(n_10163),
.Y(n_10328)
);

INVx1_ASAP7_75t_SL g10329 ( 
.A(n_10006),
.Y(n_10329)
);

AND2x2_ASAP7_75t_L g10330 ( 
.A(n_10156),
.B(n_9647),
.Y(n_10330)
);

INVx2_ASAP7_75t_L g10331 ( 
.A(n_10142),
.Y(n_10331)
);

OA21x2_ASAP7_75t_L g10332 ( 
.A1(n_9989),
.A2(n_9752),
.B(n_9743),
.Y(n_10332)
);

INVx1_ASAP7_75t_L g10333 ( 
.A(n_10180),
.Y(n_10333)
);

OAI21x1_ASAP7_75t_L g10334 ( 
.A1(n_9941),
.A2(n_9852),
.B(n_9745),
.Y(n_10334)
);

OAI21x1_ASAP7_75t_L g10335 ( 
.A1(n_9972),
.A2(n_9838),
.B(n_9638),
.Y(n_10335)
);

INVx4_ASAP7_75t_L g10336 ( 
.A(n_10083),
.Y(n_10336)
);

CKINVDCx5p33_ASAP7_75t_R g10337 ( 
.A(n_9942),
.Y(n_10337)
);

AO21x1_ASAP7_75t_SL g10338 ( 
.A1(n_9952),
.A2(n_9809),
.B(n_9672),
.Y(n_10338)
);

INVx2_ASAP7_75t_L g10339 ( 
.A(n_10120),
.Y(n_10339)
);

OR2x2_ASAP7_75t_L g10340 ( 
.A(n_9932),
.B(n_9691),
.Y(n_10340)
);

OAI21x1_ASAP7_75t_L g10341 ( 
.A1(n_9893),
.A2(n_9705),
.B(n_9714),
.Y(n_10341)
);

OAI22xp5_ASAP7_75t_L g10342 ( 
.A1(n_9880),
.A2(n_9672),
.B1(n_9830),
.B2(n_9865),
.Y(n_10342)
);

INVx2_ASAP7_75t_SL g10343 ( 
.A(n_10108),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_10068),
.Y(n_10344)
);

HB1xp67_ASAP7_75t_L g10345 ( 
.A(n_10051),
.Y(n_10345)
);

OAI21x1_ASAP7_75t_L g10346 ( 
.A1(n_10039),
.A2(n_1137),
.B(n_1138),
.Y(n_10346)
);

AND2x2_ASAP7_75t_L g10347 ( 
.A(n_10035),
.B(n_1139),
.Y(n_10347)
);

INVx2_ASAP7_75t_L g10348 ( 
.A(n_10157),
.Y(n_10348)
);

HB1xp67_ASAP7_75t_L g10349 ( 
.A(n_9927),
.Y(n_10349)
);

HB1xp67_ASAP7_75t_L g10350 ( 
.A(n_10060),
.Y(n_10350)
);

INVx1_ASAP7_75t_L g10351 ( 
.A(n_9940),
.Y(n_10351)
);

INVx2_ASAP7_75t_L g10352 ( 
.A(n_10144),
.Y(n_10352)
);

INVx1_ASAP7_75t_L g10353 ( 
.A(n_10170),
.Y(n_10353)
);

INVx2_ASAP7_75t_SL g10354 ( 
.A(n_9926),
.Y(n_10354)
);

AO21x2_ASAP7_75t_L g10355 ( 
.A1(n_10085),
.A2(n_1139),
.B(n_1140),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_10164),
.Y(n_10356)
);

CKINVDCx5p33_ASAP7_75t_R g10357 ( 
.A(n_9933),
.Y(n_10357)
);

INVx2_ASAP7_75t_SL g10358 ( 
.A(n_9926),
.Y(n_10358)
);

INVx2_ASAP7_75t_L g10359 ( 
.A(n_10144),
.Y(n_10359)
);

NAND2x1p5_ASAP7_75t_L g10360 ( 
.A(n_10011),
.B(n_1140),
.Y(n_10360)
);

INVx1_ASAP7_75t_L g10361 ( 
.A(n_10059),
.Y(n_10361)
);

INVx2_ASAP7_75t_SL g10362 ( 
.A(n_10121),
.Y(n_10362)
);

INVx6_ASAP7_75t_L g10363 ( 
.A(n_9929),
.Y(n_10363)
);

OAI22xp5_ASAP7_75t_L g10364 ( 
.A1(n_10160),
.A2(n_1144),
.B1(n_1142),
.B2(n_1143),
.Y(n_10364)
);

AOI21x1_ASAP7_75t_L g10365 ( 
.A1(n_10032),
.A2(n_1142),
.B(n_1143),
.Y(n_10365)
);

INVx2_ASAP7_75t_SL g10366 ( 
.A(n_10121),
.Y(n_10366)
);

INVx1_ASAP7_75t_L g10367 ( 
.A(n_10064),
.Y(n_10367)
);

AND2x2_ASAP7_75t_L g10368 ( 
.A(n_10066),
.B(n_1144),
.Y(n_10368)
);

AND2x2_ASAP7_75t_L g10369 ( 
.A(n_10138),
.B(n_1145),
.Y(n_10369)
);

INVx1_ASAP7_75t_L g10370 ( 
.A(n_10099),
.Y(n_10370)
);

AND2x4_ASAP7_75t_L g10371 ( 
.A(n_10147),
.B(n_1145),
.Y(n_10371)
);

AOI22xp5_ASAP7_75t_L g10372 ( 
.A1(n_10040),
.A2(n_1148),
.B1(n_1146),
.B2(n_1147),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_10111),
.Y(n_10373)
);

BUFx2_ASAP7_75t_L g10374 ( 
.A(n_10171),
.Y(n_10374)
);

BUFx6f_ASAP7_75t_L g10375 ( 
.A(n_10024),
.Y(n_10375)
);

INVx2_ASAP7_75t_L g10376 ( 
.A(n_10174),
.Y(n_10376)
);

BUFx2_ASAP7_75t_L g10377 ( 
.A(n_9995),
.Y(n_10377)
);

INVx1_ASAP7_75t_L g10378 ( 
.A(n_10162),
.Y(n_10378)
);

AOI21x1_ASAP7_75t_L g10379 ( 
.A1(n_9913),
.A2(n_1147),
.B(n_1149),
.Y(n_10379)
);

INVx2_ASAP7_75t_L g10380 ( 
.A(n_10080),
.Y(n_10380)
);

INVx3_ASAP7_75t_L g10381 ( 
.A(n_9998),
.Y(n_10381)
);

INVx2_ASAP7_75t_L g10382 ( 
.A(n_10127),
.Y(n_10382)
);

AOI21x1_ASAP7_75t_L g10383 ( 
.A1(n_10158),
.A2(n_10016),
.B(n_9961),
.Y(n_10383)
);

INVx2_ASAP7_75t_L g10384 ( 
.A(n_10127),
.Y(n_10384)
);

OA21x2_ASAP7_75t_L g10385 ( 
.A1(n_9967),
.A2(n_1150),
.B(n_1151),
.Y(n_10385)
);

BUFx2_ASAP7_75t_L g10386 ( 
.A(n_10050),
.Y(n_10386)
);

INVx1_ASAP7_75t_L g10387 ( 
.A(n_10145),
.Y(n_10387)
);

INVx2_ASAP7_75t_L g10388 ( 
.A(n_10145),
.Y(n_10388)
);

INVxp67_ASAP7_75t_L g10389 ( 
.A(n_10045),
.Y(n_10389)
);

INVx2_ASAP7_75t_L g10390 ( 
.A(n_10003),
.Y(n_10390)
);

INVx2_ASAP7_75t_L g10391 ( 
.A(n_10003),
.Y(n_10391)
);

INVx1_ASAP7_75t_L g10392 ( 
.A(n_9931),
.Y(n_10392)
);

INVx1_ASAP7_75t_L g10393 ( 
.A(n_10007),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_10007),
.Y(n_10394)
);

INVx1_ASAP7_75t_L g10395 ( 
.A(n_10009),
.Y(n_10395)
);

INVx1_ASAP7_75t_L g10396 ( 
.A(n_10009),
.Y(n_10396)
);

INVx1_ASAP7_75t_L g10397 ( 
.A(n_10038),
.Y(n_10397)
);

INVx1_ASAP7_75t_L g10398 ( 
.A(n_10038),
.Y(n_10398)
);

INVx2_ASAP7_75t_L g10399 ( 
.A(n_10069),
.Y(n_10399)
);

INVx2_ASAP7_75t_L g10400 ( 
.A(n_10069),
.Y(n_10400)
);

INVx1_ASAP7_75t_L g10401 ( 
.A(n_10087),
.Y(n_10401)
);

AOI21x1_ASAP7_75t_L g10402 ( 
.A1(n_9937),
.A2(n_1150),
.B(n_1151),
.Y(n_10402)
);

INVx1_ASAP7_75t_L g10403 ( 
.A(n_10087),
.Y(n_10403)
);

INVx1_ASAP7_75t_L g10404 ( 
.A(n_10165),
.Y(n_10404)
);

BUFx4f_ASAP7_75t_SL g10405 ( 
.A(n_9886),
.Y(n_10405)
);

INVx1_ASAP7_75t_L g10406 ( 
.A(n_9974),
.Y(n_10406)
);

INVx2_ASAP7_75t_L g10407 ( 
.A(n_10132),
.Y(n_10407)
);

AOI22xp33_ASAP7_75t_SL g10408 ( 
.A1(n_9907),
.A2(n_1154),
.B1(n_1152),
.B2(n_1153),
.Y(n_10408)
);

OA21x2_ASAP7_75t_L g10409 ( 
.A1(n_10125),
.A2(n_1153),
.B(n_1155),
.Y(n_10409)
);

AOI22xp33_ASAP7_75t_SL g10410 ( 
.A1(n_10018),
.A2(n_1157),
.B1(n_1155),
.B2(n_1156),
.Y(n_10410)
);

BUFx2_ASAP7_75t_L g10411 ( 
.A(n_9973),
.Y(n_10411)
);

INVx2_ASAP7_75t_L g10412 ( 
.A(n_10132),
.Y(n_10412)
);

BUFx6f_ASAP7_75t_L g10413 ( 
.A(n_10098),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_9923),
.Y(n_10414)
);

INVx1_ASAP7_75t_L g10415 ( 
.A(n_9923),
.Y(n_10415)
);

INVx1_ASAP7_75t_L g10416 ( 
.A(n_9959),
.Y(n_10416)
);

INVx2_ASAP7_75t_L g10417 ( 
.A(n_9959),
.Y(n_10417)
);

NAND2xp5_ASAP7_75t_L g10418 ( 
.A(n_9969),
.B(n_1158),
.Y(n_10418)
);

INVx1_ASAP7_75t_L g10419 ( 
.A(n_10062),
.Y(n_10419)
);

INVx1_ASAP7_75t_L g10420 ( 
.A(n_10079),
.Y(n_10420)
);

INVx1_ASAP7_75t_L g10421 ( 
.A(n_9965),
.Y(n_10421)
);

HB1xp67_ASAP7_75t_L g10422 ( 
.A(n_9962),
.Y(n_10422)
);

INVx2_ASAP7_75t_L g10423 ( 
.A(n_10117),
.Y(n_10423)
);

INVx2_ASAP7_75t_L g10424 ( 
.A(n_10155),
.Y(n_10424)
);

BUFx12f_ASAP7_75t_L g10425 ( 
.A(n_10104),
.Y(n_10425)
);

INVx2_ASAP7_75t_L g10426 ( 
.A(n_10070),
.Y(n_10426)
);

INVx1_ASAP7_75t_L g10427 ( 
.A(n_9955),
.Y(n_10427)
);

INVx2_ASAP7_75t_L g10428 ( 
.A(n_10177),
.Y(n_10428)
);

BUFx8_ASAP7_75t_SL g10429 ( 
.A(n_10044),
.Y(n_10429)
);

INVx2_ASAP7_75t_L g10430 ( 
.A(n_10084),
.Y(n_10430)
);

HB1xp67_ASAP7_75t_L g10431 ( 
.A(n_9957),
.Y(n_10431)
);

INVx3_ASAP7_75t_L g10432 ( 
.A(n_10086),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_9922),
.Y(n_10433)
);

INVx1_ASAP7_75t_L g10434 ( 
.A(n_10129),
.Y(n_10434)
);

BUFx6f_ASAP7_75t_L g10435 ( 
.A(n_10122),
.Y(n_10435)
);

INVx1_ASAP7_75t_L g10436 ( 
.A(n_10118),
.Y(n_10436)
);

HB1xp67_ASAP7_75t_L g10437 ( 
.A(n_9981),
.Y(n_10437)
);

INVx6_ASAP7_75t_L g10438 ( 
.A(n_9976),
.Y(n_10438)
);

BUFx2_ASAP7_75t_L g10439 ( 
.A(n_10114),
.Y(n_10439)
);

INVx2_ASAP7_75t_L g10440 ( 
.A(n_10141),
.Y(n_10440)
);

HB1xp67_ASAP7_75t_L g10441 ( 
.A(n_10054),
.Y(n_10441)
);

INVx2_ASAP7_75t_L g10442 ( 
.A(n_10082),
.Y(n_10442)
);

INVx2_ASAP7_75t_L g10443 ( 
.A(n_9888),
.Y(n_10443)
);

AND2x2_ASAP7_75t_L g10444 ( 
.A(n_9960),
.B(n_1158),
.Y(n_10444)
);

BUFx4f_ASAP7_75t_SL g10445 ( 
.A(n_10106),
.Y(n_10445)
);

BUFx6f_ASAP7_75t_L g10446 ( 
.A(n_10151),
.Y(n_10446)
);

BUFx3_ASAP7_75t_L g10447 ( 
.A(n_10000),
.Y(n_10447)
);

OAI21x1_ASAP7_75t_L g10448 ( 
.A1(n_9947),
.A2(n_1159),
.B(n_1160),
.Y(n_10448)
);

BUFx3_ASAP7_75t_L g10449 ( 
.A(n_10140),
.Y(n_10449)
);

AOI22xp33_ASAP7_75t_L g10450 ( 
.A1(n_9881),
.A2(n_1164),
.B1(n_1161),
.B2(n_1163),
.Y(n_10450)
);

INVx3_ASAP7_75t_L g10451 ( 
.A(n_9945),
.Y(n_10451)
);

INVx2_ASAP7_75t_L g10452 ( 
.A(n_10102),
.Y(n_10452)
);

INVx2_ASAP7_75t_L g10453 ( 
.A(n_10172),
.Y(n_10453)
);

AOI22xp33_ASAP7_75t_L g10454 ( 
.A1(n_10019),
.A2(n_1165),
.B1(n_1163),
.B2(n_1164),
.Y(n_10454)
);

INVx2_ASAP7_75t_L g10455 ( 
.A(n_10078),
.Y(n_10455)
);

AND2x2_ASAP7_75t_L g10456 ( 
.A(n_9991),
.B(n_1165),
.Y(n_10456)
);

INVx1_ASAP7_75t_SL g10457 ( 
.A(n_9895),
.Y(n_10457)
);

INVx2_ASAP7_75t_SL g10458 ( 
.A(n_9918),
.Y(n_10458)
);

OR2x2_ASAP7_75t_L g10459 ( 
.A(n_9978),
.B(n_1166),
.Y(n_10459)
);

INVx1_ASAP7_75t_L g10460 ( 
.A(n_10097),
.Y(n_10460)
);

NAND2x1p5_ASAP7_75t_L g10461 ( 
.A(n_10028),
.B(n_1167),
.Y(n_10461)
);

AND2x4_ASAP7_75t_L g10462 ( 
.A(n_10123),
.B(n_1168),
.Y(n_10462)
);

INVx1_ASAP7_75t_L g10463 ( 
.A(n_10043),
.Y(n_10463)
);

INVx1_ASAP7_75t_L g10464 ( 
.A(n_10152),
.Y(n_10464)
);

OA21x2_ASAP7_75t_L g10465 ( 
.A1(n_9948),
.A2(n_1168),
.B(n_1169),
.Y(n_10465)
);

AND2x2_ASAP7_75t_L g10466 ( 
.A(n_9979),
.B(n_9928),
.Y(n_10466)
);

AOI22xp33_ASAP7_75t_L g10467 ( 
.A1(n_10134),
.A2(n_10181),
.B1(n_10119),
.B2(n_10092),
.Y(n_10467)
);

INVx2_ASAP7_75t_L g10468 ( 
.A(n_10112),
.Y(n_10468)
);

INVxp67_ASAP7_75t_SL g10469 ( 
.A(n_10176),
.Y(n_10469)
);

AOI22xp33_ASAP7_75t_SL g10470 ( 
.A1(n_10075),
.A2(n_1173),
.B1(n_1169),
.B2(n_1172),
.Y(n_10470)
);

INVx2_ASAP7_75t_L g10471 ( 
.A(n_9997),
.Y(n_10471)
);

CKINVDCx5p33_ASAP7_75t_R g10472 ( 
.A(n_10021),
.Y(n_10472)
);

BUFx3_ASAP7_75t_L g10473 ( 
.A(n_10169),
.Y(n_10473)
);

INVx3_ASAP7_75t_L g10474 ( 
.A(n_10124),
.Y(n_10474)
);

INVx3_ASAP7_75t_L g10475 ( 
.A(n_9925),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_10013),
.Y(n_10476)
);

INVx1_ASAP7_75t_L g10477 ( 
.A(n_10094),
.Y(n_10477)
);

INVx3_ASAP7_75t_L g10478 ( 
.A(n_10076),
.Y(n_10478)
);

INVx1_ASAP7_75t_L g10479 ( 
.A(n_10200),
.Y(n_10479)
);

INVx1_ASAP7_75t_L g10480 ( 
.A(n_10261),
.Y(n_10480)
);

INVx1_ASAP7_75t_L g10481 ( 
.A(n_10182),
.Y(n_10481)
);

INVx1_ASAP7_75t_L g10482 ( 
.A(n_10183),
.Y(n_10482)
);

OAI21x1_ASAP7_75t_L g10483 ( 
.A1(n_10198),
.A2(n_10116),
.B(n_10074),
.Y(n_10483)
);

AO21x1_ASAP7_75t_L g10484 ( 
.A1(n_10271),
.A2(n_10037),
.B(n_10149),
.Y(n_10484)
);

BUFx3_ASAP7_75t_L g10485 ( 
.A(n_10425),
.Y(n_10485)
);

OAI21x1_ASAP7_75t_L g10486 ( 
.A1(n_10192),
.A2(n_10091),
.B(n_10143),
.Y(n_10486)
);

INVx1_ASAP7_75t_L g10487 ( 
.A(n_10203),
.Y(n_10487)
);

INVx1_ASAP7_75t_L g10488 ( 
.A(n_10216),
.Y(n_10488)
);

INVx3_ASAP7_75t_L g10489 ( 
.A(n_10336),
.Y(n_10489)
);

INVx1_ASAP7_75t_L g10490 ( 
.A(n_10225),
.Y(n_10490)
);

AND2x4_ASAP7_75t_L g10491 ( 
.A(n_10377),
.B(n_10194),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_10226),
.Y(n_10492)
);

INVx2_ASAP7_75t_L g10493 ( 
.A(n_10228),
.Y(n_10493)
);

BUFx2_ASAP7_75t_L g10494 ( 
.A(n_10411),
.Y(n_10494)
);

INVx1_ASAP7_75t_L g10495 ( 
.A(n_10231),
.Y(n_10495)
);

BUFx6f_ASAP7_75t_L g10496 ( 
.A(n_10217),
.Y(n_10496)
);

NAND2xp5_ASAP7_75t_L g10497 ( 
.A(n_10243),
.B(n_10133),
.Y(n_10497)
);

OAI21xp5_ASAP7_75t_L g10498 ( 
.A1(n_10233),
.A2(n_10146),
.B(n_10027),
.Y(n_10498)
);

HB1xp67_ASAP7_75t_SL g10499 ( 
.A(n_10184),
.Y(n_10499)
);

INVx2_ASAP7_75t_L g10500 ( 
.A(n_10224),
.Y(n_10500)
);

AND2x2_ASAP7_75t_L g10501 ( 
.A(n_10234),
.B(n_10001),
.Y(n_10501)
);

HB1xp67_ASAP7_75t_L g10502 ( 
.A(n_10245),
.Y(n_10502)
);

INVx1_ASAP7_75t_L g10503 ( 
.A(n_10236),
.Y(n_10503)
);

INVx1_ASAP7_75t_L g10504 ( 
.A(n_10237),
.Y(n_10504)
);

INVx1_ASAP7_75t_L g10505 ( 
.A(n_10240),
.Y(n_10505)
);

OA21x2_ASAP7_75t_L g10506 ( 
.A1(n_10433),
.A2(n_10128),
.B(n_1173),
.Y(n_10506)
);

BUFx3_ASAP7_75t_L g10507 ( 
.A(n_10217),
.Y(n_10507)
);

INVx3_ASAP7_75t_L g10508 ( 
.A(n_10246),
.Y(n_10508)
);

OR2x2_ASAP7_75t_L g10509 ( 
.A(n_10275),
.B(n_1174),
.Y(n_10509)
);

INVx2_ASAP7_75t_L g10510 ( 
.A(n_10331),
.Y(n_10510)
);

OR2x6_ASAP7_75t_L g10511 ( 
.A(n_10212),
.B(n_10304),
.Y(n_10511)
);

INVx2_ASAP7_75t_L g10512 ( 
.A(n_10285),
.Y(n_10512)
);

BUFx2_ASAP7_75t_L g10513 ( 
.A(n_10268),
.Y(n_10513)
);

INVx1_ASAP7_75t_L g10514 ( 
.A(n_10247),
.Y(n_10514)
);

AND2x2_ASAP7_75t_L g10515 ( 
.A(n_10188),
.B(n_1174),
.Y(n_10515)
);

INVx1_ASAP7_75t_L g10516 ( 
.A(n_10250),
.Y(n_10516)
);

BUFx6f_ASAP7_75t_L g10517 ( 
.A(n_10304),
.Y(n_10517)
);

AOI21x1_ASAP7_75t_L g10518 ( 
.A1(n_10325),
.A2(n_1175),
.B(n_1176),
.Y(n_10518)
);

INVx1_ASAP7_75t_L g10519 ( 
.A(n_10252),
.Y(n_10519)
);

BUFx2_ASAP7_75t_L g10520 ( 
.A(n_10259),
.Y(n_10520)
);

OR2x2_ASAP7_75t_L g10521 ( 
.A(n_10199),
.B(n_1175),
.Y(n_10521)
);

OAI21xp5_ASAP7_75t_L g10522 ( 
.A1(n_10230),
.A2(n_1176),
.B(n_1178),
.Y(n_10522)
);

INVx1_ASAP7_75t_L g10523 ( 
.A(n_10253),
.Y(n_10523)
);

INVx2_ASAP7_75t_L g10524 ( 
.A(n_10407),
.Y(n_10524)
);

BUFx2_ASAP7_75t_L g10525 ( 
.A(n_10260),
.Y(n_10525)
);

HB1xp67_ASAP7_75t_L g10526 ( 
.A(n_10204),
.Y(n_10526)
);

AO31x2_ASAP7_75t_L g10527 ( 
.A1(n_10434),
.A2(n_1180),
.A3(n_1178),
.B(n_1179),
.Y(n_10527)
);

INVx2_ASAP7_75t_L g10528 ( 
.A(n_10412),
.Y(n_10528)
);

INVx1_ASAP7_75t_L g10529 ( 
.A(n_10185),
.Y(n_10529)
);

INVx1_ASAP7_75t_L g10530 ( 
.A(n_10273),
.Y(n_10530)
);

INVx1_ASAP7_75t_L g10531 ( 
.A(n_10277),
.Y(n_10531)
);

INVx2_ASAP7_75t_L g10532 ( 
.A(n_10326),
.Y(n_10532)
);

INVx2_ASAP7_75t_L g10533 ( 
.A(n_10328),
.Y(n_10533)
);

AND2x2_ASAP7_75t_L g10534 ( 
.A(n_10352),
.B(n_1180),
.Y(n_10534)
);

INVx2_ASAP7_75t_L g10535 ( 
.A(n_10238),
.Y(n_10535)
);

INVx2_ASAP7_75t_L g10536 ( 
.A(n_10359),
.Y(n_10536)
);

INVx2_ASAP7_75t_L g10537 ( 
.A(n_10335),
.Y(n_10537)
);

INVx2_ASAP7_75t_L g10538 ( 
.A(n_10264),
.Y(n_10538)
);

INVx1_ASAP7_75t_L g10539 ( 
.A(n_10282),
.Y(n_10539)
);

OAI21x1_ASAP7_75t_L g10540 ( 
.A1(n_10201),
.A2(n_1181),
.B(n_1182),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_10318),
.Y(n_10541)
);

INVx2_ASAP7_75t_L g10542 ( 
.A(n_10269),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_10297),
.Y(n_10543)
);

AND2x2_ASAP7_75t_L g10544 ( 
.A(n_10293),
.B(n_1181),
.Y(n_10544)
);

INVx1_ASAP7_75t_L g10545 ( 
.A(n_10298),
.Y(n_10545)
);

INVx1_ASAP7_75t_L g10546 ( 
.A(n_10299),
.Y(n_10546)
);

INVx2_ASAP7_75t_L g10547 ( 
.A(n_10279),
.Y(n_10547)
);

INVx2_ASAP7_75t_L g10548 ( 
.A(n_10254),
.Y(n_10548)
);

INVx1_ASAP7_75t_SL g10549 ( 
.A(n_10265),
.Y(n_10549)
);

INVx2_ASAP7_75t_L g10550 ( 
.A(n_10255),
.Y(n_10550)
);

NAND2xp5_ASAP7_75t_L g10551 ( 
.A(n_10251),
.B(n_10219),
.Y(n_10551)
);

INVx3_ASAP7_75t_L g10552 ( 
.A(n_10305),
.Y(n_10552)
);

INVx2_ASAP7_75t_L g10553 ( 
.A(n_10256),
.Y(n_10553)
);

AOI21xp33_ASAP7_75t_L g10554 ( 
.A1(n_10186),
.A2(n_1183),
.B(n_1184),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_10362),
.B(n_1183),
.Y(n_10555)
);

OR2x6_ASAP7_75t_L g10556 ( 
.A(n_10305),
.B(n_1184),
.Y(n_10556)
);

INVx2_ASAP7_75t_L g10557 ( 
.A(n_10262),
.Y(n_10557)
);

INVx2_ASAP7_75t_L g10558 ( 
.A(n_10189),
.Y(n_10558)
);

AND2x2_ASAP7_75t_L g10559 ( 
.A(n_10366),
.B(n_1185),
.Y(n_10559)
);

OAI21x1_ASAP7_75t_L g10560 ( 
.A1(n_10287),
.A2(n_1185),
.B(n_1186),
.Y(n_10560)
);

AND2x4_ASAP7_75t_L g10561 ( 
.A(n_10223),
.B(n_1186),
.Y(n_10561)
);

INVx1_ASAP7_75t_L g10562 ( 
.A(n_10218),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_10197),
.Y(n_10563)
);

INVx1_ASAP7_75t_L g10564 ( 
.A(n_10283),
.Y(n_10564)
);

AND2x4_ASAP7_75t_L g10565 ( 
.A(n_10257),
.B(n_10419),
.Y(n_10565)
);

AO21x1_ASAP7_75t_SL g10566 ( 
.A1(n_10427),
.A2(n_1187),
.B(n_1188),
.Y(n_10566)
);

HB1xp67_ASAP7_75t_L g10567 ( 
.A(n_10206),
.Y(n_10567)
);

BUFx3_ASAP7_75t_L g10568 ( 
.A(n_10429),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_10284),
.Y(n_10569)
);

INVx2_ASAP7_75t_L g10570 ( 
.A(n_10208),
.Y(n_10570)
);

INVx1_ASAP7_75t_L g10571 ( 
.A(n_10288),
.Y(n_10571)
);

BUFx3_ASAP7_75t_L g10572 ( 
.A(n_10375),
.Y(n_10572)
);

AO21x2_ASAP7_75t_L g10573 ( 
.A1(n_10422),
.A2(n_1187),
.B(n_1189),
.Y(n_10573)
);

INVx2_ASAP7_75t_L g10574 ( 
.A(n_10209),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_10267),
.Y(n_10575)
);

AND2x2_ASAP7_75t_L g10576 ( 
.A(n_10220),
.B(n_1189),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_10301),
.Y(n_10577)
);

INVx1_ASAP7_75t_L g10578 ( 
.A(n_10302),
.Y(n_10578)
);

INVx1_ASAP7_75t_L g10579 ( 
.A(n_10310),
.Y(n_10579)
);

INVx2_ASAP7_75t_L g10580 ( 
.A(n_10210),
.Y(n_10580)
);

OR2x2_ASAP7_75t_L g10581 ( 
.A(n_10290),
.B(n_1190),
.Y(n_10581)
);

BUFx2_ASAP7_75t_L g10582 ( 
.A(n_10374),
.Y(n_10582)
);

INVx1_ASAP7_75t_L g10583 ( 
.A(n_10190),
.Y(n_10583)
);

AND2x2_ASAP7_75t_L g10584 ( 
.A(n_10195),
.B(n_1190),
.Y(n_10584)
);

INVx2_ASAP7_75t_L g10585 ( 
.A(n_10211),
.Y(n_10585)
);

INVx3_ASAP7_75t_L g10586 ( 
.A(n_10375),
.Y(n_10586)
);

AND2x2_ASAP7_75t_L g10587 ( 
.A(n_10390),
.B(n_1191),
.Y(n_10587)
);

HB1xp67_ASAP7_75t_L g10588 ( 
.A(n_10187),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_10213),
.Y(n_10589)
);

OAI21x1_ASAP7_75t_L g10590 ( 
.A1(n_10248),
.A2(n_1191),
.B(n_1192),
.Y(n_10590)
);

INVx2_ASAP7_75t_L g10591 ( 
.A(n_10215),
.Y(n_10591)
);

INVx1_ASAP7_75t_L g10592 ( 
.A(n_10321),
.Y(n_10592)
);

INVx1_ASAP7_75t_L g10593 ( 
.A(n_10249),
.Y(n_10593)
);

INVxp67_ASAP7_75t_L g10594 ( 
.A(n_10409),
.Y(n_10594)
);

BUFx2_ASAP7_75t_L g10595 ( 
.A(n_10349),
.Y(n_10595)
);

HB1xp67_ASAP7_75t_L g10596 ( 
.A(n_10345),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_10289),
.Y(n_10597)
);

INVx2_ASAP7_75t_L g10598 ( 
.A(n_10229),
.Y(n_10598)
);

INVx1_ASAP7_75t_L g10599 ( 
.A(n_10291),
.Y(n_10599)
);

HB1xp67_ASAP7_75t_L g10600 ( 
.A(n_10196),
.Y(n_10600)
);

INVx4_ASAP7_75t_L g10601 ( 
.A(n_10413),
.Y(n_10601)
);

INVx1_ASAP7_75t_L g10602 ( 
.A(n_10295),
.Y(n_10602)
);

INVx2_ASAP7_75t_L g10603 ( 
.A(n_10239),
.Y(n_10603)
);

OAI21xp5_ASAP7_75t_L g10604 ( 
.A1(n_10232),
.A2(n_1192),
.B(n_1193),
.Y(n_10604)
);

INVx4_ASAP7_75t_L g10605 ( 
.A(n_10413),
.Y(n_10605)
);

CKINVDCx14_ASAP7_75t_R g10606 ( 
.A(n_10244),
.Y(n_10606)
);

HB1xp67_ASAP7_75t_L g10607 ( 
.A(n_10350),
.Y(n_10607)
);

INVx2_ASAP7_75t_SL g10608 ( 
.A(n_10222),
.Y(n_10608)
);

AND2x2_ASAP7_75t_L g10609 ( 
.A(n_10391),
.B(n_1194),
.Y(n_10609)
);

INVx2_ASAP7_75t_L g10610 ( 
.A(n_10241),
.Y(n_10610)
);

INVx1_ASAP7_75t_L g10611 ( 
.A(n_10306),
.Y(n_10611)
);

OR2x2_ASAP7_75t_L g10612 ( 
.A(n_10351),
.B(n_10340),
.Y(n_10612)
);

AO21x2_ASAP7_75t_L g10613 ( 
.A1(n_10378),
.A2(n_10420),
.B(n_10383),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_10309),
.Y(n_10614)
);

INVx1_ASAP7_75t_L g10615 ( 
.A(n_10320),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_10227),
.Y(n_10616)
);

INVx1_ASAP7_75t_L g10617 ( 
.A(n_10333),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_10281),
.Y(n_10618)
);

AND2x2_ASAP7_75t_L g10619 ( 
.A(n_10399),
.B(n_1194),
.Y(n_10619)
);

AOI21x1_ASAP7_75t_L g10620 ( 
.A1(n_10439),
.A2(n_1195),
.B(n_1196),
.Y(n_10620)
);

INVx2_ASAP7_75t_L g10621 ( 
.A(n_10339),
.Y(n_10621)
);

HB1xp67_ASAP7_75t_L g10622 ( 
.A(n_10332),
.Y(n_10622)
);

BUFx2_ASAP7_75t_L g10623 ( 
.A(n_10311),
.Y(n_10623)
);

OR2x2_ASAP7_75t_L g10624 ( 
.A(n_10312),
.B(n_1195),
.Y(n_10624)
);

INVx1_ASAP7_75t_L g10625 ( 
.A(n_10334),
.Y(n_10625)
);

INVx1_ASAP7_75t_L g10626 ( 
.A(n_10356),
.Y(n_10626)
);

INVxp67_ASAP7_75t_SL g10627 ( 
.A(n_10389),
.Y(n_10627)
);

NOR2xp33_ASAP7_75t_L g10628 ( 
.A(n_10292),
.B(n_1197),
.Y(n_10628)
);

INVx1_ASAP7_75t_L g10629 ( 
.A(n_10207),
.Y(n_10629)
);

INVx2_ASAP7_75t_L g10630 ( 
.A(n_10400),
.Y(n_10630)
);

INVx1_ASAP7_75t_L g10631 ( 
.A(n_10221),
.Y(n_10631)
);

HB1xp67_ASAP7_75t_L g10632 ( 
.A(n_10276),
.Y(n_10632)
);

BUFx6f_ASAP7_75t_L g10633 ( 
.A(n_10193),
.Y(n_10633)
);

INVx1_ASAP7_75t_L g10634 ( 
.A(n_10263),
.Y(n_10634)
);

INVx1_ASAP7_75t_L g10635 ( 
.A(n_10464),
.Y(n_10635)
);

INVx1_ASAP7_75t_L g10636 ( 
.A(n_10300),
.Y(n_10636)
);

AO21x2_ASAP7_75t_L g10637 ( 
.A1(n_10402),
.A2(n_1197),
.B(n_1198),
.Y(n_10637)
);

OAI21x1_ASAP7_75t_L g10638 ( 
.A1(n_10344),
.A2(n_1199),
.B(n_1200),
.Y(n_10638)
);

BUFx2_ASAP7_75t_L g10639 ( 
.A(n_10314),
.Y(n_10639)
);

OAI21xp5_ASAP7_75t_L g10640 ( 
.A1(n_10274),
.A2(n_1200),
.B(n_1201),
.Y(n_10640)
);

INVx3_ASAP7_75t_L g10641 ( 
.A(n_10242),
.Y(n_10641)
);

AO21x2_ASAP7_75t_L g10642 ( 
.A1(n_10404),
.A2(n_1202),
.B(n_1203),
.Y(n_10642)
);

BUFx3_ASAP7_75t_L g10643 ( 
.A(n_10266),
.Y(n_10643)
);

AND2x2_ASAP7_75t_L g10644 ( 
.A(n_10191),
.B(n_10406),
.Y(n_10644)
);

INVx1_ASAP7_75t_L g10645 ( 
.A(n_10463),
.Y(n_10645)
);

INVx2_ASAP7_75t_L g10646 ( 
.A(n_10443),
.Y(n_10646)
);

INVx1_ASAP7_75t_L g10647 ( 
.A(n_10286),
.Y(n_10647)
);

AND2x2_ASAP7_75t_L g10648 ( 
.A(n_10393),
.B(n_1202),
.Y(n_10648)
);

OAI21x1_ASAP7_75t_L g10649 ( 
.A1(n_10341),
.A2(n_1203),
.B(n_1204),
.Y(n_10649)
);

INVx1_ASAP7_75t_L g10650 ( 
.A(n_10353),
.Y(n_10650)
);

INVx2_ASAP7_75t_L g10651 ( 
.A(n_10348),
.Y(n_10651)
);

AND3x2_ASAP7_75t_L g10652 ( 
.A(n_10431),
.B(n_10441),
.C(n_10437),
.Y(n_10652)
);

HB1xp67_ASAP7_75t_L g10653 ( 
.A(n_10258),
.Y(n_10653)
);

INVx1_ASAP7_75t_L g10654 ( 
.A(n_10361),
.Y(n_10654)
);

NAND2xp5_ASAP7_75t_L g10655 ( 
.A(n_10466),
.B(n_1204),
.Y(n_10655)
);

INVx3_ASAP7_75t_L g10656 ( 
.A(n_10363),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_10367),
.Y(n_10657)
);

NAND2xp5_ASAP7_75t_L g10658 ( 
.A(n_10458),
.B(n_1205),
.Y(n_10658)
);

HB1xp67_ASAP7_75t_SL g10659 ( 
.A(n_10473),
.Y(n_10659)
);

INVx1_ASAP7_75t_L g10660 ( 
.A(n_10460),
.Y(n_10660)
);

AND2x2_ASAP7_75t_L g10661 ( 
.A(n_10394),
.B(n_10395),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_10330),
.Y(n_10662)
);

INVx4_ASAP7_75t_L g10663 ( 
.A(n_10435),
.Y(n_10663)
);

OA21x2_ASAP7_75t_L g10664 ( 
.A1(n_10457),
.A2(n_1206),
.B(n_1207),
.Y(n_10664)
);

INVx2_ASAP7_75t_L g10665 ( 
.A(n_10396),
.Y(n_10665)
);

INVx2_ASAP7_75t_L g10666 ( 
.A(n_10397),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_10398),
.Y(n_10667)
);

HB1xp67_ASAP7_75t_L g10668 ( 
.A(n_10278),
.Y(n_10668)
);

INVx1_ASAP7_75t_L g10669 ( 
.A(n_10401),
.Y(n_10669)
);

INVx1_ASAP7_75t_L g10670 ( 
.A(n_10403),
.Y(n_10670)
);

INVx1_ASAP7_75t_L g10671 ( 
.A(n_10414),
.Y(n_10671)
);

BUFx6f_ASAP7_75t_L g10672 ( 
.A(n_10435),
.Y(n_10672)
);

INVx5_ASAP7_75t_L g10673 ( 
.A(n_10322),
.Y(n_10673)
);

INVx1_ASAP7_75t_L g10674 ( 
.A(n_10415),
.Y(n_10674)
);

INVx1_ASAP7_75t_L g10675 ( 
.A(n_10416),
.Y(n_10675)
);

INVx1_ASAP7_75t_L g10676 ( 
.A(n_10392),
.Y(n_10676)
);

INVx1_ASAP7_75t_L g10677 ( 
.A(n_10421),
.Y(n_10677)
);

INVxp67_ASAP7_75t_L g10678 ( 
.A(n_10446),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_10455),
.Y(n_10679)
);

INVx1_ASAP7_75t_L g10680 ( 
.A(n_10417),
.Y(n_10680)
);

OAI21x1_ASAP7_75t_L g10681 ( 
.A1(n_10376),
.A2(n_1206),
.B(n_1207),
.Y(n_10681)
);

OA21x2_ASAP7_75t_L g10682 ( 
.A1(n_10205),
.A2(n_1208),
.B(n_1209),
.Y(n_10682)
);

AO31x2_ASAP7_75t_L g10683 ( 
.A1(n_10342),
.A2(n_1212),
.A3(n_1209),
.B(n_1210),
.Y(n_10683)
);

INVx4_ASAP7_75t_L g10684 ( 
.A(n_10357),
.Y(n_10684)
);

AND2x2_ASAP7_75t_L g10685 ( 
.A(n_10235),
.B(n_1210),
.Y(n_10685)
);

AO21x1_ASAP7_75t_L g10686 ( 
.A1(n_10294),
.A2(n_1212),
.B(n_1213),
.Y(n_10686)
);

OAI21x1_ASAP7_75t_L g10687 ( 
.A1(n_10370),
.A2(n_1213),
.B(n_1215),
.Y(n_10687)
);

AND2x2_ASAP7_75t_L g10688 ( 
.A(n_10316),
.B(n_1215),
.Y(n_10688)
);

NOR2x1_ASAP7_75t_L g10689 ( 
.A(n_10451),
.B(n_1216),
.Y(n_10689)
);

NAND2xp5_ASAP7_75t_L g10690 ( 
.A(n_10453),
.B(n_1216),
.Y(n_10690)
);

NOR2x1_ASAP7_75t_SL g10691 ( 
.A(n_10202),
.B(n_1217),
.Y(n_10691)
);

INVx1_ASAP7_75t_L g10692 ( 
.A(n_10347),
.Y(n_10692)
);

BUFx2_ASAP7_75t_L g10693 ( 
.A(n_10440),
.Y(n_10693)
);

NAND2xp5_ASAP7_75t_L g10694 ( 
.A(n_10452),
.B(n_1217),
.Y(n_10694)
);

AND2x4_ASAP7_75t_L g10695 ( 
.A(n_10343),
.B(n_1218),
.Y(n_10695)
);

INVx1_ASAP7_75t_L g10696 ( 
.A(n_10280),
.Y(n_10696)
);

AND2x2_ASAP7_75t_L g10697 ( 
.A(n_10317),
.B(n_10382),
.Y(n_10697)
);

OAI21xp5_ASAP7_75t_L g10698 ( 
.A1(n_10469),
.A2(n_1219),
.B(n_1221),
.Y(n_10698)
);

BUFx2_ASAP7_75t_L g10699 ( 
.A(n_10307),
.Y(n_10699)
);

INVx1_ASAP7_75t_L g10700 ( 
.A(n_10387),
.Y(n_10700)
);

BUFx2_ASAP7_75t_L g10701 ( 
.A(n_10308),
.Y(n_10701)
);

INVxp67_ASAP7_75t_L g10702 ( 
.A(n_10446),
.Y(n_10702)
);

AND2x2_ASAP7_75t_L g10703 ( 
.A(n_10384),
.B(n_1219),
.Y(n_10703)
);

AO21x1_ASAP7_75t_SL g10704 ( 
.A1(n_10296),
.A2(n_1222),
.B(n_1223),
.Y(n_10704)
);

OA21x2_ASAP7_75t_L g10705 ( 
.A1(n_10388),
.A2(n_1223),
.B(n_1224),
.Y(n_10705)
);

BUFx3_ASAP7_75t_R g10706 ( 
.A(n_10386),
.Y(n_10706)
);

AND2x2_ASAP7_75t_L g10707 ( 
.A(n_10327),
.B(n_1225),
.Y(n_10707)
);

INVx1_ASAP7_75t_L g10708 ( 
.A(n_10373),
.Y(n_10708)
);

INVx1_ASAP7_75t_L g10709 ( 
.A(n_10365),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_10380),
.Y(n_10710)
);

INVx1_ASAP7_75t_L g10711 ( 
.A(n_10436),
.Y(n_10711)
);

INVx2_ASAP7_75t_L g10712 ( 
.A(n_10354),
.Y(n_10712)
);

INVx2_ASAP7_75t_L g10713 ( 
.A(n_10358),
.Y(n_10713)
);

NAND2xp5_ASAP7_75t_L g10714 ( 
.A(n_10475),
.B(n_1225),
.Y(n_10714)
);

INVx1_ASAP7_75t_L g10715 ( 
.A(n_10368),
.Y(n_10715)
);

INVx2_ASAP7_75t_L g10716 ( 
.A(n_10315),
.Y(n_10716)
);

INVx2_ASAP7_75t_L g10717 ( 
.A(n_10428),
.Y(n_10717)
);

HB1xp67_ASAP7_75t_L g10718 ( 
.A(n_10379),
.Y(n_10718)
);

BUFx3_ASAP7_75t_L g10719 ( 
.A(n_10426),
.Y(n_10719)
);

INVx1_ASAP7_75t_L g10720 ( 
.A(n_10471),
.Y(n_10720)
);

INVx1_ASAP7_75t_L g10721 ( 
.A(n_10468),
.Y(n_10721)
);

BUFx6f_ASAP7_75t_L g10722 ( 
.A(n_10323),
.Y(n_10722)
);

INVx1_ASAP7_75t_L g10723 ( 
.A(n_10319),
.Y(n_10723)
);

OR2x2_ASAP7_75t_L g10724 ( 
.A(n_10477),
.B(n_1226),
.Y(n_10724)
);

OR2x2_ASAP7_75t_L g10725 ( 
.A(n_10476),
.B(n_1227),
.Y(n_10725)
);

INVx3_ASAP7_75t_L g10726 ( 
.A(n_10381),
.Y(n_10726)
);

INVx1_ASAP7_75t_L g10727 ( 
.A(n_10385),
.Y(n_10727)
);

INVx1_ASAP7_75t_L g10728 ( 
.A(n_10346),
.Y(n_10728)
);

HB1xp67_ASAP7_75t_L g10729 ( 
.A(n_10465),
.Y(n_10729)
);

AND2x4_ASAP7_75t_L g10730 ( 
.A(n_10442),
.B(n_1227),
.Y(n_10730)
);

INVx2_ASAP7_75t_SL g10731 ( 
.A(n_10214),
.Y(n_10731)
);

BUFx2_ASAP7_75t_L g10732 ( 
.A(n_10445),
.Y(n_10732)
);

AO21x2_ASAP7_75t_L g10733 ( 
.A1(n_10418),
.A2(n_1228),
.B(n_1229),
.Y(n_10733)
);

AO21x2_ASAP7_75t_L g10734 ( 
.A1(n_10369),
.A2(n_1229),
.B(n_1230),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_10459),
.Y(n_10735)
);

AOI21x1_ASAP7_75t_L g10736 ( 
.A1(n_10423),
.A2(n_1231),
.B(n_1232),
.Y(n_10736)
);

AND2x2_ASAP7_75t_L g10737 ( 
.A(n_10329),
.B(n_1231),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_10449),
.Y(n_10738)
);

INVx2_ASAP7_75t_L g10739 ( 
.A(n_10371),
.Y(n_10739)
);

AND2x4_ASAP7_75t_L g10740 ( 
.A(n_10430),
.B(n_1232),
.Y(n_10740)
);

INVx2_ASAP7_75t_L g10741 ( 
.A(n_10447),
.Y(n_10741)
);

NAND2xp5_ASAP7_75t_L g10742 ( 
.A(n_10478),
.B(n_1233),
.Y(n_10742)
);

INVx2_ASAP7_75t_L g10743 ( 
.A(n_10432),
.Y(n_10743)
);

INVx2_ASAP7_75t_L g10744 ( 
.A(n_10438),
.Y(n_10744)
);

AO21x2_ASAP7_75t_L g10745 ( 
.A1(n_10355),
.A2(n_10456),
.B(n_10424),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_10448),
.Y(n_10746)
);

INVx1_ASAP7_75t_L g10747 ( 
.A(n_10444),
.Y(n_10747)
);

INVx3_ASAP7_75t_L g10748 ( 
.A(n_10405),
.Y(n_10748)
);

AND2x2_ASAP7_75t_L g10749 ( 
.A(n_10270),
.B(n_10313),
.Y(n_10749)
);

INVx1_ASAP7_75t_L g10750 ( 
.A(n_10474),
.Y(n_10750)
);

OAI21x1_ASAP7_75t_L g10751 ( 
.A1(n_10360),
.A2(n_1233),
.B(n_1235),
.Y(n_10751)
);

HB1xp67_ASAP7_75t_L g10752 ( 
.A(n_10462),
.Y(n_10752)
);

INVx1_ASAP7_75t_L g10753 ( 
.A(n_10303),
.Y(n_10753)
);

AND2x2_ASAP7_75t_L g10754 ( 
.A(n_10324),
.B(n_1235),
.Y(n_10754)
);

AND2x2_ASAP7_75t_L g10755 ( 
.A(n_10337),
.B(n_1237),
.Y(n_10755)
);

BUFx2_ASAP7_75t_L g10756 ( 
.A(n_10472),
.Y(n_10756)
);

AO31x2_ASAP7_75t_L g10757 ( 
.A1(n_10364),
.A2(n_1240),
.A3(n_1237),
.B(n_1238),
.Y(n_10757)
);

BUFx3_ASAP7_75t_L g10758 ( 
.A(n_10461),
.Y(n_10758)
);

OAI21x1_ASAP7_75t_L g10759 ( 
.A1(n_10272),
.A2(n_1241),
.B(n_1242),
.Y(n_10759)
);

INVx2_ASAP7_75t_L g10760 ( 
.A(n_10372),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_10338),
.Y(n_10761)
);

AND2x2_ASAP7_75t_L g10762 ( 
.A(n_10408),
.B(n_1241),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_10410),
.Y(n_10763)
);

BUFx2_ASAP7_75t_L g10764 ( 
.A(n_10450),
.Y(n_10764)
);

INVx1_ASAP7_75t_L g10765 ( 
.A(n_10467),
.Y(n_10765)
);

AND2x4_ASAP7_75t_L g10766 ( 
.A(n_10454),
.B(n_1243),
.Y(n_10766)
);

INVx1_ASAP7_75t_L g10767 ( 
.A(n_10470),
.Y(n_10767)
);

AND2x2_ASAP7_75t_L g10768 ( 
.A(n_10377),
.B(n_1243),
.Y(n_10768)
);

INVx1_ASAP7_75t_L g10769 ( 
.A(n_10200),
.Y(n_10769)
);

INVx2_ASAP7_75t_L g10770 ( 
.A(n_10377),
.Y(n_10770)
);

INVx1_ASAP7_75t_L g10771 ( 
.A(n_10200),
.Y(n_10771)
);

BUFx3_ASAP7_75t_L g10772 ( 
.A(n_10425),
.Y(n_10772)
);

OA21x2_ASAP7_75t_L g10773 ( 
.A1(n_10271),
.A2(n_1244),
.B(n_1245),
.Y(n_10773)
);

AND2x2_ASAP7_75t_L g10774 ( 
.A(n_10377),
.B(n_1244),
.Y(n_10774)
);

AND2x2_ASAP7_75t_L g10775 ( 
.A(n_10377),
.B(n_1245),
.Y(n_10775)
);

BUFx12f_ASAP7_75t_L g10776 ( 
.A(n_10244),
.Y(n_10776)
);

INVx1_ASAP7_75t_L g10777 ( 
.A(n_10200),
.Y(n_10777)
);

HB1xp67_ASAP7_75t_L g10778 ( 
.A(n_10245),
.Y(n_10778)
);

INVx3_ASAP7_75t_L g10779 ( 
.A(n_10336),
.Y(n_10779)
);

INVx1_ASAP7_75t_L g10780 ( 
.A(n_10200),
.Y(n_10780)
);

INVx2_ASAP7_75t_L g10781 ( 
.A(n_10377),
.Y(n_10781)
);

BUFx3_ASAP7_75t_L g10782 ( 
.A(n_10425),
.Y(n_10782)
);

INVx3_ASAP7_75t_L g10783 ( 
.A(n_10336),
.Y(n_10783)
);

OR2x2_ASAP7_75t_L g10784 ( 
.A(n_10275),
.B(n_1246),
.Y(n_10784)
);

HB1xp67_ASAP7_75t_L g10785 ( 
.A(n_10245),
.Y(n_10785)
);

AND2x2_ASAP7_75t_L g10786 ( 
.A(n_10377),
.B(n_1247),
.Y(n_10786)
);

AND2x2_ASAP7_75t_L g10787 ( 
.A(n_10377),
.B(n_1247),
.Y(n_10787)
);

INVx2_ASAP7_75t_L g10788 ( 
.A(n_10377),
.Y(n_10788)
);

INVx1_ASAP7_75t_L g10789 ( 
.A(n_10200),
.Y(n_10789)
);

BUFx12f_ASAP7_75t_L g10790 ( 
.A(n_10244),
.Y(n_10790)
);

INVx3_ASAP7_75t_L g10791 ( 
.A(n_10336),
.Y(n_10791)
);

INVx1_ASAP7_75t_L g10792 ( 
.A(n_10200),
.Y(n_10792)
);

OAI222xp33_ASAP7_75t_L g10793 ( 
.A1(n_10325),
.A2(n_1250),
.B1(n_1253),
.B2(n_1248),
.C1(n_1249),
.C2(n_1251),
.Y(n_10793)
);

INVx2_ASAP7_75t_L g10794 ( 
.A(n_10377),
.Y(n_10794)
);

AND2x2_ASAP7_75t_L g10795 ( 
.A(n_10377),
.B(n_1248),
.Y(n_10795)
);

NOR2xp33_ASAP7_75t_L g10796 ( 
.A(n_10606),
.B(n_1250),
.Y(n_10796)
);

INVx1_ASAP7_75t_L g10797 ( 
.A(n_10607),
.Y(n_10797)
);

A2O1A1Ixp33_ASAP7_75t_L g10798 ( 
.A1(n_10604),
.A2(n_1254),
.B(n_1251),
.C(n_1253),
.Y(n_10798)
);

AND2x2_ASAP7_75t_L g10799 ( 
.A(n_10582),
.B(n_1255),
.Y(n_10799)
);

INVx1_ASAP7_75t_L g10800 ( 
.A(n_10596),
.Y(n_10800)
);

OR2x2_ASAP7_75t_L g10801 ( 
.A(n_10595),
.B(n_1255),
.Y(n_10801)
);

AND2x2_ASAP7_75t_L g10802 ( 
.A(n_10494),
.B(n_1257),
.Y(n_10802)
);

INVx1_ASAP7_75t_L g10803 ( 
.A(n_10479),
.Y(n_10803)
);

NOR2xp33_ASAP7_75t_L g10804 ( 
.A(n_10499),
.B(n_1257),
.Y(n_10804)
);

OAI22xp5_ASAP7_75t_L g10805 ( 
.A1(n_10659),
.A2(n_1260),
.B1(n_1258),
.B2(n_1259),
.Y(n_10805)
);

INVx1_ASAP7_75t_L g10806 ( 
.A(n_10480),
.Y(n_10806)
);

INVx2_ASAP7_75t_L g10807 ( 
.A(n_10693),
.Y(n_10807)
);

BUFx3_ASAP7_75t_L g10808 ( 
.A(n_10776),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_10481),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_10482),
.Y(n_10810)
);

INVxp67_ASAP7_75t_L g10811 ( 
.A(n_10566),
.Y(n_10811)
);

AND2x4_ASAP7_75t_L g10812 ( 
.A(n_10491),
.B(n_1258),
.Y(n_10812)
);

AND2x4_ASAP7_75t_L g10813 ( 
.A(n_10508),
.B(n_1259),
.Y(n_10813)
);

AOI221xp5_ASAP7_75t_L g10814 ( 
.A1(n_10522),
.A2(n_1262),
.B1(n_1260),
.B2(n_1261),
.C(n_1263),
.Y(n_10814)
);

AOI21xp5_ASAP7_75t_L g10815 ( 
.A1(n_10484),
.A2(n_1261),
.B(n_1262),
.Y(n_10815)
);

INVx3_ASAP7_75t_L g10816 ( 
.A(n_10790),
.Y(n_10816)
);

AND2x4_ASAP7_75t_L g10817 ( 
.A(n_10513),
.B(n_1263),
.Y(n_10817)
);

AOI221xp5_ASAP7_75t_L g10818 ( 
.A1(n_10653),
.A2(n_1267),
.B1(n_1264),
.B2(n_1265),
.C(n_1268),
.Y(n_10818)
);

O2A1O1Ixp33_ASAP7_75t_L g10819 ( 
.A1(n_10594),
.A2(n_1268),
.B(n_1264),
.C(n_1267),
.Y(n_10819)
);

NAND2xp33_ASAP7_75t_R g10820 ( 
.A(n_10652),
.B(n_10773),
.Y(n_10820)
);

OAI21xp5_ASAP7_75t_L g10821 ( 
.A1(n_10640),
.A2(n_1269),
.B(n_1271),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_10487),
.Y(n_10822)
);

AOI21xp5_ASAP7_75t_L g10823 ( 
.A1(n_10497),
.A2(n_1269),
.B(n_1271),
.Y(n_10823)
);

OAI21xp5_ASAP7_75t_L g10824 ( 
.A1(n_10622),
.A2(n_1272),
.B(n_1273),
.Y(n_10824)
);

AND2x2_ASAP7_75t_L g10825 ( 
.A(n_10623),
.B(n_1272),
.Y(n_10825)
);

AOI22xp5_ASAP7_75t_L g10826 ( 
.A1(n_10686),
.A2(n_1275),
.B1(n_1273),
.B2(n_1274),
.Y(n_10826)
);

O2A1O1Ixp33_ASAP7_75t_L g10827 ( 
.A1(n_10729),
.A2(n_10793),
.B(n_10632),
.C(n_10718),
.Y(n_10827)
);

BUFx6f_ASAP7_75t_L g10828 ( 
.A(n_10496),
.Y(n_10828)
);

NAND2xp5_ASAP7_75t_L g10829 ( 
.A(n_10727),
.B(n_1276),
.Y(n_10829)
);

AND2x4_ASAP7_75t_L g10830 ( 
.A(n_10489),
.B(n_1276),
.Y(n_10830)
);

AND2x2_ASAP7_75t_L g10831 ( 
.A(n_10520),
.B(n_1277),
.Y(n_10831)
);

NAND2xp5_ASAP7_75t_L g10832 ( 
.A(n_10745),
.B(n_1277),
.Y(n_10832)
);

INVx2_ASAP7_75t_L g10833 ( 
.A(n_10719),
.Y(n_10833)
);

NOR2xp33_ASAP7_75t_L g10834 ( 
.A(n_10601),
.B(n_1278),
.Y(n_10834)
);

AO32x2_ASAP7_75t_L g10835 ( 
.A1(n_10706),
.A2(n_1281),
.A3(n_1279),
.B1(n_1280),
.B2(n_1282),
.Y(n_10835)
);

AND2x2_ASAP7_75t_L g10836 ( 
.A(n_10525),
.B(n_1279),
.Y(n_10836)
);

CKINVDCx5p33_ASAP7_75t_R g10837 ( 
.A(n_10568),
.Y(n_10837)
);

AO32x2_ASAP7_75t_L g10838 ( 
.A1(n_10731),
.A2(n_1282),
.A3(n_1280),
.B1(n_1281),
.B2(n_1283),
.Y(n_10838)
);

INVx2_ASAP7_75t_L g10839 ( 
.A(n_10639),
.Y(n_10839)
);

BUFx3_ASAP7_75t_L g10840 ( 
.A(n_10485),
.Y(n_10840)
);

INVx3_ASAP7_75t_L g10841 ( 
.A(n_10605),
.Y(n_10841)
);

OAI22xp5_ASAP7_75t_L g10842 ( 
.A1(n_10761),
.A2(n_1285),
.B1(n_1283),
.B2(n_1284),
.Y(n_10842)
);

INVx2_ASAP7_75t_SL g10843 ( 
.A(n_10496),
.Y(n_10843)
);

AND2x2_ASAP7_75t_L g10844 ( 
.A(n_10779),
.B(n_1285),
.Y(n_10844)
);

INVx2_ASAP7_75t_L g10845 ( 
.A(n_10783),
.Y(n_10845)
);

OA21x2_ASAP7_75t_L g10846 ( 
.A1(n_10551),
.A2(n_1286),
.B(n_1287),
.Y(n_10846)
);

NOR2xp33_ASAP7_75t_SL g10847 ( 
.A(n_10549),
.B(n_1287),
.Y(n_10847)
);

AND2x2_ASAP7_75t_L g10848 ( 
.A(n_10791),
.B(n_1289),
.Y(n_10848)
);

AO32x2_ASAP7_75t_L g10849 ( 
.A1(n_10663),
.A2(n_1291),
.A3(n_1289),
.B1(n_1290),
.B2(n_1292),
.Y(n_10849)
);

NOR2x1_ASAP7_75t_SL g10850 ( 
.A(n_10613),
.B(n_1290),
.Y(n_10850)
);

AND2x2_ASAP7_75t_L g10851 ( 
.A(n_10699),
.B(n_10701),
.Y(n_10851)
);

O2A1O1Ixp33_ASAP7_75t_L g10852 ( 
.A1(n_10554),
.A2(n_1295),
.B(n_1293),
.C(n_1294),
.Y(n_10852)
);

AND2x4_ASAP7_75t_L g10853 ( 
.A(n_10726),
.B(n_1293),
.Y(n_10853)
);

A2O1A1Ixp33_ASAP7_75t_L g10854 ( 
.A1(n_10689),
.A2(n_1298),
.B(n_1294),
.C(n_1296),
.Y(n_10854)
);

OAI22xp5_ASAP7_75t_L g10855 ( 
.A1(n_10627),
.A2(n_1299),
.B1(n_1296),
.B2(n_1298),
.Y(n_10855)
);

AND2x2_ASAP7_75t_L g10856 ( 
.A(n_10770),
.B(n_10781),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_10488),
.Y(n_10857)
);

AND2x2_ASAP7_75t_L g10858 ( 
.A(n_10788),
.B(n_1300),
.Y(n_10858)
);

NAND2xp5_ASAP7_75t_L g10859 ( 
.A(n_10738),
.B(n_10741),
.Y(n_10859)
);

A2O1A1Ixp33_ASAP7_75t_L g10860 ( 
.A1(n_10486),
.A2(n_1303),
.B(n_1301),
.C(n_1302),
.Y(n_10860)
);

INVxp67_ASAP7_75t_L g10861 ( 
.A(n_10756),
.Y(n_10861)
);

NAND2xp5_ASAP7_75t_L g10862 ( 
.A(n_10683),
.B(n_1301),
.Y(n_10862)
);

INVx2_ASAP7_75t_L g10863 ( 
.A(n_10565),
.Y(n_10863)
);

AND2x2_ASAP7_75t_L g10864 ( 
.A(n_10794),
.B(n_1302),
.Y(n_10864)
);

AND2x2_ASAP7_75t_L g10865 ( 
.A(n_10644),
.B(n_1303),
.Y(n_10865)
);

CKINVDCx20_ASAP7_75t_R g10866 ( 
.A(n_10772),
.Y(n_10866)
);

OAI21xp5_ASAP7_75t_L g10867 ( 
.A1(n_10518),
.A2(n_1304),
.B(n_1305),
.Y(n_10867)
);

O2A1O1Ixp33_ASAP7_75t_SL g10868 ( 
.A1(n_10763),
.A2(n_1307),
.B(n_1305),
.C(n_1306),
.Y(n_10868)
);

AOI21xp5_ASAP7_75t_L g10869 ( 
.A1(n_10691),
.A2(n_1306),
.B(n_1308),
.Y(n_10869)
);

BUFx6f_ASAP7_75t_L g10870 ( 
.A(n_10517),
.Y(n_10870)
);

INVx2_ASAP7_75t_L g10871 ( 
.A(n_10511),
.Y(n_10871)
);

AND2x2_ASAP7_75t_L g10872 ( 
.A(n_10493),
.B(n_1309),
.Y(n_10872)
);

OR2x2_ASAP7_75t_L g10873 ( 
.A(n_10612),
.B(n_1309),
.Y(n_10873)
);

INVxp67_ASAP7_75t_L g10874 ( 
.A(n_10682),
.Y(n_10874)
);

NAND2xp5_ASAP7_75t_L g10875 ( 
.A(n_10683),
.B(n_1310),
.Y(n_10875)
);

AOI22xp5_ASAP7_75t_L g10876 ( 
.A1(n_10678),
.A2(n_1313),
.B1(n_1310),
.B2(n_1312),
.Y(n_10876)
);

O2A1O1Ixp33_ASAP7_75t_L g10877 ( 
.A1(n_10702),
.A2(n_1314),
.B(n_1312),
.C(n_1313),
.Y(n_10877)
);

AOI221xp5_ASAP7_75t_L g10878 ( 
.A1(n_10765),
.A2(n_1316),
.B1(n_1314),
.B2(n_1315),
.C(n_1317),
.Y(n_10878)
);

BUFx3_ASAP7_75t_L g10879 ( 
.A(n_10782),
.Y(n_10879)
);

AND2x4_ASAP7_75t_L g10880 ( 
.A(n_10656),
.B(n_1315),
.Y(n_10880)
);

AND2x2_ASAP7_75t_L g10881 ( 
.A(n_10668),
.B(n_1316),
.Y(n_10881)
);

AO32x2_ASAP7_75t_L g10882 ( 
.A1(n_10502),
.A2(n_1319),
.A3(n_1317),
.B1(n_1318),
.B2(n_1320),
.Y(n_10882)
);

INVx2_ASAP7_75t_L g10883 ( 
.A(n_10511),
.Y(n_10883)
);

AND2x2_ASAP7_75t_L g10884 ( 
.A(n_10630),
.B(n_1318),
.Y(n_10884)
);

OR2x6_ASAP7_75t_L g10885 ( 
.A(n_10732),
.B(n_1321),
.Y(n_10885)
);

HB1xp67_ASAP7_75t_L g10886 ( 
.A(n_10778),
.Y(n_10886)
);

INVx2_ASAP7_75t_L g10887 ( 
.A(n_10712),
.Y(n_10887)
);

BUFx3_ASAP7_75t_L g10888 ( 
.A(n_10507),
.Y(n_10888)
);

AND2x4_ASAP7_75t_L g10889 ( 
.A(n_10713),
.B(n_1321),
.Y(n_10889)
);

AND2x2_ASAP7_75t_L g10890 ( 
.A(n_10716),
.B(n_1322),
.Y(n_10890)
);

A2O1A1Ixp33_ASAP7_75t_L g10891 ( 
.A1(n_10698),
.A2(n_1324),
.B(n_1322),
.C(n_1323),
.Y(n_10891)
);

BUFx12f_ASAP7_75t_L g10892 ( 
.A(n_10556),
.Y(n_10892)
);

AND2x2_ASAP7_75t_L g10893 ( 
.A(n_10524),
.B(n_1324),
.Y(n_10893)
);

AOI22xp33_ASAP7_75t_L g10894 ( 
.A1(n_10764),
.A2(n_1327),
.B1(n_1325),
.B2(n_1326),
.Y(n_10894)
);

AND2x2_ASAP7_75t_L g10895 ( 
.A(n_10528),
.B(n_1325),
.Y(n_10895)
);

INVx1_ASAP7_75t_L g10896 ( 
.A(n_10490),
.Y(n_10896)
);

INVx4_ASAP7_75t_L g10897 ( 
.A(n_10517),
.Y(n_10897)
);

OAI21x1_ASAP7_75t_L g10898 ( 
.A1(n_10629),
.A2(n_1328),
.B(n_1329),
.Y(n_10898)
);

AOI21xp5_ASAP7_75t_L g10899 ( 
.A1(n_10498),
.A2(n_1328),
.B(n_1330),
.Y(n_10899)
);

OAI22xp5_ASAP7_75t_L g10900 ( 
.A1(n_10750),
.A2(n_1333),
.B1(n_1330),
.B2(n_1331),
.Y(n_10900)
);

AND2x2_ASAP7_75t_L g10901 ( 
.A(n_10536),
.B(n_1331),
.Y(n_10901)
);

AND2x4_ASAP7_75t_SL g10902 ( 
.A(n_10748),
.B(n_1333),
.Y(n_10902)
);

INVx1_ASAP7_75t_L g10903 ( 
.A(n_10492),
.Y(n_10903)
);

AND2x2_ASAP7_75t_L g10904 ( 
.A(n_10500),
.B(n_1334),
.Y(n_10904)
);

OAI22xp5_ASAP7_75t_L g10905 ( 
.A1(n_10746),
.A2(n_1337),
.B1(n_1335),
.B2(n_1336),
.Y(n_10905)
);

AND2x2_ASAP7_75t_L g10906 ( 
.A(n_10660),
.B(n_1335),
.Y(n_10906)
);

AND2x4_ASAP7_75t_L g10907 ( 
.A(n_10743),
.B(n_1337),
.Y(n_10907)
);

NAND2xp5_ASAP7_75t_L g10908 ( 
.A(n_10679),
.B(n_1338),
.Y(n_10908)
);

A2O1A1Ixp33_ASAP7_75t_L g10909 ( 
.A1(n_10759),
.A2(n_1341),
.B(n_1339),
.C(n_1340),
.Y(n_10909)
);

CKINVDCx5p33_ASAP7_75t_R g10910 ( 
.A(n_10643),
.Y(n_10910)
);

OAI221xp5_ASAP7_75t_L g10911 ( 
.A1(n_10631),
.A2(n_1341),
.B1(n_1339),
.B2(n_1340),
.C(n_1342),
.Y(n_10911)
);

INVx2_ASAP7_75t_L g10912 ( 
.A(n_10697),
.Y(n_10912)
);

AND2x4_ASAP7_75t_L g10913 ( 
.A(n_10744),
.B(n_1342),
.Y(n_10913)
);

NOR2x1_ASAP7_75t_SL g10914 ( 
.A(n_10573),
.B(n_1343),
.Y(n_10914)
);

NOR2x1_ASAP7_75t_L g10915 ( 
.A(n_10664),
.B(n_1343),
.Y(n_10915)
);

OR2x6_ASAP7_75t_L g10916 ( 
.A(n_10556),
.B(n_1344),
.Y(n_10916)
);

A2O1A1Ixp33_ASAP7_75t_L g10917 ( 
.A1(n_10483),
.A2(n_1347),
.B(n_1344),
.C(n_1345),
.Y(n_10917)
);

OAI21xp5_ASAP7_75t_L g10918 ( 
.A1(n_10560),
.A2(n_1348),
.B(n_1349),
.Y(n_10918)
);

AND2x4_ASAP7_75t_L g10919 ( 
.A(n_10646),
.B(n_1348),
.Y(n_10919)
);

OR2x2_ASAP7_75t_L g10920 ( 
.A(n_10785),
.B(n_1349),
.Y(n_10920)
);

AOI221xp5_ASAP7_75t_L g10921 ( 
.A1(n_10618),
.A2(n_1353),
.B1(n_1351),
.B2(n_1352),
.C(n_1354),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_10495),
.Y(n_10922)
);

NOR2xp33_ASAP7_75t_L g10923 ( 
.A(n_10673),
.B(n_1353),
.Y(n_10923)
);

AND2x2_ASAP7_75t_L g10924 ( 
.A(n_10661),
.B(n_1354),
.Y(n_10924)
);

NAND2xp5_ASAP7_75t_L g10925 ( 
.A(n_10711),
.B(n_1355),
.Y(n_10925)
);

AND2x2_ASAP7_75t_L g10926 ( 
.A(n_10635),
.B(n_1356),
.Y(n_10926)
);

AND2x2_ASAP7_75t_L g10927 ( 
.A(n_10645),
.B(n_1357),
.Y(n_10927)
);

AO21x2_ASAP7_75t_L g10928 ( 
.A1(n_10709),
.A2(n_1357),
.B(n_1359),
.Y(n_10928)
);

AO32x2_ASAP7_75t_L g10929 ( 
.A1(n_10684),
.A2(n_1361),
.A3(n_1359),
.B1(n_1360),
.B2(n_1362),
.Y(n_10929)
);

INVx1_ASAP7_75t_L g10930 ( 
.A(n_10503),
.Y(n_10930)
);

BUFx12f_ASAP7_75t_L g10931 ( 
.A(n_10672),
.Y(n_10931)
);

OR2x2_ASAP7_75t_L g10932 ( 
.A(n_10616),
.B(n_1360),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_10504),
.Y(n_10933)
);

OR2x2_ASAP7_75t_L g10934 ( 
.A(n_10526),
.B(n_1361),
.Y(n_10934)
);

NOR2x1_ASAP7_75t_L g10935 ( 
.A(n_10509),
.B(n_1362),
.Y(n_10935)
);

AND2x4_ASAP7_75t_L g10936 ( 
.A(n_10749),
.B(n_1363),
.Y(n_10936)
);

AND2x2_ASAP7_75t_L g10937 ( 
.A(n_10696),
.B(n_10662),
.Y(n_10937)
);

AND2x2_ASAP7_75t_L g10938 ( 
.A(n_10723),
.B(n_1363),
.Y(n_10938)
);

AO32x2_ASAP7_75t_L g10939 ( 
.A1(n_10600),
.A2(n_10608),
.A3(n_10588),
.B1(n_10567),
.B2(n_10626),
.Y(n_10939)
);

AOI21xp5_ASAP7_75t_L g10940 ( 
.A1(n_10742),
.A2(n_10655),
.B(n_10714),
.Y(n_10940)
);

AOI211xp5_ASAP7_75t_L g10941 ( 
.A1(n_10762),
.A2(n_1366),
.B(n_1364),
.C(n_1365),
.Y(n_10941)
);

INVx3_ASAP7_75t_L g10942 ( 
.A(n_10633),
.Y(n_10942)
);

A2O1A1Ixp33_ASAP7_75t_L g10943 ( 
.A1(n_10767),
.A2(n_1366),
.B(n_1364),
.C(n_1365),
.Y(n_10943)
);

AND2x2_ASAP7_75t_L g10944 ( 
.A(n_10634),
.B(n_1367),
.Y(n_10944)
);

AND2x2_ASAP7_75t_L g10945 ( 
.A(n_10665),
.B(n_10666),
.Y(n_10945)
);

A2O1A1Ixp33_ASAP7_75t_L g10946 ( 
.A1(n_10758),
.A2(n_1370),
.B(n_1368),
.C(n_1369),
.Y(n_10946)
);

AND2x4_ASAP7_75t_L g10947 ( 
.A(n_10641),
.B(n_1368),
.Y(n_10947)
);

OAI21xp5_ASAP7_75t_L g10948 ( 
.A1(n_10625),
.A2(n_10540),
.B(n_10760),
.Y(n_10948)
);

NAND2xp5_ASAP7_75t_L g10949 ( 
.A(n_10728),
.B(n_1370),
.Y(n_10949)
);

AND2x2_ASAP7_75t_L g10950 ( 
.A(n_10647),
.B(n_1371),
.Y(n_10950)
);

NOR2xp33_ASAP7_75t_L g10951 ( 
.A(n_10673),
.B(n_10552),
.Y(n_10951)
);

AND2x2_ASAP7_75t_L g10952 ( 
.A(n_10720),
.B(n_1372),
.Y(n_10952)
);

OR2x2_ASAP7_75t_L g10953 ( 
.A(n_10677),
.B(n_1372),
.Y(n_10953)
);

INVx1_ASAP7_75t_L g10954 ( 
.A(n_10505),
.Y(n_10954)
);

INVx3_ASAP7_75t_L g10955 ( 
.A(n_10633),
.Y(n_10955)
);

AND2x2_ASAP7_75t_L g10956 ( 
.A(n_10721),
.B(n_1373),
.Y(n_10956)
);

AND2x4_ASAP7_75t_L g10957 ( 
.A(n_10717),
.B(n_1373),
.Y(n_10957)
);

AND2x2_ASAP7_75t_L g10958 ( 
.A(n_10752),
.B(n_1374),
.Y(n_10958)
);

NAND2x1p5_ASAP7_75t_L g10959 ( 
.A(n_10649),
.B(n_10705),
.Y(n_10959)
);

INVx1_ASAP7_75t_L g10960 ( 
.A(n_10514),
.Y(n_10960)
);

AND2x2_ASAP7_75t_L g10961 ( 
.A(n_10651),
.B(n_1375),
.Y(n_10961)
);

OA21x2_ASAP7_75t_L g10962 ( 
.A1(n_10537),
.A2(n_1375),
.B(n_1376),
.Y(n_10962)
);

NOR2xp33_ASAP7_75t_L g10963 ( 
.A(n_10586),
.B(n_1376),
.Y(n_10963)
);

O2A1O1Ixp33_ASAP7_75t_SL g10964 ( 
.A1(n_10784),
.A2(n_1379),
.B(n_1377),
.C(n_1378),
.Y(n_10964)
);

BUFx12f_ASAP7_75t_L g10965 ( 
.A(n_10672),
.Y(n_10965)
);

NAND2xp5_ASAP7_75t_L g10966 ( 
.A(n_10735),
.B(n_10671),
.Y(n_10966)
);

AO32x2_ASAP7_75t_L g10967 ( 
.A1(n_10753),
.A2(n_1379),
.A3(n_1377),
.B1(n_1378),
.B2(n_1380),
.Y(n_10967)
);

OAI22xp5_ASAP7_75t_SL g10968 ( 
.A1(n_10506),
.A2(n_1382),
.B1(n_1380),
.B2(n_1381),
.Y(n_10968)
);

INVx2_ASAP7_75t_SL g10969 ( 
.A(n_10572),
.Y(n_10969)
);

NOR2xp33_ASAP7_75t_L g10970 ( 
.A(n_10722),
.B(n_1381),
.Y(n_10970)
);

OAI22xp5_ASAP7_75t_L g10971 ( 
.A1(n_10747),
.A2(n_1384),
.B1(n_1382),
.B2(n_1383),
.Y(n_10971)
);

AND2x4_ASAP7_75t_L g10972 ( 
.A(n_10710),
.B(n_1383),
.Y(n_10972)
);

OA21x2_ASAP7_75t_L g10973 ( 
.A1(n_10636),
.A2(n_1384),
.B(n_1385),
.Y(n_10973)
);

INVx2_ASAP7_75t_L g10974 ( 
.A(n_10722),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_10516),
.Y(n_10975)
);

AND2x2_ASAP7_75t_L g10976 ( 
.A(n_10501),
.B(n_1385),
.Y(n_10976)
);

NOR2x1_ASAP7_75t_SL g10977 ( 
.A(n_10642),
.B(n_1386),
.Y(n_10977)
);

AO32x2_ASAP7_75t_L g10978 ( 
.A1(n_10676),
.A2(n_1388),
.A3(n_1386),
.B1(n_1387),
.B2(n_1389),
.Y(n_10978)
);

OR2x6_ASAP7_75t_L g10979 ( 
.A(n_10751),
.B(n_1387),
.Y(n_10979)
);

NAND4xp25_ASAP7_75t_L g10980 ( 
.A(n_10628),
.B(n_1391),
.C(n_1388),
.D(n_1390),
.Y(n_10980)
);

AND2x4_ASAP7_75t_L g10981 ( 
.A(n_10667),
.B(n_1390),
.Y(n_10981)
);

AO22x2_ASAP7_75t_L g10982 ( 
.A1(n_10708),
.A2(n_1393),
.B1(n_1391),
.B2(n_1392),
.Y(n_10982)
);

NAND2xp5_ASAP7_75t_L g10983 ( 
.A(n_10674),
.B(n_1392),
.Y(n_10983)
);

AND2x2_ASAP7_75t_L g10984 ( 
.A(n_10669),
.B(n_10670),
.Y(n_10984)
);

AND2x2_ASAP7_75t_L g10985 ( 
.A(n_10512),
.B(n_1393),
.Y(n_10985)
);

AND2x2_ASAP7_75t_L g10986 ( 
.A(n_10680),
.B(n_1394),
.Y(n_10986)
);

AND2x2_ASAP7_75t_L g10987 ( 
.A(n_10535),
.B(n_1394),
.Y(n_10987)
);

NOR2x1_ASAP7_75t_SL g10988 ( 
.A(n_10734),
.B(n_1395),
.Y(n_10988)
);

AND2x2_ASAP7_75t_L g10989 ( 
.A(n_10621),
.B(n_10700),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_10519),
.Y(n_10990)
);

A2O1A1Ixp33_ASAP7_75t_L g10991 ( 
.A1(n_10687),
.A2(n_10766),
.B(n_10725),
.C(n_10724),
.Y(n_10991)
);

AND2x4_ASAP7_75t_L g10992 ( 
.A(n_10739),
.B(n_1395),
.Y(n_10992)
);

OAI21xp5_ASAP7_75t_L g10993 ( 
.A1(n_10620),
.A2(n_1396),
.B(n_1397),
.Y(n_10993)
);

INVx1_ASAP7_75t_L g10994 ( 
.A(n_10523),
.Y(n_10994)
);

A2O1A1Ixp33_ASAP7_75t_L g10995 ( 
.A1(n_10681),
.A2(n_1398),
.B(n_1396),
.C(n_1397),
.Y(n_10995)
);

AND2x2_ASAP7_75t_L g10996 ( 
.A(n_10675),
.B(n_1398),
.Y(n_10996)
);

AND2x2_ASAP7_75t_L g10997 ( 
.A(n_10715),
.B(n_1399),
.Y(n_10997)
);

AND2x4_ASAP7_75t_L g10998 ( 
.A(n_10692),
.B(n_1399),
.Y(n_10998)
);

NAND2xp5_ASAP7_75t_L g10999 ( 
.A(n_10733),
.B(n_1400),
.Y(n_10999)
);

BUFx3_ASAP7_75t_L g11000 ( 
.A(n_10730),
.Y(n_11000)
);

OAI22xp5_ASAP7_75t_L g11001 ( 
.A1(n_10521),
.A2(n_1403),
.B1(n_1401),
.B2(n_1402),
.Y(n_11001)
);

NOR2x1_ASAP7_75t_SL g11002 ( 
.A(n_10583),
.B(n_1401),
.Y(n_11002)
);

INVx1_ASAP7_75t_L g11003 ( 
.A(n_10530),
.Y(n_11003)
);

BUFx6f_ASAP7_75t_L g11004 ( 
.A(n_10561),
.Y(n_11004)
);

NOR2xp33_ASAP7_75t_L g11005 ( 
.A(n_10690),
.B(n_10694),
.Y(n_11005)
);

INVx1_ASAP7_75t_L g11006 ( 
.A(n_10531),
.Y(n_11006)
);

NOR2xp33_ASAP7_75t_SL g11007 ( 
.A(n_10768),
.B(n_1404),
.Y(n_11007)
);

INVx1_ASAP7_75t_L g11008 ( 
.A(n_10539),
.Y(n_11008)
);

NOR2xp33_ASAP7_75t_L g11009 ( 
.A(n_10581),
.B(n_1404),
.Y(n_11009)
);

AND2x4_ASAP7_75t_L g11010 ( 
.A(n_10617),
.B(n_1405),
.Y(n_11010)
);

AND2x2_ASAP7_75t_L g11011 ( 
.A(n_10515),
.B(n_1405),
.Y(n_11011)
);

AND2x2_ASAP7_75t_L g11012 ( 
.A(n_10576),
.B(n_1406),
.Y(n_11012)
);

OAI22xp5_ASAP7_75t_L g11013 ( 
.A1(n_10650),
.A2(n_1409),
.B1(n_1407),
.B2(n_1408),
.Y(n_11013)
);

AND2x2_ASAP7_75t_L g11014 ( 
.A(n_10584),
.B(n_1407),
.Y(n_11014)
);

OR2x6_ASAP7_75t_L g11015 ( 
.A(n_10774),
.B(n_1408),
.Y(n_11015)
);

AND2x2_ASAP7_75t_L g11016 ( 
.A(n_10654),
.B(n_1409),
.Y(n_11016)
);

BUFx3_ASAP7_75t_L g11017 ( 
.A(n_10695),
.Y(n_11017)
);

OR2x2_ASAP7_75t_L g11018 ( 
.A(n_10562),
.B(n_1410),
.Y(n_11018)
);

AND2x2_ASAP7_75t_L g11019 ( 
.A(n_10657),
.B(n_1410),
.Y(n_11019)
);

AOI22xp33_ASAP7_75t_L g11020 ( 
.A1(n_10637),
.A2(n_1413),
.B1(n_1411),
.B2(n_1412),
.Y(n_11020)
);

NAND2xp5_ASAP7_75t_L g11021 ( 
.A(n_10527),
.B(n_1411),
.Y(n_11021)
);

AND2x4_ASAP7_75t_L g11022 ( 
.A(n_10685),
.B(n_1414),
.Y(n_11022)
);

AOI21xp5_ASAP7_75t_SL g11023 ( 
.A1(n_10740),
.A2(n_1414),
.B(n_1415),
.Y(n_11023)
);

OAI21xp5_ASAP7_75t_L g11024 ( 
.A1(n_10638),
.A2(n_1415),
.B(n_1416),
.Y(n_11024)
);

INVx2_ASAP7_75t_L g11025 ( 
.A(n_10510),
.Y(n_11025)
);

AND2x2_ASAP7_75t_L g11026 ( 
.A(n_10532),
.B(n_1416),
.Y(n_11026)
);

INVx1_ASAP7_75t_L g11027 ( 
.A(n_10541),
.Y(n_11027)
);

INVx1_ASAP7_75t_L g11028 ( 
.A(n_10543),
.Y(n_11028)
);

AND2x2_ASAP7_75t_L g11029 ( 
.A(n_10533),
.B(n_1417),
.Y(n_11029)
);

AND2x2_ASAP7_75t_L g11030 ( 
.A(n_10538),
.B(n_1417),
.Y(n_11030)
);

AND2x2_ASAP7_75t_L g11031 ( 
.A(n_10542),
.B(n_1418),
.Y(n_11031)
);

OR2x2_ASAP7_75t_L g11032 ( 
.A(n_10558),
.B(n_1418),
.Y(n_11032)
);

NAND2xp5_ASAP7_75t_L g11033 ( 
.A(n_10527),
.B(n_1419),
.Y(n_11033)
);

AND2x2_ASAP7_75t_L g11034 ( 
.A(n_10547),
.B(n_1420),
.Y(n_11034)
);

INVx2_ASAP7_75t_L g11035 ( 
.A(n_10548),
.Y(n_11035)
);

A2O1A1Ixp33_ASAP7_75t_L g11036 ( 
.A1(n_10658),
.A2(n_1423),
.B(n_1421),
.C(n_1422),
.Y(n_11036)
);

NAND2xp5_ASAP7_75t_L g11037 ( 
.A(n_10775),
.B(n_1423),
.Y(n_11037)
);

NAND2xp5_ASAP7_75t_L g11038 ( 
.A(n_10786),
.B(n_1424),
.Y(n_11038)
);

AND2x2_ASAP7_75t_L g11039 ( 
.A(n_10550),
.B(n_1424),
.Y(n_11039)
);

A2O1A1Ixp33_ASAP7_75t_L g11040 ( 
.A1(n_10590),
.A2(n_10787),
.B(n_10795),
.C(n_10737),
.Y(n_11040)
);

AO32x2_ASAP7_75t_L g11041 ( 
.A1(n_10592),
.A2(n_1427),
.A3(n_1425),
.B1(n_1426),
.B2(n_1428),
.Y(n_11041)
);

CKINVDCx20_ASAP7_75t_R g11042 ( 
.A(n_10754),
.Y(n_11042)
);

A2O1A1Ixp33_ASAP7_75t_L g11043 ( 
.A1(n_10624),
.A2(n_1428),
.B(n_1426),
.C(n_1427),
.Y(n_11043)
);

NOR2xp33_ASAP7_75t_SL g11044 ( 
.A(n_10555),
.B(n_1429),
.Y(n_11044)
);

NOR2x1_ASAP7_75t_SL g11045 ( 
.A(n_10704),
.B(n_1429),
.Y(n_11045)
);

AND2x4_ASAP7_75t_L g11046 ( 
.A(n_10559),
.B(n_1430),
.Y(n_11046)
);

OR2x2_ASAP7_75t_L g11047 ( 
.A(n_10563),
.B(n_1430),
.Y(n_11047)
);

OAI22xp5_ASAP7_75t_L g11048 ( 
.A1(n_10545),
.A2(n_1434),
.B1(n_1431),
.B2(n_1432),
.Y(n_11048)
);

INVx2_ASAP7_75t_L g11049 ( 
.A(n_10553),
.Y(n_11049)
);

AND2x2_ASAP7_75t_L g11050 ( 
.A(n_10557),
.B(n_1431),
.Y(n_11050)
);

INVx1_ASAP7_75t_L g11051 ( 
.A(n_10546),
.Y(n_11051)
);

OR2x2_ASAP7_75t_L g11052 ( 
.A(n_10570),
.B(n_1432),
.Y(n_11052)
);

AOI22xp33_ASAP7_75t_L g11053 ( 
.A1(n_10574),
.A2(n_1436),
.B1(n_1434),
.B2(n_1435),
.Y(n_11053)
);

OAI22xp5_ASAP7_75t_L g11054 ( 
.A1(n_10769),
.A2(n_1437),
.B1(n_1435),
.B2(n_1436),
.Y(n_11054)
);

AND2x4_ASAP7_75t_L g11055 ( 
.A(n_10544),
.B(n_1437),
.Y(n_11055)
);

OR2x2_ASAP7_75t_L g11056 ( 
.A(n_10580),
.B(n_1438),
.Y(n_11056)
);

NAND3xp33_ASAP7_75t_L g11057 ( 
.A(n_10615),
.B(n_1438),
.C(n_1439),
.Y(n_11057)
);

OAI21xp5_ASAP7_75t_L g11058 ( 
.A1(n_10736),
.A2(n_1439),
.B(n_1440),
.Y(n_11058)
);

AND2x2_ASAP7_75t_L g11059 ( 
.A(n_10585),
.B(n_1440),
.Y(n_11059)
);

NOR2xp33_ASAP7_75t_L g11060 ( 
.A(n_10755),
.B(n_1441),
.Y(n_11060)
);

AND2x2_ASAP7_75t_L g11061 ( 
.A(n_10589),
.B(n_1442),
.Y(n_11061)
);

NAND2xp5_ASAP7_75t_L g11062 ( 
.A(n_10534),
.B(n_1442),
.Y(n_11062)
);

OA21x2_ASAP7_75t_L g11063 ( 
.A1(n_10575),
.A2(n_1443),
.B(n_1444),
.Y(n_11063)
);

OR2x6_ASAP7_75t_L g11064 ( 
.A(n_10707),
.B(n_1443),
.Y(n_11064)
);

AOI221xp5_ASAP7_75t_L g11065 ( 
.A1(n_10792),
.A2(n_1446),
.B1(n_1444),
.B2(n_1445),
.C(n_1447),
.Y(n_11065)
);

CKINVDCx14_ASAP7_75t_R g11066 ( 
.A(n_10648),
.Y(n_11066)
);

OR2x2_ASAP7_75t_L g11067 ( 
.A(n_10591),
.B(n_1446),
.Y(n_11067)
);

AOI22xp5_ASAP7_75t_L g11068 ( 
.A1(n_10771),
.A2(n_1450),
.B1(n_1447),
.B2(n_1449),
.Y(n_11068)
);

AND2x2_ASAP7_75t_L g11069 ( 
.A(n_10598),
.B(n_1449),
.Y(n_11069)
);

INVx1_ASAP7_75t_L g11070 ( 
.A(n_10777),
.Y(n_11070)
);

OAI21x1_ASAP7_75t_SL g11071 ( 
.A1(n_10780),
.A2(n_1450),
.B(n_1451),
.Y(n_11071)
);

INVx1_ASAP7_75t_L g11072 ( 
.A(n_10789),
.Y(n_11072)
);

A2O1A1Ixp33_ASAP7_75t_L g11073 ( 
.A1(n_10577),
.A2(n_1453),
.B(n_1451),
.C(n_1452),
.Y(n_11073)
);

OAI22xp5_ASAP7_75t_L g11074 ( 
.A1(n_10578),
.A2(n_1456),
.B1(n_1454),
.B2(n_1455),
.Y(n_11074)
);

AND2x4_ASAP7_75t_L g11075 ( 
.A(n_10688),
.B(n_1454),
.Y(n_11075)
);

OR2x2_ASAP7_75t_L g11076 ( 
.A(n_10603),
.B(n_1456),
.Y(n_11076)
);

AND2x2_ASAP7_75t_L g11077 ( 
.A(n_10610),
.B(n_1457),
.Y(n_11077)
);

OA21x2_ASAP7_75t_L g11078 ( 
.A1(n_10579),
.A2(n_10564),
.B(n_10529),
.Y(n_11078)
);

AND2x2_ASAP7_75t_L g11079 ( 
.A(n_10569),
.B(n_1457),
.Y(n_11079)
);

NOR2xp33_ASAP7_75t_L g11080 ( 
.A(n_10587),
.B(n_1458),
.Y(n_11080)
);

AND2x2_ASAP7_75t_L g11081 ( 
.A(n_10571),
.B(n_1458),
.Y(n_11081)
);

INVx1_ASAP7_75t_L g11082 ( 
.A(n_10593),
.Y(n_11082)
);

OR2x2_ASAP7_75t_L g11083 ( 
.A(n_10597),
.B(n_1459),
.Y(n_11083)
);

O2A1O1Ixp33_ASAP7_75t_SL g11084 ( 
.A1(n_10599),
.A2(n_1461),
.B(n_1459),
.C(n_1460),
.Y(n_11084)
);

INVxp67_ASAP7_75t_L g11085 ( 
.A(n_10609),
.Y(n_11085)
);

NOR2xp33_ASAP7_75t_SL g11086 ( 
.A(n_10619),
.B(n_1460),
.Y(n_11086)
);

INVx2_ASAP7_75t_L g11087 ( 
.A(n_10602),
.Y(n_11087)
);

NAND2xp5_ASAP7_75t_L g11088 ( 
.A(n_10703),
.B(n_1461),
.Y(n_11088)
);

NOR2x1_ASAP7_75t_SL g11089 ( 
.A(n_10611),
.B(n_1462),
.Y(n_11089)
);

AND2x2_ASAP7_75t_L g11090 ( 
.A(n_10614),
.B(n_1462),
.Y(n_11090)
);

AND2x4_ASAP7_75t_L g11091 ( 
.A(n_10757),
.B(n_1463),
.Y(n_11091)
);

AND2x4_ASAP7_75t_SL g11092 ( 
.A(n_10757),
.B(n_1463),
.Y(n_11092)
);

INVx1_ASAP7_75t_L g11093 ( 
.A(n_10607),
.Y(n_11093)
);

OA21x2_ASAP7_75t_L g11094 ( 
.A1(n_10594),
.A2(n_1464),
.B(n_1465),
.Y(n_11094)
);

AO21x2_ASAP7_75t_L g11095 ( 
.A1(n_10653),
.A2(n_1464),
.B(n_1465),
.Y(n_11095)
);

A2O1A1Ixp33_ASAP7_75t_L g11096 ( 
.A1(n_10604),
.A2(n_1468),
.B(n_1466),
.C(n_1467),
.Y(n_11096)
);

OAI21x1_ASAP7_75t_SL g11097 ( 
.A1(n_10691),
.A2(n_1466),
.B(n_1468),
.Y(n_11097)
);

AOI22xp5_ASAP7_75t_L g11098 ( 
.A1(n_10484),
.A2(n_1471),
.B1(n_1469),
.B2(n_1470),
.Y(n_11098)
);

AND2x2_ASAP7_75t_L g11099 ( 
.A(n_10582),
.B(n_1469),
.Y(n_11099)
);

NAND2xp5_ASAP7_75t_L g11100 ( 
.A(n_10594),
.B(n_1470),
.Y(n_11100)
);

NAND2xp5_ASAP7_75t_L g11101 ( 
.A(n_10594),
.B(n_1472),
.Y(n_11101)
);

OA21x2_ASAP7_75t_L g11102 ( 
.A1(n_10594),
.A2(n_1473),
.B(n_1474),
.Y(n_11102)
);

INVx1_ASAP7_75t_L g11103 ( 
.A(n_10607),
.Y(n_11103)
);

INVx3_ASAP7_75t_L g11104 ( 
.A(n_10776),
.Y(n_11104)
);

AND2x2_ASAP7_75t_L g11105 ( 
.A(n_10582),
.B(n_1473),
.Y(n_11105)
);

OR2x2_ASAP7_75t_L g11106 ( 
.A(n_10596),
.B(n_1474),
.Y(n_11106)
);

A2O1A1Ixp33_ASAP7_75t_L g11107 ( 
.A1(n_10604),
.A2(n_1477),
.B(n_1475),
.C(n_1476),
.Y(n_11107)
);

NOR2x1_ASAP7_75t_SL g11108 ( 
.A(n_10566),
.B(n_1476),
.Y(n_11108)
);

INVx1_ASAP7_75t_L g11109 ( 
.A(n_10607),
.Y(n_11109)
);

OR2x2_ASAP7_75t_L g11110 ( 
.A(n_10596),
.B(n_1477),
.Y(n_11110)
);

AND2x2_ASAP7_75t_L g11111 ( 
.A(n_10582),
.B(n_1478),
.Y(n_11111)
);

OR2x2_ASAP7_75t_L g11112 ( 
.A(n_10596),
.B(n_1479),
.Y(n_11112)
);

A2O1A1Ixp33_ASAP7_75t_L g11113 ( 
.A1(n_10604),
.A2(n_1481),
.B(n_1479),
.C(n_1480),
.Y(n_11113)
);

AND2x2_ASAP7_75t_L g11114 ( 
.A(n_10582),
.B(n_1480),
.Y(n_11114)
);

NOR2xp33_ASAP7_75t_L g11115 ( 
.A(n_10606),
.B(n_1481),
.Y(n_11115)
);

NOR2xp67_ASAP7_75t_SL g11116 ( 
.A(n_10776),
.B(n_1482),
.Y(n_11116)
);

INVx2_ASAP7_75t_L g11117 ( 
.A(n_10693),
.Y(n_11117)
);

NAND3xp33_ASAP7_75t_L g11118 ( 
.A(n_10653),
.B(n_1482),
.C(n_1484),
.Y(n_11118)
);

NOR3xp33_ASAP7_75t_SL g11119 ( 
.A(n_10793),
.B(n_1485),
.C(n_1486),
.Y(n_11119)
);

AOI22xp5_ASAP7_75t_L g11120 ( 
.A1(n_10484),
.A2(n_1487),
.B1(n_1485),
.B2(n_1486),
.Y(n_11120)
);

AND2x2_ASAP7_75t_L g11121 ( 
.A(n_10582),
.B(n_1488),
.Y(n_11121)
);

AND2x4_ASAP7_75t_L g11122 ( 
.A(n_10491),
.B(n_1489),
.Y(n_11122)
);

AND2x2_ASAP7_75t_L g11123 ( 
.A(n_10582),
.B(n_1489),
.Y(n_11123)
);

AND2x2_ASAP7_75t_L g11124 ( 
.A(n_10582),
.B(n_1490),
.Y(n_11124)
);

BUFx6f_ASAP7_75t_L g11125 ( 
.A(n_10776),
.Y(n_11125)
);

AND2x2_ASAP7_75t_L g11126 ( 
.A(n_10582),
.B(n_1490),
.Y(n_11126)
);

OR2x6_ASAP7_75t_L g11127 ( 
.A(n_10776),
.B(n_1492),
.Y(n_11127)
);

NOR2x1_ASAP7_75t_SL g11128 ( 
.A(n_10566),
.B(n_1492),
.Y(n_11128)
);

AO22x2_ASAP7_75t_L g11129 ( 
.A1(n_10770),
.A2(n_1495),
.B1(n_1493),
.B2(n_1494),
.Y(n_11129)
);

AND2x2_ASAP7_75t_L g11130 ( 
.A(n_10871),
.B(n_1493),
.Y(n_11130)
);

INVx2_ASAP7_75t_L g11131 ( 
.A(n_10888),
.Y(n_11131)
);

BUFx2_ASAP7_75t_L g11132 ( 
.A(n_10892),
.Y(n_11132)
);

AOI22xp33_ASAP7_75t_L g11133 ( 
.A1(n_10815),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_11133)
);

AND2x4_ASAP7_75t_L g11134 ( 
.A(n_10816),
.B(n_1496),
.Y(n_11134)
);

INVxp67_ASAP7_75t_SL g11135 ( 
.A(n_11108),
.Y(n_11135)
);

AND2x2_ASAP7_75t_L g11136 ( 
.A(n_10883),
.B(n_1497),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_L g11137 ( 
.A(n_10874),
.B(n_1497),
.Y(n_11137)
);

NAND2xp5_ASAP7_75t_L g11138 ( 
.A(n_11098),
.B(n_11120),
.Y(n_11138)
);

INVx1_ASAP7_75t_L g11139 ( 
.A(n_10886),
.Y(n_11139)
);

NAND2xp5_ASAP7_75t_L g11140 ( 
.A(n_10839),
.B(n_1499),
.Y(n_11140)
);

INVx1_ASAP7_75t_L g11141 ( 
.A(n_10803),
.Y(n_11141)
);

INVx2_ASAP7_75t_L g11142 ( 
.A(n_10840),
.Y(n_11142)
);

AND2x4_ASAP7_75t_L g11143 ( 
.A(n_11104),
.B(n_1499),
.Y(n_11143)
);

BUFx2_ASAP7_75t_L g11144 ( 
.A(n_10841),
.Y(n_11144)
);

INVx2_ASAP7_75t_L g11145 ( 
.A(n_10879),
.Y(n_11145)
);

AND2x2_ASAP7_75t_L g11146 ( 
.A(n_10851),
.B(n_1500),
.Y(n_11146)
);

OR2x2_ASAP7_75t_L g11147 ( 
.A(n_10800),
.B(n_1500),
.Y(n_11147)
);

OR2x2_ASAP7_75t_L g11148 ( 
.A(n_10807),
.B(n_1501),
.Y(n_11148)
);

AND2x2_ASAP7_75t_L g11149 ( 
.A(n_10833),
.B(n_1501),
.Y(n_11149)
);

INVx1_ASAP7_75t_L g11150 ( 
.A(n_10806),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_10809),
.Y(n_11151)
);

AND2x2_ASAP7_75t_L g11152 ( 
.A(n_11117),
.B(n_1502),
.Y(n_11152)
);

OR2x2_ASAP7_75t_L g11153 ( 
.A(n_10797),
.B(n_1502),
.Y(n_11153)
);

INVx1_ASAP7_75t_L g11154 ( 
.A(n_10810),
.Y(n_11154)
);

INVx1_ASAP7_75t_L g11155 ( 
.A(n_10822),
.Y(n_11155)
);

AND2x2_ASAP7_75t_L g11156 ( 
.A(n_10863),
.B(n_1503),
.Y(n_11156)
);

INVx1_ASAP7_75t_L g11157 ( 
.A(n_10857),
.Y(n_11157)
);

OAI22xp5_ASAP7_75t_L g11158 ( 
.A1(n_10917),
.A2(n_1505),
.B1(n_1503),
.B2(n_1504),
.Y(n_11158)
);

INVx2_ASAP7_75t_L g11159 ( 
.A(n_10942),
.Y(n_11159)
);

OR2x2_ASAP7_75t_L g11160 ( 
.A(n_11093),
.B(n_11103),
.Y(n_11160)
);

INVx1_ASAP7_75t_L g11161 ( 
.A(n_10896),
.Y(n_11161)
);

INVx1_ASAP7_75t_L g11162 ( 
.A(n_10903),
.Y(n_11162)
);

INVx1_ASAP7_75t_L g11163 ( 
.A(n_10922),
.Y(n_11163)
);

NOR2x1_ASAP7_75t_L g11164 ( 
.A(n_10915),
.B(n_1504),
.Y(n_11164)
);

INVx2_ASAP7_75t_L g11165 ( 
.A(n_10955),
.Y(n_11165)
);

INVx1_ASAP7_75t_L g11166 ( 
.A(n_10930),
.Y(n_11166)
);

INVx1_ASAP7_75t_L g11167 ( 
.A(n_10933),
.Y(n_11167)
);

OR2x2_ASAP7_75t_L g11168 ( 
.A(n_11109),
.B(n_1506),
.Y(n_11168)
);

AND2x2_ASAP7_75t_L g11169 ( 
.A(n_10969),
.B(n_1507),
.Y(n_11169)
);

INVx3_ASAP7_75t_L g11170 ( 
.A(n_10931),
.Y(n_11170)
);

INVx1_ASAP7_75t_L g11171 ( 
.A(n_10954),
.Y(n_11171)
);

INVx2_ASAP7_75t_L g11172 ( 
.A(n_10828),
.Y(n_11172)
);

OR2x6_ASAP7_75t_L g11173 ( 
.A(n_11125),
.B(n_1507),
.Y(n_11173)
);

AND2x2_ASAP7_75t_L g11174 ( 
.A(n_10861),
.B(n_1508),
.Y(n_11174)
);

AND2x2_ASAP7_75t_L g11175 ( 
.A(n_10951),
.B(n_1508),
.Y(n_11175)
);

AND2x2_ASAP7_75t_L g11176 ( 
.A(n_10856),
.B(n_1510),
.Y(n_11176)
);

NAND2xp5_ASAP7_75t_L g11177 ( 
.A(n_10860),
.B(n_1510),
.Y(n_11177)
);

OR2x2_ASAP7_75t_L g11178 ( 
.A(n_10887),
.B(n_10966),
.Y(n_11178)
);

AND2x2_ASAP7_75t_L g11179 ( 
.A(n_10845),
.B(n_1511),
.Y(n_11179)
);

AND2x2_ASAP7_75t_L g11180 ( 
.A(n_10974),
.B(n_1511),
.Y(n_11180)
);

INVx1_ASAP7_75t_SL g11181 ( 
.A(n_11042),
.Y(n_11181)
);

INVx2_ASAP7_75t_L g11182 ( 
.A(n_10828),
.Y(n_11182)
);

NOR2x1_ASAP7_75t_SL g11183 ( 
.A(n_11095),
.B(n_1512),
.Y(n_11183)
);

INVx2_ASAP7_75t_L g11184 ( 
.A(n_10870),
.Y(n_11184)
);

OR2x2_ASAP7_75t_L g11185 ( 
.A(n_10873),
.B(n_1513),
.Y(n_11185)
);

AND2x2_ASAP7_75t_L g11186 ( 
.A(n_10912),
.B(n_1513),
.Y(n_11186)
);

AND2x2_ASAP7_75t_L g11187 ( 
.A(n_11085),
.B(n_1514),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_10870),
.Y(n_11188)
);

HB1xp67_ASAP7_75t_L g11189 ( 
.A(n_11078),
.Y(n_11189)
);

NOR2xp33_ASAP7_75t_L g11190 ( 
.A(n_11125),
.B(n_1514),
.Y(n_11190)
);

BUFx3_ASAP7_75t_L g11191 ( 
.A(n_10808),
.Y(n_11191)
);

INVx1_ASAP7_75t_L g11192 ( 
.A(n_10960),
.Y(n_11192)
);

OR2x2_ASAP7_75t_L g11193 ( 
.A(n_10859),
.B(n_1515),
.Y(n_11193)
);

AND2x2_ASAP7_75t_L g11194 ( 
.A(n_11066),
.B(n_1516),
.Y(n_11194)
);

INVx1_ASAP7_75t_L g11195 ( 
.A(n_10975),
.Y(n_11195)
);

HB1xp67_ASAP7_75t_L g11196 ( 
.A(n_10962),
.Y(n_11196)
);

AOI22xp33_ASAP7_75t_L g11197 ( 
.A1(n_10899),
.A2(n_1520),
.B1(n_1518),
.B2(n_1519),
.Y(n_11197)
);

AND2x4_ASAP7_75t_SL g11198 ( 
.A(n_10866),
.B(n_1518),
.Y(n_11198)
);

AND2x2_ASAP7_75t_L g11199 ( 
.A(n_10811),
.B(n_10843),
.Y(n_11199)
);

INVx1_ASAP7_75t_L g11200 ( 
.A(n_10990),
.Y(n_11200)
);

AND2x2_ASAP7_75t_L g11201 ( 
.A(n_10897),
.B(n_1519),
.Y(n_11201)
);

INVx2_ASAP7_75t_L g11202 ( 
.A(n_11000),
.Y(n_11202)
);

BUFx2_ASAP7_75t_L g11203 ( 
.A(n_10939),
.Y(n_11203)
);

INVx1_ASAP7_75t_L g11204 ( 
.A(n_10994),
.Y(n_11204)
);

INVx2_ASAP7_75t_L g11205 ( 
.A(n_11004),
.Y(n_11205)
);

BUFx6f_ASAP7_75t_L g11206 ( 
.A(n_10965),
.Y(n_11206)
);

AOI22xp33_ASAP7_75t_L g11207 ( 
.A1(n_10821),
.A2(n_1523),
.B1(n_1520),
.B2(n_1521),
.Y(n_11207)
);

AND2x2_ASAP7_75t_L g11208 ( 
.A(n_10937),
.B(n_1521),
.Y(n_11208)
);

INVx1_ASAP7_75t_L g11209 ( 
.A(n_11003),
.Y(n_11209)
);

AND2x2_ASAP7_75t_L g11210 ( 
.A(n_10976),
.B(n_1524),
.Y(n_11210)
);

BUFx12f_ASAP7_75t_L g11211 ( 
.A(n_11127),
.Y(n_11211)
);

INVx3_ASAP7_75t_L g11212 ( 
.A(n_11004),
.Y(n_11212)
);

AND2x2_ASAP7_75t_SL g11213 ( 
.A(n_11092),
.B(n_1524),
.Y(n_11213)
);

NOR2xp33_ASAP7_75t_L g11214 ( 
.A(n_10837),
.B(n_1525),
.Y(n_11214)
);

AND2x2_ASAP7_75t_L g11215 ( 
.A(n_11017),
.B(n_10945),
.Y(n_11215)
);

INVx2_ASAP7_75t_L g11216 ( 
.A(n_11128),
.Y(n_11216)
);

AND2x2_ASAP7_75t_L g11217 ( 
.A(n_10959),
.B(n_1525),
.Y(n_11217)
);

AND2x4_ASAP7_75t_L g11218 ( 
.A(n_10812),
.B(n_1526),
.Y(n_11218)
);

BUFx2_ASAP7_75t_L g11219 ( 
.A(n_10939),
.Y(n_11219)
);

AND2x4_ASAP7_75t_L g11220 ( 
.A(n_11122),
.B(n_1526),
.Y(n_11220)
);

OR2x2_ASAP7_75t_L g11221 ( 
.A(n_10829),
.B(n_1527),
.Y(n_11221)
);

OR2x2_ASAP7_75t_L g11222 ( 
.A(n_11025),
.B(n_1527),
.Y(n_11222)
);

AND2x2_ASAP7_75t_L g11223 ( 
.A(n_10865),
.B(n_10989),
.Y(n_11223)
);

INVx2_ASAP7_75t_L g11224 ( 
.A(n_11089),
.Y(n_11224)
);

NAND2xp5_ASAP7_75t_L g11225 ( 
.A(n_10823),
.B(n_1528),
.Y(n_11225)
);

INVx3_ASAP7_75t_L g11226 ( 
.A(n_10910),
.Y(n_11226)
);

INVx5_ASAP7_75t_L g11227 ( 
.A(n_11127),
.Y(n_11227)
);

OR2x2_ASAP7_75t_L g11228 ( 
.A(n_11035),
.B(n_11049),
.Y(n_11228)
);

INVx1_ASAP7_75t_SL g11229 ( 
.A(n_10916),
.Y(n_11229)
);

HB1xp67_ASAP7_75t_L g11230 ( 
.A(n_10973),
.Y(n_11230)
);

INVxp67_ASAP7_75t_SL g11231 ( 
.A(n_10850),
.Y(n_11231)
);

INVx1_ASAP7_75t_L g11232 ( 
.A(n_11006),
.Y(n_11232)
);

BUFx2_ASAP7_75t_L g11233 ( 
.A(n_10835),
.Y(n_11233)
);

INVx2_ASAP7_75t_L g11234 ( 
.A(n_11032),
.Y(n_11234)
);

OR2x2_ASAP7_75t_L g11235 ( 
.A(n_10832),
.B(n_1528),
.Y(n_11235)
);

HB1xp67_ASAP7_75t_L g11236 ( 
.A(n_10846),
.Y(n_11236)
);

INVx1_ASAP7_75t_L g11237 ( 
.A(n_11008),
.Y(n_11237)
);

INVx2_ASAP7_75t_L g11238 ( 
.A(n_11047),
.Y(n_11238)
);

HB1xp67_ASAP7_75t_L g11239 ( 
.A(n_11094),
.Y(n_11239)
);

OAI21xp5_ASAP7_75t_L g11240 ( 
.A1(n_10827),
.A2(n_1529),
.B(n_1530),
.Y(n_11240)
);

AND2x2_ASAP7_75t_L g11241 ( 
.A(n_11040),
.B(n_1530),
.Y(n_11241)
);

AND2x2_ASAP7_75t_L g11242 ( 
.A(n_10938),
.B(n_1531),
.Y(n_11242)
);

NOR2xp33_ASAP7_75t_L g11243 ( 
.A(n_10804),
.B(n_1532),
.Y(n_11243)
);

INVx1_ASAP7_75t_L g11244 ( 
.A(n_11027),
.Y(n_11244)
);

OR2x2_ASAP7_75t_L g11245 ( 
.A(n_10949),
.B(n_1532),
.Y(n_11245)
);

INVx2_ASAP7_75t_L g11246 ( 
.A(n_11052),
.Y(n_11246)
);

AND2x2_ASAP7_75t_L g11247 ( 
.A(n_10950),
.B(n_1533),
.Y(n_11247)
);

INVx2_ASAP7_75t_L g11248 ( 
.A(n_11056),
.Y(n_11248)
);

INVx2_ASAP7_75t_SL g11249 ( 
.A(n_10817),
.Y(n_11249)
);

INVx2_ASAP7_75t_L g11250 ( 
.A(n_11067),
.Y(n_11250)
);

INVx2_ASAP7_75t_L g11251 ( 
.A(n_11076),
.Y(n_11251)
);

AND2x2_ASAP7_75t_L g11252 ( 
.A(n_10944),
.B(n_1534),
.Y(n_11252)
);

AND2x2_ASAP7_75t_L g11253 ( 
.A(n_10958),
.B(n_10997),
.Y(n_11253)
);

OR2x2_ASAP7_75t_L g11254 ( 
.A(n_10908),
.B(n_1535),
.Y(n_11254)
);

INVx1_ASAP7_75t_L g11255 ( 
.A(n_11028),
.Y(n_11255)
);

INVx2_ASAP7_75t_SL g11256 ( 
.A(n_10853),
.Y(n_11256)
);

INVx2_ASAP7_75t_L g11257 ( 
.A(n_11002),
.Y(n_11257)
);

INVx1_ASAP7_75t_L g11258 ( 
.A(n_11051),
.Y(n_11258)
);

AND2x2_ASAP7_75t_L g11259 ( 
.A(n_11005),
.B(n_1535),
.Y(n_11259)
);

INVx2_ASAP7_75t_L g11260 ( 
.A(n_11083),
.Y(n_11260)
);

AND2x2_ASAP7_75t_L g11261 ( 
.A(n_10825),
.B(n_1536),
.Y(n_11261)
);

AND2x2_ASAP7_75t_L g11262 ( 
.A(n_10831),
.B(n_1536),
.Y(n_11262)
);

OAI33xp33_ASAP7_75t_L g11263 ( 
.A1(n_10968),
.A2(n_1540),
.A3(n_1542),
.B1(n_1538),
.B2(n_1539),
.B3(n_1541),
.Y(n_11263)
);

OR2x2_ASAP7_75t_L g11264 ( 
.A(n_10801),
.B(n_1539),
.Y(n_11264)
);

INVx2_ASAP7_75t_L g11265 ( 
.A(n_10984),
.Y(n_11265)
);

AND2x2_ASAP7_75t_L g11266 ( 
.A(n_10836),
.B(n_1540),
.Y(n_11266)
);

AO31x2_ASAP7_75t_L g11267 ( 
.A1(n_11100),
.A2(n_11101),
.A3(n_10914),
.B(n_10977),
.Y(n_11267)
);

INVx1_ASAP7_75t_L g11268 ( 
.A(n_11070),
.Y(n_11268)
);

INVx2_ASAP7_75t_L g11269 ( 
.A(n_11018),
.Y(n_11269)
);

AND2x2_ASAP7_75t_L g11270 ( 
.A(n_10802),
.B(n_1541),
.Y(n_11270)
);

INVx1_ASAP7_75t_L g11271 ( 
.A(n_11072),
.Y(n_11271)
);

BUFx3_ASAP7_75t_L g11272 ( 
.A(n_10902),
.Y(n_11272)
);

NOR2xp33_ASAP7_75t_L g11273 ( 
.A(n_10796),
.B(n_1542),
.Y(n_11273)
);

AO21x2_ASAP7_75t_L g11274 ( 
.A1(n_10948),
.A2(n_1543),
.B(n_1545),
.Y(n_11274)
);

AOI21xp5_ASAP7_75t_L g11275 ( 
.A1(n_10988),
.A2(n_1543),
.B(n_1545),
.Y(n_11275)
);

INVx1_ASAP7_75t_L g11276 ( 
.A(n_11087),
.Y(n_11276)
);

AND2x2_ASAP7_75t_L g11277 ( 
.A(n_10991),
.B(n_1546),
.Y(n_11277)
);

OR2x2_ASAP7_75t_L g11278 ( 
.A(n_10932),
.B(n_1547),
.Y(n_11278)
);

AND2x2_ASAP7_75t_L g11279 ( 
.A(n_10799),
.B(n_1547),
.Y(n_11279)
);

OR2x2_ASAP7_75t_L g11280 ( 
.A(n_10925),
.B(n_1548),
.Y(n_11280)
);

HB1xp67_ASAP7_75t_L g11281 ( 
.A(n_11102),
.Y(n_11281)
);

INVx2_ASAP7_75t_L g11282 ( 
.A(n_10986),
.Y(n_11282)
);

INVx2_ASAP7_75t_L g11283 ( 
.A(n_11079),
.Y(n_11283)
);

INVx2_ASAP7_75t_L g11284 ( 
.A(n_11081),
.Y(n_11284)
);

INVx2_ASAP7_75t_L g11285 ( 
.A(n_11090),
.Y(n_11285)
);

OR2x2_ASAP7_75t_L g11286 ( 
.A(n_10983),
.B(n_1549),
.Y(n_11286)
);

AND2x2_ASAP7_75t_L g11287 ( 
.A(n_11099),
.B(n_1549),
.Y(n_11287)
);

CKINVDCx11_ASAP7_75t_R g11288 ( 
.A(n_10916),
.Y(n_11288)
);

AND2x4_ASAP7_75t_L g11289 ( 
.A(n_10844),
.B(n_1550),
.Y(n_11289)
);

AOI221xp5_ASAP7_75t_L g11290 ( 
.A1(n_10824),
.A2(n_1552),
.B1(n_1550),
.B2(n_1551),
.C(n_1553),
.Y(n_11290)
);

OR2x2_ASAP7_75t_L g11291 ( 
.A(n_10953),
.B(n_1551),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_11082),
.Y(n_11292)
);

INVxp67_ASAP7_75t_SL g11293 ( 
.A(n_10820),
.Y(n_11293)
);

INVx2_ASAP7_75t_L g11294 ( 
.A(n_11026),
.Y(n_11294)
);

INVx5_ASAP7_75t_SL g11295 ( 
.A(n_10885),
.Y(n_11295)
);

INVx5_ASAP7_75t_SL g11296 ( 
.A(n_10885),
.Y(n_11296)
);

AOI22xp33_ASAP7_75t_L g11297 ( 
.A1(n_10814),
.A2(n_1556),
.B1(n_1554),
.B2(n_1555),
.Y(n_11297)
);

INVx1_ASAP7_75t_L g11298 ( 
.A(n_11029),
.Y(n_11298)
);

INVx2_ASAP7_75t_L g11299 ( 
.A(n_11030),
.Y(n_11299)
);

AND2x2_ASAP7_75t_L g11300 ( 
.A(n_11105),
.B(n_1555),
.Y(n_11300)
);

INVx2_ASAP7_75t_L g11301 ( 
.A(n_11031),
.Y(n_11301)
);

INVx4_ASAP7_75t_L g11302 ( 
.A(n_10880),
.Y(n_11302)
);

INVx1_ASAP7_75t_L g11303 ( 
.A(n_11034),
.Y(n_11303)
);

INVx2_ASAP7_75t_SL g11304 ( 
.A(n_10830),
.Y(n_11304)
);

INVx1_ASAP7_75t_L g11305 ( 
.A(n_11039),
.Y(n_11305)
);

INVx1_ASAP7_75t_L g11306 ( 
.A(n_11050),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_11111),
.B(n_1556),
.Y(n_11307)
);

INVx2_ASAP7_75t_L g11308 ( 
.A(n_11059),
.Y(n_11308)
);

INVx3_ASAP7_75t_L g11309 ( 
.A(n_10813),
.Y(n_11309)
);

INVx2_ASAP7_75t_L g11310 ( 
.A(n_11061),
.Y(n_11310)
);

INVx2_ASAP7_75t_L g11311 ( 
.A(n_11069),
.Y(n_11311)
);

NOR2x1_ASAP7_75t_R g11312 ( 
.A(n_10936),
.B(n_1557),
.Y(n_11312)
);

AND2x2_ASAP7_75t_L g11313 ( 
.A(n_11114),
.B(n_1557),
.Y(n_11313)
);

AND2x2_ASAP7_75t_L g11314 ( 
.A(n_11121),
.B(n_1558),
.Y(n_11314)
);

NAND2xp5_ASAP7_75t_L g11315 ( 
.A(n_10940),
.B(n_1558),
.Y(n_11315)
);

INVx1_ASAP7_75t_L g11316 ( 
.A(n_11077),
.Y(n_11316)
);

INVx2_ASAP7_75t_L g11317 ( 
.A(n_10985),
.Y(n_11317)
);

INVx2_ASAP7_75t_L g11318 ( 
.A(n_10987),
.Y(n_11318)
);

AND2x2_ASAP7_75t_L g11319 ( 
.A(n_11123),
.B(n_1559),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_10934),
.Y(n_11320)
);

INVx2_ASAP7_75t_L g11321 ( 
.A(n_11097),
.Y(n_11321)
);

INVx2_ASAP7_75t_SL g11322 ( 
.A(n_10889),
.Y(n_11322)
);

AND2x2_ASAP7_75t_L g11323 ( 
.A(n_11124),
.B(n_1559),
.Y(n_11323)
);

INVx2_ASAP7_75t_L g11324 ( 
.A(n_10961),
.Y(n_11324)
);

INVxp67_ASAP7_75t_L g11325 ( 
.A(n_10847),
.Y(n_11325)
);

BUFx2_ASAP7_75t_L g11326 ( 
.A(n_10835),
.Y(n_11326)
);

AND2x2_ASAP7_75t_L g11327 ( 
.A(n_11126),
.B(n_1560),
.Y(n_11327)
);

INVx3_ASAP7_75t_L g11328 ( 
.A(n_10972),
.Y(n_11328)
);

AND2x2_ASAP7_75t_L g11329 ( 
.A(n_10924),
.B(n_1560),
.Y(n_11329)
);

AND2x2_ASAP7_75t_L g11330 ( 
.A(n_10881),
.B(n_1563),
.Y(n_11330)
);

INVxp67_ASAP7_75t_SL g11331 ( 
.A(n_11045),
.Y(n_11331)
);

INVx2_ASAP7_75t_L g11332 ( 
.A(n_10872),
.Y(n_11332)
);

OR2x2_ASAP7_75t_L g11333 ( 
.A(n_11106),
.B(n_1563),
.Y(n_11333)
);

INVx1_ASAP7_75t_L g11334 ( 
.A(n_11063),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_L g11335 ( 
.A(n_11091),
.B(n_1564),
.Y(n_11335)
);

INVx1_ASAP7_75t_L g11336 ( 
.A(n_10920),
.Y(n_11336)
);

OR2x2_ASAP7_75t_L g11337 ( 
.A(n_11110),
.B(n_11112),
.Y(n_11337)
);

AND2x2_ASAP7_75t_L g11338 ( 
.A(n_10858),
.B(n_1564),
.Y(n_11338)
);

INVx1_ASAP7_75t_L g11339 ( 
.A(n_10884),
.Y(n_11339)
);

AND2x2_ASAP7_75t_L g11340 ( 
.A(n_10864),
.B(n_1565),
.Y(n_11340)
);

INVxp67_ASAP7_75t_SL g11341 ( 
.A(n_10935),
.Y(n_11341)
);

BUFx2_ASAP7_75t_L g11342 ( 
.A(n_11064),
.Y(n_11342)
);

OR2x2_ASAP7_75t_L g11343 ( 
.A(n_10906),
.B(n_1565),
.Y(n_11343)
);

INVx2_ASAP7_75t_L g11344 ( 
.A(n_10893),
.Y(n_11344)
);

NAND2xp5_ASAP7_75t_L g11345 ( 
.A(n_11129),
.B(n_1566),
.Y(n_11345)
);

INVx1_ASAP7_75t_L g11346 ( 
.A(n_10895),
.Y(n_11346)
);

HB1xp67_ASAP7_75t_L g11347 ( 
.A(n_10928),
.Y(n_11347)
);

AND2x2_ASAP7_75t_L g11348 ( 
.A(n_11064),
.B(n_1566),
.Y(n_11348)
);

INVx2_ASAP7_75t_L g11349 ( 
.A(n_10901),
.Y(n_11349)
);

AND2x4_ASAP7_75t_L g11350 ( 
.A(n_10848),
.B(n_10890),
.Y(n_11350)
);

INVx2_ASAP7_75t_L g11351 ( 
.A(n_11010),
.Y(n_11351)
);

HB1xp67_ASAP7_75t_L g11352 ( 
.A(n_11015),
.Y(n_11352)
);

INVx2_ASAP7_75t_L g11353 ( 
.A(n_10981),
.Y(n_11353)
);

AND2x2_ASAP7_75t_L g11354 ( 
.A(n_10926),
.B(n_1567),
.Y(n_11354)
);

INVx2_ASAP7_75t_L g11355 ( 
.A(n_10919),
.Y(n_11355)
);

AOI22xp5_ASAP7_75t_L g11356 ( 
.A1(n_11119),
.A2(n_1570),
.B1(n_1568),
.B2(n_1569),
.Y(n_11356)
);

BUFx2_ASAP7_75t_L g11357 ( 
.A(n_11015),
.Y(n_11357)
);

BUFx2_ASAP7_75t_L g11358 ( 
.A(n_10979),
.Y(n_11358)
);

AND2x2_ASAP7_75t_L g11359 ( 
.A(n_10927),
.B(n_1569),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_11016),
.Y(n_11360)
);

INVx2_ASAP7_75t_L g11361 ( 
.A(n_10996),
.Y(n_11361)
);

INVx2_ASAP7_75t_L g11362 ( 
.A(n_11019),
.Y(n_11362)
);

INVx1_ASAP7_75t_L g11363 ( 
.A(n_10952),
.Y(n_11363)
);

HB1xp67_ASAP7_75t_L g11364 ( 
.A(n_10898),
.Y(n_11364)
);

INVx1_ASAP7_75t_L g11365 ( 
.A(n_10956),
.Y(n_11365)
);

AO21x2_ASAP7_75t_L g11366 ( 
.A1(n_10862),
.A2(n_1570),
.B(n_1571),
.Y(n_11366)
);

NAND2xp5_ASAP7_75t_L g11367 ( 
.A(n_11009),
.B(n_1571),
.Y(n_11367)
);

AND2x2_ASAP7_75t_L g11368 ( 
.A(n_11011),
.B(n_1572),
.Y(n_11368)
);

AND2x2_ASAP7_75t_L g11369 ( 
.A(n_10904),
.B(n_1572),
.Y(n_11369)
);

AND2x2_ASAP7_75t_L g11370 ( 
.A(n_11012),
.B(n_1573),
.Y(n_11370)
);

AND2x2_ASAP7_75t_L g11371 ( 
.A(n_11014),
.B(n_1573),
.Y(n_11371)
);

CKINVDCx16_ASAP7_75t_R g11372 ( 
.A(n_11007),
.Y(n_11372)
);

NAND2xp5_ASAP7_75t_L g11373 ( 
.A(n_10869),
.B(n_1574),
.Y(n_11373)
);

NAND2xp5_ASAP7_75t_L g11374 ( 
.A(n_10826),
.B(n_1574),
.Y(n_11374)
);

NAND2xp5_ASAP7_75t_L g11375 ( 
.A(n_10957),
.B(n_10982),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_10978),
.Y(n_11376)
);

BUFx2_ASAP7_75t_L g11377 ( 
.A(n_10979),
.Y(n_11377)
);

NAND2xp5_ASAP7_75t_L g11378 ( 
.A(n_10999),
.B(n_1575),
.Y(n_11378)
);

INVx1_ASAP7_75t_L g11379 ( 
.A(n_10978),
.Y(n_11379)
);

NAND3xp33_ASAP7_75t_L g11380 ( 
.A(n_11240),
.B(n_10818),
.C(n_10798),
.Y(n_11380)
);

NAND3xp33_ASAP7_75t_L g11381 ( 
.A(n_11347),
.B(n_11107),
.C(n_11096),
.Y(n_11381)
);

OAI21xp5_ASAP7_75t_SL g11382 ( 
.A1(n_11233),
.A2(n_11113),
.B(n_10819),
.Y(n_11382)
);

NAND2xp5_ASAP7_75t_L g11383 ( 
.A(n_11326),
.B(n_10923),
.Y(n_11383)
);

NAND3xp33_ASAP7_75t_L g11384 ( 
.A(n_11203),
.B(n_10941),
.C(n_10921),
.Y(n_11384)
);

NAND2xp5_ASAP7_75t_L g11385 ( 
.A(n_11229),
.B(n_10868),
.Y(n_11385)
);

AND2x2_ASAP7_75t_L g11386 ( 
.A(n_11132),
.B(n_11115),
.Y(n_11386)
);

NAND2xp5_ASAP7_75t_L g11387 ( 
.A(n_11376),
.B(n_11021),
.Y(n_11387)
);

NAND2xp5_ASAP7_75t_L g11388 ( 
.A(n_11379),
.B(n_11033),
.Y(n_11388)
);

NAND2xp5_ASAP7_75t_L g11389 ( 
.A(n_11293),
.B(n_11080),
.Y(n_11389)
);

AND2x2_ASAP7_75t_L g11390 ( 
.A(n_11295),
.B(n_10834),
.Y(n_11390)
);

NOR2xp33_ASAP7_75t_SL g11391 ( 
.A(n_11227),
.B(n_11116),
.Y(n_11391)
);

AND2x2_ASAP7_75t_L g11392 ( 
.A(n_11295),
.B(n_11046),
.Y(n_11392)
);

NAND2xp5_ASAP7_75t_L g11393 ( 
.A(n_11341),
.B(n_10943),
.Y(n_11393)
);

NAND3xp33_ASAP7_75t_L g11394 ( 
.A(n_11219),
.B(n_11230),
.C(n_11236),
.Y(n_11394)
);

AND2x2_ASAP7_75t_L g11395 ( 
.A(n_11296),
.B(n_11075),
.Y(n_11395)
);

AOI22xp5_ASAP7_75t_L g11396 ( 
.A1(n_11372),
.A2(n_10878),
.B1(n_10805),
.B2(n_10980),
.Y(n_11396)
);

NAND2xp5_ASAP7_75t_SL g11397 ( 
.A(n_11227),
.B(n_10993),
.Y(n_11397)
);

NOR2xp33_ASAP7_75t_L g11398 ( 
.A(n_11206),
.B(n_11086),
.Y(n_11398)
);

OAI21xp5_ASAP7_75t_SL g11399 ( 
.A1(n_11138),
.A2(n_10891),
.B(n_10894),
.Y(n_11399)
);

NAND2xp5_ASAP7_75t_L g11400 ( 
.A(n_11181),
.B(n_10875),
.Y(n_11400)
);

NAND3xp33_ASAP7_75t_L g11401 ( 
.A(n_11334),
.B(n_10854),
.C(n_11065),
.Y(n_11401)
);

NAND2xp5_ASAP7_75t_L g11402 ( 
.A(n_11357),
.B(n_10907),
.Y(n_11402)
);

NAND2xp5_ASAP7_75t_L g11403 ( 
.A(n_11352),
.B(n_10992),
.Y(n_11403)
);

AOI22xp33_ASAP7_75t_SL g11404 ( 
.A1(n_11231),
.A2(n_10867),
.B1(n_11118),
.B2(n_11057),
.Y(n_11404)
);

NAND3xp33_ASAP7_75t_L g11405 ( 
.A(n_11239),
.B(n_11020),
.C(n_10852),
.Y(n_11405)
);

OA211x2_ASAP7_75t_L g11406 ( 
.A1(n_11325),
.A2(n_11044),
.B(n_11058),
.C(n_10918),
.Y(n_11406)
);

NAND3xp33_ASAP7_75t_L g11407 ( 
.A(n_11281),
.B(n_11196),
.C(n_11189),
.Y(n_11407)
);

OAI21xp5_ASAP7_75t_SL g11408 ( 
.A1(n_11356),
.A2(n_10877),
.B(n_10876),
.Y(n_11408)
);

NAND3xp33_ASAP7_75t_L g11409 ( 
.A(n_11164),
.B(n_10946),
.C(n_11073),
.Y(n_11409)
);

NAND2xp5_ASAP7_75t_L g11410 ( 
.A(n_11135),
.B(n_10998),
.Y(n_11410)
);

OAI21xp5_ASAP7_75t_SL g11411 ( 
.A1(n_11241),
.A2(n_11068),
.B(n_10911),
.Y(n_11411)
);

NAND2xp5_ASAP7_75t_L g11412 ( 
.A(n_11342),
.B(n_11036),
.Y(n_11412)
);

OAI221xp5_ASAP7_75t_L g11413 ( 
.A1(n_11331),
.A2(n_11043),
.B1(n_11024),
.B2(n_10909),
.C(n_10905),
.Y(n_11413)
);

NAND2xp5_ASAP7_75t_SL g11414 ( 
.A(n_11257),
.B(n_10947),
.Y(n_11414)
);

OAI21xp5_ASAP7_75t_SL g11415 ( 
.A1(n_11277),
.A2(n_11053),
.B(n_10855),
.Y(n_11415)
);

OAI22xp5_ASAP7_75t_L g11416 ( 
.A1(n_11133),
.A2(n_10995),
.B1(n_11023),
.B2(n_11013),
.Y(n_11416)
);

NAND2xp5_ASAP7_75t_L g11417 ( 
.A(n_11253),
.B(n_11060),
.Y(n_11417)
);

NOR2xp33_ASAP7_75t_R g11418 ( 
.A(n_11288),
.B(n_10970),
.Y(n_11418)
);

AND2x2_ASAP7_75t_L g11419 ( 
.A(n_11296),
.B(n_11055),
.Y(n_11419)
);

AND2x2_ASAP7_75t_L g11420 ( 
.A(n_11199),
.B(n_11022),
.Y(n_11420)
);

AND2x2_ASAP7_75t_L g11421 ( 
.A(n_11191),
.B(n_10963),
.Y(n_11421)
);

NAND2xp5_ASAP7_75t_L g11422 ( 
.A(n_11322),
.B(n_10913),
.Y(n_11422)
);

NAND3xp33_ASAP7_75t_L g11423 ( 
.A(n_11290),
.B(n_10964),
.C(n_10842),
.Y(n_11423)
);

NAND2x1p5_ASAP7_75t_L g11424 ( 
.A(n_11144),
.B(n_11037),
.Y(n_11424)
);

NAND3xp33_ASAP7_75t_L g11425 ( 
.A(n_11364),
.B(n_11084),
.C(n_10900),
.Y(n_11425)
);

AND2x2_ASAP7_75t_L g11426 ( 
.A(n_11170),
.B(n_11038),
.Y(n_11426)
);

NAND2xp5_ASAP7_75t_L g11427 ( 
.A(n_11216),
.B(n_11001),
.Y(n_11427)
);

NAND2xp5_ASAP7_75t_L g11428 ( 
.A(n_11183),
.B(n_11088),
.Y(n_11428)
);

NAND3xp33_ASAP7_75t_L g11429 ( 
.A(n_11297),
.B(n_10971),
.C(n_11048),
.Y(n_11429)
);

AND2x2_ASAP7_75t_L g11430 ( 
.A(n_11142),
.B(n_11062),
.Y(n_11430)
);

OAI22xp5_ASAP7_75t_L g11431 ( 
.A1(n_11197),
.A2(n_11054),
.B1(n_11074),
.B2(n_10882),
.Y(n_11431)
);

OAI22xp5_ASAP7_75t_L g11432 ( 
.A1(n_11375),
.A2(n_10882),
.B1(n_10929),
.B2(n_10967),
.Y(n_11432)
);

NAND2xp5_ASAP7_75t_L g11433 ( 
.A(n_11358),
.B(n_11071),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_11377),
.B(n_1575),
.Y(n_11434)
);

NAND3xp33_ASAP7_75t_L g11435 ( 
.A(n_11139),
.B(n_10929),
.C(n_10849),
.Y(n_11435)
);

NAND4xp25_ASAP7_75t_L g11436 ( 
.A(n_11160),
.B(n_10849),
.C(n_10967),
.D(n_10838),
.Y(n_11436)
);

NOR3xp33_ASAP7_75t_L g11437 ( 
.A(n_11374),
.B(n_10838),
.C(n_11041),
.Y(n_11437)
);

OAI22xp5_ASAP7_75t_L g11438 ( 
.A1(n_11207),
.A2(n_11041),
.B1(n_1578),
.B2(n_1576),
.Y(n_11438)
);

NAND2xp5_ASAP7_75t_L g11439 ( 
.A(n_11321),
.B(n_1577),
.Y(n_11439)
);

NAND3xp33_ASAP7_75t_L g11440 ( 
.A(n_11158),
.B(n_1577),
.C(n_1578),
.Y(n_11440)
);

OAI21xp5_ASAP7_75t_SL g11441 ( 
.A1(n_11177),
.A2(n_1579),
.B(n_1581),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_L g11442 ( 
.A(n_11217),
.B(n_1579),
.Y(n_11442)
);

NOR3xp33_ASAP7_75t_L g11443 ( 
.A(n_11315),
.B(n_1581),
.C(n_1582),
.Y(n_11443)
);

NAND2xp5_ASAP7_75t_L g11444 ( 
.A(n_11223),
.B(n_1583),
.Y(n_11444)
);

NOR3xp33_ASAP7_75t_L g11445 ( 
.A(n_11212),
.B(n_1583),
.C(n_1584),
.Y(n_11445)
);

AND2x2_ASAP7_75t_L g11446 ( 
.A(n_11145),
.B(n_1584),
.Y(n_11446)
);

AND2x2_ASAP7_75t_L g11447 ( 
.A(n_11302),
.B(n_1585),
.Y(n_11447)
);

NAND3xp33_ASAP7_75t_L g11448 ( 
.A(n_11275),
.B(n_1585),
.C(n_1586),
.Y(n_11448)
);

AOI22xp33_ASAP7_75t_SL g11449 ( 
.A1(n_11274),
.A2(n_1588),
.B1(n_1586),
.B2(n_1587),
.Y(n_11449)
);

AND2x2_ASAP7_75t_L g11450 ( 
.A(n_11309),
.B(n_1587),
.Y(n_11450)
);

AND2x2_ASAP7_75t_L g11451 ( 
.A(n_11131),
.B(n_1589),
.Y(n_11451)
);

NAND2xp5_ASAP7_75t_L g11452 ( 
.A(n_11202),
.B(n_1589),
.Y(n_11452)
);

OA21x2_ASAP7_75t_L g11453 ( 
.A1(n_11137),
.A2(n_1590),
.B(n_1591),
.Y(n_11453)
);

NAND3xp33_ASAP7_75t_L g11454 ( 
.A(n_11225),
.B(n_1590),
.C(n_1592),
.Y(n_11454)
);

AOI22xp33_ASAP7_75t_L g11455 ( 
.A1(n_11215),
.A2(n_1594),
.B1(n_1592),
.B2(n_1593),
.Y(n_11455)
);

OAI221xp5_ASAP7_75t_L g11456 ( 
.A1(n_11224),
.A2(n_1595),
.B1(n_1593),
.B2(n_1594),
.C(n_1596),
.Y(n_11456)
);

NAND2xp5_ASAP7_75t_SL g11457 ( 
.A(n_11350),
.B(n_1595),
.Y(n_11457)
);

INVx1_ASAP7_75t_L g11458 ( 
.A(n_11222),
.Y(n_11458)
);

NAND2xp5_ASAP7_75t_L g11459 ( 
.A(n_11249),
.B(n_11267),
.Y(n_11459)
);

OAI221xp5_ASAP7_75t_SL g11460 ( 
.A1(n_11345),
.A2(n_1598),
.B1(n_1596),
.B2(n_1597),
.C(n_1599),
.Y(n_11460)
);

NAND2xp5_ASAP7_75t_SL g11461 ( 
.A(n_11304),
.B(n_1597),
.Y(n_11461)
);

NAND2xp5_ASAP7_75t_L g11462 ( 
.A(n_11267),
.B(n_1598),
.Y(n_11462)
);

NAND2xp5_ASAP7_75t_L g11463 ( 
.A(n_11355),
.B(n_1600),
.Y(n_11463)
);

NAND3xp33_ASAP7_75t_L g11464 ( 
.A(n_11159),
.B(n_1601),
.C(n_1602),
.Y(n_11464)
);

NOR3xp33_ASAP7_75t_SL g11465 ( 
.A(n_11263),
.B(n_1602),
.C(n_1603),
.Y(n_11465)
);

NAND3xp33_ASAP7_75t_L g11466 ( 
.A(n_11165),
.B(n_1603),
.C(n_1605),
.Y(n_11466)
);

OA21x2_ASAP7_75t_L g11467 ( 
.A1(n_11205),
.A2(n_1606),
.B(n_1607),
.Y(n_11467)
);

NAND2xp5_ASAP7_75t_SL g11468 ( 
.A(n_11328),
.B(n_1606),
.Y(n_11468)
);

NAND4xp25_ASAP7_75t_L g11469 ( 
.A(n_11360),
.B(n_1609),
.C(n_1607),
.D(n_1608),
.Y(n_11469)
);

NAND4xp25_ASAP7_75t_L g11470 ( 
.A(n_11363),
.B(n_1611),
.C(n_1608),
.D(n_1610),
.Y(n_11470)
);

NAND2xp5_ASAP7_75t_L g11471 ( 
.A(n_11332),
.B(n_1610),
.Y(n_11471)
);

OAI22xp5_ASAP7_75t_L g11472 ( 
.A1(n_11256),
.A2(n_1614),
.B1(n_1611),
.B2(n_1612),
.Y(n_11472)
);

NOR3xp33_ASAP7_75t_SL g11473 ( 
.A(n_11320),
.B(n_1612),
.C(n_1614),
.Y(n_11473)
);

AOI221xp5_ASAP7_75t_L g11474 ( 
.A1(n_11265),
.A2(n_1617),
.B1(n_1615),
.B2(n_1616),
.C(n_1618),
.Y(n_11474)
);

AND2x2_ASAP7_75t_L g11475 ( 
.A(n_11226),
.B(n_1615),
.Y(n_11475)
);

AND2x2_ASAP7_75t_L g11476 ( 
.A(n_11172),
.B(n_1616),
.Y(n_11476)
);

OAI21xp33_ASAP7_75t_L g11477 ( 
.A1(n_11234),
.A2(n_1617),
.B(n_1618),
.Y(n_11477)
);

OAI211xp5_ASAP7_75t_L g11478 ( 
.A1(n_11373),
.A2(n_11178),
.B(n_11378),
.C(n_11235),
.Y(n_11478)
);

AOI21xp5_ASAP7_75t_SL g11479 ( 
.A1(n_11312),
.A2(n_1619),
.B(n_1620),
.Y(n_11479)
);

AND2x2_ASAP7_75t_L g11480 ( 
.A(n_11182),
.B(n_1620),
.Y(n_11480)
);

AND2x2_ASAP7_75t_L g11481 ( 
.A(n_11184),
.B(n_1621),
.Y(n_11481)
);

NAND2xp5_ASAP7_75t_L g11482 ( 
.A(n_11351),
.B(n_1621),
.Y(n_11482)
);

NAND4xp25_ASAP7_75t_L g11483 ( 
.A(n_11365),
.B(n_1624),
.C(n_1622),
.D(n_1623),
.Y(n_11483)
);

NAND2xp5_ASAP7_75t_L g11484 ( 
.A(n_11353),
.B(n_1622),
.Y(n_11484)
);

AND2x2_ASAP7_75t_L g11485 ( 
.A(n_11188),
.B(n_1624),
.Y(n_11485)
);

AOI21xp5_ASAP7_75t_SL g11486 ( 
.A1(n_11366),
.A2(n_1625),
.B(n_1626),
.Y(n_11486)
);

OAI21xp33_ASAP7_75t_L g11487 ( 
.A1(n_11238),
.A2(n_1625),
.B(n_1626),
.Y(n_11487)
);

AND2x2_ASAP7_75t_L g11488 ( 
.A(n_11206),
.B(n_1627),
.Y(n_11488)
);

AND2x2_ASAP7_75t_L g11489 ( 
.A(n_11211),
.B(n_1627),
.Y(n_11489)
);

NAND3xp33_ASAP7_75t_L g11490 ( 
.A(n_11336),
.B(n_1628),
.C(n_1629),
.Y(n_11490)
);

AND2x2_ASAP7_75t_L g11491 ( 
.A(n_11272),
.B(n_1628),
.Y(n_11491)
);

OAI221xp5_ASAP7_75t_SL g11492 ( 
.A1(n_11173),
.A2(n_1632),
.B1(n_1630),
.B2(n_1631),
.C(n_1633),
.Y(n_11492)
);

AND2x2_ASAP7_75t_SL g11493 ( 
.A(n_11213),
.B(n_1631),
.Y(n_11493)
);

AND2x2_ASAP7_75t_L g11494 ( 
.A(n_11282),
.B(n_1633),
.Y(n_11494)
);

OAI22xp5_ASAP7_75t_L g11495 ( 
.A1(n_11337),
.A2(n_1636),
.B1(n_1634),
.B2(n_1635),
.Y(n_11495)
);

AND2x2_ASAP7_75t_L g11496 ( 
.A(n_11283),
.B(n_1634),
.Y(n_11496)
);

NAND3xp33_ASAP7_75t_L g11497 ( 
.A(n_11269),
.B(n_1635),
.C(n_1636),
.Y(n_11497)
);

NAND2xp5_ASAP7_75t_SL g11498 ( 
.A(n_11260),
.B(n_1637),
.Y(n_11498)
);

NAND2xp5_ASAP7_75t_SL g11499 ( 
.A(n_11284),
.B(n_1637),
.Y(n_11499)
);

NAND3xp33_ASAP7_75t_L g11500 ( 
.A(n_11228),
.B(n_1638),
.C(n_1639),
.Y(n_11500)
);

AOI22xp33_ASAP7_75t_L g11501 ( 
.A1(n_11246),
.A2(n_11248),
.B1(n_11251),
.B2(n_11250),
.Y(n_11501)
);

NAND2xp5_ASAP7_75t_L g11502 ( 
.A(n_11361),
.B(n_1638),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_11285),
.B(n_1639),
.Y(n_11503)
);

NOR2xp33_ASAP7_75t_L g11504 ( 
.A(n_11193),
.B(n_1640),
.Y(n_11504)
);

AOI22xp33_ASAP7_75t_SL g11505 ( 
.A1(n_11194),
.A2(n_1643),
.B1(n_1641),
.B2(n_1642),
.Y(n_11505)
);

AND2x2_ASAP7_75t_L g11506 ( 
.A(n_11362),
.B(n_1643),
.Y(n_11506)
);

NOR3xp33_ASAP7_75t_L g11507 ( 
.A(n_11140),
.B(n_1644),
.C(n_1645),
.Y(n_11507)
);

AND2x2_ASAP7_75t_L g11508 ( 
.A(n_11294),
.B(n_1645),
.Y(n_11508)
);

NOR3xp33_ASAP7_75t_L g11509 ( 
.A(n_11273),
.B(n_1646),
.C(n_1647),
.Y(n_11509)
);

NAND2xp5_ASAP7_75t_L g11510 ( 
.A(n_11298),
.B(n_1646),
.Y(n_11510)
);

AND2x2_ASAP7_75t_L g11511 ( 
.A(n_11299),
.B(n_1647),
.Y(n_11511)
);

NAND2x1p5_ASAP7_75t_L g11512 ( 
.A(n_11201),
.B(n_1648),
.Y(n_11512)
);

NAND2xp5_ASAP7_75t_L g11513 ( 
.A(n_11303),
.B(n_1649),
.Y(n_11513)
);

AOI22xp5_ASAP7_75t_L g11514 ( 
.A1(n_11305),
.A2(n_1651),
.B1(n_1649),
.B2(n_1650),
.Y(n_11514)
);

NAND2xp5_ASAP7_75t_L g11515 ( 
.A(n_11306),
.B(n_1652),
.Y(n_11515)
);

NAND2xp5_ASAP7_75t_SL g11516 ( 
.A(n_11301),
.B(n_1652),
.Y(n_11516)
);

NAND3xp33_ASAP7_75t_L g11517 ( 
.A(n_11276),
.B(n_1653),
.C(n_1654),
.Y(n_11517)
);

AND2x2_ASAP7_75t_L g11518 ( 
.A(n_11308),
.B(n_11310),
.Y(n_11518)
);

OAI22xp5_ASAP7_75t_L g11519 ( 
.A1(n_11316),
.A2(n_1656),
.B1(n_1654),
.B2(n_1655),
.Y(n_11519)
);

NAND2xp5_ASAP7_75t_L g11520 ( 
.A(n_11339),
.B(n_1656),
.Y(n_11520)
);

NAND2xp5_ASAP7_75t_L g11521 ( 
.A(n_11346),
.B(n_1657),
.Y(n_11521)
);

OAI21xp5_ASAP7_75t_L g11522 ( 
.A1(n_11243),
.A2(n_1657),
.B(n_1658),
.Y(n_11522)
);

OAI22xp5_ASAP7_75t_L g11523 ( 
.A1(n_11311),
.A2(n_1660),
.B1(n_1658),
.B2(n_1659),
.Y(n_11523)
);

NAND2xp5_ASAP7_75t_SL g11524 ( 
.A(n_11317),
.B(n_1659),
.Y(n_11524)
);

AND2x2_ASAP7_75t_L g11525 ( 
.A(n_11318),
.B(n_1660),
.Y(n_11525)
);

NAND2xp5_ASAP7_75t_L g11526 ( 
.A(n_11324),
.B(n_11344),
.Y(n_11526)
);

NAND2xp5_ASAP7_75t_L g11527 ( 
.A(n_11349),
.B(n_1661),
.Y(n_11527)
);

NAND3xp33_ASAP7_75t_L g11528 ( 
.A(n_11292),
.B(n_1661),
.C(n_1662),
.Y(n_11528)
);

AOI21xp5_ASAP7_75t_SL g11529 ( 
.A1(n_11173),
.A2(n_11335),
.B(n_11148),
.Y(n_11529)
);

NAND2xp5_ASAP7_75t_SL g11530 ( 
.A(n_11146),
.B(n_1662),
.Y(n_11530)
);

NAND3xp33_ASAP7_75t_L g11531 ( 
.A(n_11141),
.B(n_1663),
.C(n_1664),
.Y(n_11531)
);

AND2x2_ASAP7_75t_L g11532 ( 
.A(n_11175),
.B(n_1665),
.Y(n_11532)
);

INVxp33_ASAP7_75t_L g11533 ( 
.A(n_11190),
.Y(n_11533)
);

NAND2xp5_ASAP7_75t_L g11534 ( 
.A(n_11176),
.B(n_1665),
.Y(n_11534)
);

NAND2xp5_ASAP7_75t_SL g11535 ( 
.A(n_11289),
.B(n_1666),
.Y(n_11535)
);

OA21x2_ASAP7_75t_L g11536 ( 
.A1(n_11150),
.A2(n_1666),
.B(n_1667),
.Y(n_11536)
);

NOR3xp33_ASAP7_75t_L g11537 ( 
.A(n_11367),
.B(n_1668),
.C(n_1669),
.Y(n_11537)
);

OAI22xp5_ASAP7_75t_L g11538 ( 
.A1(n_11147),
.A2(n_1671),
.B1(n_1669),
.B2(n_1670),
.Y(n_11538)
);

AND2x2_ASAP7_75t_L g11539 ( 
.A(n_11130),
.B(n_1671),
.Y(n_11539)
);

NAND2xp5_ASAP7_75t_L g11540 ( 
.A(n_11152),
.B(n_1672),
.Y(n_11540)
);

OAI221xp5_ASAP7_75t_SL g11541 ( 
.A1(n_11221),
.A2(n_1674),
.B1(n_1672),
.B2(n_1673),
.C(n_1675),
.Y(n_11541)
);

OAI221xp5_ASAP7_75t_SL g11542 ( 
.A1(n_11245),
.A2(n_1675),
.B1(n_1673),
.B2(n_1674),
.C(n_1676),
.Y(n_11542)
);

INVx2_ASAP7_75t_L g11543 ( 
.A(n_11136),
.Y(n_11543)
);

AOI221xp5_ASAP7_75t_L g11544 ( 
.A1(n_11151),
.A2(n_1679),
.B1(n_1677),
.B2(n_1678),
.C(n_1681),
.Y(n_11544)
);

NAND3xp33_ASAP7_75t_L g11545 ( 
.A(n_11154),
.B(n_1679),
.C(n_1681),
.Y(n_11545)
);

NAND2xp5_ASAP7_75t_L g11546 ( 
.A(n_11208),
.B(n_1682),
.Y(n_11546)
);

NOR2xp33_ASAP7_75t_R g11547 ( 
.A(n_11348),
.B(n_11270),
.Y(n_11547)
);

AOI221xp5_ASAP7_75t_L g11548 ( 
.A1(n_11155),
.A2(n_1685),
.B1(n_1682),
.B2(n_1683),
.C(n_1686),
.Y(n_11548)
);

NAND2xp5_ASAP7_75t_L g11549 ( 
.A(n_11259),
.B(n_1685),
.Y(n_11549)
);

NAND2xp5_ASAP7_75t_L g11550 ( 
.A(n_11187),
.B(n_1686),
.Y(n_11550)
);

NAND2xp5_ASAP7_75t_L g11551 ( 
.A(n_11174),
.B(n_1687),
.Y(n_11551)
);

NAND2xp5_ASAP7_75t_L g11552 ( 
.A(n_11186),
.B(n_1688),
.Y(n_11552)
);

OAI22xp5_ASAP7_75t_L g11553 ( 
.A1(n_11153),
.A2(n_1691),
.B1(n_1689),
.B2(n_1690),
.Y(n_11553)
);

NAND2xp5_ASAP7_75t_L g11554 ( 
.A(n_11179),
.B(n_1689),
.Y(n_11554)
);

OA21x2_ASAP7_75t_L g11555 ( 
.A1(n_11157),
.A2(n_1690),
.B(n_1692),
.Y(n_11555)
);

OAI22xp5_ASAP7_75t_L g11556 ( 
.A1(n_11168),
.A2(n_11162),
.B1(n_11163),
.B2(n_11161),
.Y(n_11556)
);

NAND2xp5_ASAP7_75t_L g11557 ( 
.A(n_11156),
.B(n_1692),
.Y(n_11557)
);

AND2x2_ASAP7_75t_L g11558 ( 
.A(n_11210),
.B(n_1693),
.Y(n_11558)
);

AOI22xp33_ASAP7_75t_L g11559 ( 
.A1(n_11166),
.A2(n_1695),
.B1(n_1693),
.B2(n_1694),
.Y(n_11559)
);

NAND2xp5_ASAP7_75t_L g11560 ( 
.A(n_11169),
.B(n_1694),
.Y(n_11560)
);

AND2x2_ASAP7_75t_L g11561 ( 
.A(n_11329),
.B(n_1695),
.Y(n_11561)
);

OAI22xp5_ASAP7_75t_L g11562 ( 
.A1(n_11167),
.A2(n_1698),
.B1(n_1696),
.B2(n_1697),
.Y(n_11562)
);

AND2x2_ASAP7_75t_L g11563 ( 
.A(n_11368),
.B(n_1696),
.Y(n_11563)
);

NAND2xp5_ASAP7_75t_L g11564 ( 
.A(n_11149),
.B(n_1697),
.Y(n_11564)
);

AOI22xp33_ASAP7_75t_L g11565 ( 
.A1(n_11171),
.A2(n_1700),
.B1(n_1698),
.B2(n_1699),
.Y(n_11565)
);

NAND2xp5_ASAP7_75t_L g11566 ( 
.A(n_11354),
.B(n_1699),
.Y(n_11566)
);

NAND2xp5_ASAP7_75t_L g11567 ( 
.A(n_11359),
.B(n_1700),
.Y(n_11567)
);

AOI22xp33_ASAP7_75t_SL g11568 ( 
.A1(n_11192),
.A2(n_1703),
.B1(n_1701),
.B2(n_1702),
.Y(n_11568)
);

NAND2xp5_ASAP7_75t_L g11569 ( 
.A(n_11261),
.B(n_1702),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_L g11570 ( 
.A(n_11262),
.B(n_1703),
.Y(n_11570)
);

AND2x2_ASAP7_75t_L g11571 ( 
.A(n_11266),
.B(n_1704),
.Y(n_11571)
);

AND2x2_ASAP7_75t_L g11572 ( 
.A(n_11279),
.B(n_11287),
.Y(n_11572)
);

NAND2xp5_ASAP7_75t_L g11573 ( 
.A(n_11300),
.B(n_1704),
.Y(n_11573)
);

NAND4xp25_ASAP7_75t_L g11574 ( 
.A(n_11195),
.B(n_1707),
.C(n_1705),
.D(n_1706),
.Y(n_11574)
);

NAND2xp5_ASAP7_75t_SL g11575 ( 
.A(n_11185),
.B(n_1706),
.Y(n_11575)
);

OAI21xp5_ASAP7_75t_SL g11576 ( 
.A1(n_11198),
.A2(n_1707),
.B(n_1708),
.Y(n_11576)
);

AOI221xp5_ASAP7_75t_L g11577 ( 
.A1(n_11200),
.A2(n_1711),
.B1(n_1709),
.B2(n_1710),
.C(n_1712),
.Y(n_11577)
);

NAND3xp33_ASAP7_75t_L g11578 ( 
.A(n_11204),
.B(n_1709),
.C(n_1710),
.Y(n_11578)
);

AND2x2_ASAP7_75t_L g11579 ( 
.A(n_11307),
.B(n_1711),
.Y(n_11579)
);

AND2x2_ASAP7_75t_L g11580 ( 
.A(n_11313),
.B(n_1712),
.Y(n_11580)
);

INVx2_ASAP7_75t_L g11581 ( 
.A(n_11392),
.Y(n_11581)
);

AND2x2_ASAP7_75t_L g11582 ( 
.A(n_11386),
.B(n_11314),
.Y(n_11582)
);

AND2x4_ASAP7_75t_L g11583 ( 
.A(n_11395),
.B(n_11134),
.Y(n_11583)
);

INVx2_ASAP7_75t_L g11584 ( 
.A(n_11419),
.Y(n_11584)
);

AND2x2_ASAP7_75t_L g11585 ( 
.A(n_11420),
.B(n_11319),
.Y(n_11585)
);

INVxp67_ASAP7_75t_L g11586 ( 
.A(n_11391),
.Y(n_11586)
);

AO21x2_ASAP7_75t_L g11587 ( 
.A1(n_11394),
.A2(n_11214),
.B(n_11180),
.Y(n_11587)
);

INVx1_ASAP7_75t_SL g11588 ( 
.A(n_11493),
.Y(n_11588)
);

BUFx2_ASAP7_75t_L g11589 ( 
.A(n_11418),
.Y(n_11589)
);

INVx2_ASAP7_75t_L g11590 ( 
.A(n_11512),
.Y(n_11590)
);

INVx1_ASAP7_75t_L g11591 ( 
.A(n_11508),
.Y(n_11591)
);

NAND2xp5_ASAP7_75t_L g11592 ( 
.A(n_11437),
.B(n_11323),
.Y(n_11592)
);

AND2x2_ASAP7_75t_L g11593 ( 
.A(n_11390),
.B(n_11327),
.Y(n_11593)
);

INVx1_ASAP7_75t_L g11594 ( 
.A(n_11511),
.Y(n_11594)
);

OR2x2_ASAP7_75t_L g11595 ( 
.A(n_11383),
.B(n_11343),
.Y(n_11595)
);

INVxp67_ASAP7_75t_L g11596 ( 
.A(n_11398),
.Y(n_11596)
);

INVx1_ASAP7_75t_L g11597 ( 
.A(n_11525),
.Y(n_11597)
);

OAI31xp33_ASAP7_75t_L g11598 ( 
.A1(n_11381),
.A2(n_11264),
.A3(n_11286),
.B(n_11280),
.Y(n_11598)
);

AND2x2_ASAP7_75t_L g11599 ( 
.A(n_11421),
.B(n_11330),
.Y(n_11599)
);

OR2x2_ASAP7_75t_L g11600 ( 
.A(n_11403),
.B(n_11385),
.Y(n_11600)
);

NAND2xp5_ASAP7_75t_L g11601 ( 
.A(n_11432),
.B(n_11242),
.Y(n_11601)
);

NAND2xp5_ASAP7_75t_SL g11602 ( 
.A(n_11409),
.B(n_11143),
.Y(n_11602)
);

NAND3xp33_ASAP7_75t_L g11603 ( 
.A(n_11384),
.B(n_11232),
.C(n_11209),
.Y(n_11603)
);

AND2x2_ASAP7_75t_L g11604 ( 
.A(n_11572),
.B(n_11338),
.Y(n_11604)
);

OAI211xp5_ASAP7_75t_L g11605 ( 
.A1(n_11382),
.A2(n_11244),
.B(n_11255),
.C(n_11237),
.Y(n_11605)
);

AOI22xp5_ASAP7_75t_L g11606 ( 
.A1(n_11380),
.A2(n_11268),
.B1(n_11271),
.B2(n_11258),
.Y(n_11606)
);

INVx5_ASAP7_75t_L g11607 ( 
.A(n_11488),
.Y(n_11607)
);

AND2x2_ASAP7_75t_L g11608 ( 
.A(n_11426),
.B(n_11340),
.Y(n_11608)
);

INVx4_ASAP7_75t_L g11609 ( 
.A(n_11447),
.Y(n_11609)
);

OR2x2_ASAP7_75t_L g11610 ( 
.A(n_11389),
.B(n_11278),
.Y(n_11610)
);

AND2x4_ASAP7_75t_L g11611 ( 
.A(n_11543),
.B(n_11218),
.Y(n_11611)
);

INVx3_ASAP7_75t_L g11612 ( 
.A(n_11424),
.Y(n_11612)
);

INVxp67_ASAP7_75t_L g11613 ( 
.A(n_11489),
.Y(n_11613)
);

INVx2_ASAP7_75t_L g11614 ( 
.A(n_11491),
.Y(n_11614)
);

INVx2_ASAP7_75t_L g11615 ( 
.A(n_11450),
.Y(n_11615)
);

BUFx2_ASAP7_75t_L g11616 ( 
.A(n_11547),
.Y(n_11616)
);

NAND2xp5_ASAP7_75t_L g11617 ( 
.A(n_11404),
.B(n_11396),
.Y(n_11617)
);

INVxp67_ASAP7_75t_SL g11618 ( 
.A(n_11414),
.Y(n_11618)
);

INVx2_ASAP7_75t_L g11619 ( 
.A(n_11446),
.Y(n_11619)
);

HB1xp67_ASAP7_75t_L g11620 ( 
.A(n_11467),
.Y(n_11620)
);

INVx1_ASAP7_75t_L g11621 ( 
.A(n_11494),
.Y(n_11621)
);

NAND2xp5_ASAP7_75t_L g11622 ( 
.A(n_11465),
.B(n_11247),
.Y(n_11622)
);

INVx1_ASAP7_75t_L g11623 ( 
.A(n_11496),
.Y(n_11623)
);

INVx1_ASAP7_75t_L g11624 ( 
.A(n_11503),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_11506),
.Y(n_11625)
);

INVx1_ASAP7_75t_SL g11626 ( 
.A(n_11433),
.Y(n_11626)
);

AOI322xp5_ASAP7_75t_L g11627 ( 
.A1(n_11393),
.A2(n_11252),
.A3(n_11370),
.B1(n_11371),
.B2(n_11369),
.C1(n_11220),
.C2(n_11254),
.Y(n_11627)
);

AND2x4_ASAP7_75t_L g11628 ( 
.A(n_11518),
.B(n_11430),
.Y(n_11628)
);

INVx2_ASAP7_75t_L g11629 ( 
.A(n_11451),
.Y(n_11629)
);

NOR2xp33_ASAP7_75t_L g11630 ( 
.A(n_11533),
.B(n_11333),
.Y(n_11630)
);

AND2x2_ASAP7_75t_L g11631 ( 
.A(n_11501),
.B(n_11291),
.Y(n_11631)
);

INVx2_ASAP7_75t_L g11632 ( 
.A(n_11475),
.Y(n_11632)
);

OAI21xp5_ASAP7_75t_L g11633 ( 
.A1(n_11401),
.A2(n_1713),
.B(n_1714),
.Y(n_11633)
);

INVx1_ASAP7_75t_L g11634 ( 
.A(n_11463),
.Y(n_11634)
);

INVx1_ASAP7_75t_L g11635 ( 
.A(n_11526),
.Y(n_11635)
);

OR2x2_ASAP7_75t_L g11636 ( 
.A(n_11428),
.B(n_1713),
.Y(n_11636)
);

AND2x4_ASAP7_75t_L g11637 ( 
.A(n_11422),
.B(n_1714),
.Y(n_11637)
);

AND2x4_ASAP7_75t_L g11638 ( 
.A(n_11458),
.B(n_1715),
.Y(n_11638)
);

AO21x2_ASAP7_75t_L g11639 ( 
.A1(n_11407),
.A2(n_1715),
.B(n_1716),
.Y(n_11639)
);

AND2x2_ASAP7_75t_L g11640 ( 
.A(n_11402),
.B(n_1716),
.Y(n_11640)
);

OR2x2_ASAP7_75t_L g11641 ( 
.A(n_11412),
.B(n_1717),
.Y(n_11641)
);

BUFx2_ASAP7_75t_L g11642 ( 
.A(n_11467),
.Y(n_11642)
);

INVx1_ASAP7_75t_L g11643 ( 
.A(n_11482),
.Y(n_11643)
);

OAI31xp33_ASAP7_75t_L g11644 ( 
.A1(n_11425),
.A2(n_1719),
.A3(n_1717),
.B(n_1718),
.Y(n_11644)
);

NOR2xp33_ASAP7_75t_L g11645 ( 
.A(n_11410),
.B(n_1718),
.Y(n_11645)
);

INVx2_ASAP7_75t_L g11646 ( 
.A(n_11476),
.Y(n_11646)
);

NAND4xp25_ASAP7_75t_SL g11647 ( 
.A(n_11405),
.B(n_1721),
.C(n_1719),
.D(n_1720),
.Y(n_11647)
);

INVx1_ASAP7_75t_L g11648 ( 
.A(n_11484),
.Y(n_11648)
);

INVx1_ASAP7_75t_L g11649 ( 
.A(n_11434),
.Y(n_11649)
);

OAI22xp5_ASAP7_75t_L g11650 ( 
.A1(n_11423),
.A2(n_1722),
.B1(n_1720),
.B2(n_1721),
.Y(n_11650)
);

OAI221xp5_ASAP7_75t_L g11651 ( 
.A1(n_11399),
.A2(n_1725),
.B1(n_1723),
.B2(n_1724),
.C(n_1726),
.Y(n_11651)
);

INVx1_ASAP7_75t_L g11652 ( 
.A(n_11566),
.Y(n_11652)
);

NAND2xp5_ASAP7_75t_L g11653 ( 
.A(n_11443),
.B(n_1724),
.Y(n_11653)
);

CKINVDCx20_ASAP7_75t_R g11654 ( 
.A(n_11473),
.Y(n_11654)
);

NAND2xp5_ASAP7_75t_SL g11655 ( 
.A(n_11449),
.B(n_1725),
.Y(n_11655)
);

OAI221xp5_ASAP7_75t_SL g11656 ( 
.A1(n_11411),
.A2(n_1729),
.B1(n_1726),
.B2(n_1727),
.C(n_1730),
.Y(n_11656)
);

BUFx3_ASAP7_75t_L g11657 ( 
.A(n_11480),
.Y(n_11657)
);

INVx1_ASAP7_75t_L g11658 ( 
.A(n_11567),
.Y(n_11658)
);

AND2x2_ASAP7_75t_L g11659 ( 
.A(n_11529),
.B(n_1727),
.Y(n_11659)
);

INVx1_ASAP7_75t_L g11660 ( 
.A(n_11471),
.Y(n_11660)
);

AOI22xp33_ASAP7_75t_SL g11661 ( 
.A1(n_11413),
.A2(n_11431),
.B1(n_11435),
.B2(n_11416),
.Y(n_11661)
);

INVx1_ASAP7_75t_L g11662 ( 
.A(n_11527),
.Y(n_11662)
);

OR2x2_ASAP7_75t_L g11663 ( 
.A(n_11387),
.B(n_1729),
.Y(n_11663)
);

AOI22xp33_ASAP7_75t_L g11664 ( 
.A1(n_11406),
.A2(n_1733),
.B1(n_1731),
.B2(n_1732),
.Y(n_11664)
);

INVx2_ASAP7_75t_L g11665 ( 
.A(n_11481),
.Y(n_11665)
);

OAI33xp33_ASAP7_75t_L g11666 ( 
.A1(n_11388),
.A2(n_1734),
.A3(n_1736),
.B1(n_1731),
.B2(n_1732),
.B3(n_1735),
.Y(n_11666)
);

INVx1_ASAP7_75t_L g11667 ( 
.A(n_11569),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_11570),
.Y(n_11668)
);

INVx1_ASAP7_75t_L g11669 ( 
.A(n_11573),
.Y(n_11669)
);

NOR2xp33_ASAP7_75t_L g11670 ( 
.A(n_11441),
.B(n_1734),
.Y(n_11670)
);

OR2x6_ASAP7_75t_L g11671 ( 
.A(n_11479),
.B(n_1735),
.Y(n_11671)
);

AND2x2_ASAP7_75t_L g11672 ( 
.A(n_11532),
.B(n_1736),
.Y(n_11672)
);

INVx1_ASAP7_75t_L g11673 ( 
.A(n_11502),
.Y(n_11673)
);

OR2x6_ASAP7_75t_L g11674 ( 
.A(n_11486),
.B(n_1738),
.Y(n_11674)
);

INVx1_ASAP7_75t_L g11675 ( 
.A(n_11452),
.Y(n_11675)
);

INVx2_ASAP7_75t_L g11676 ( 
.A(n_11485),
.Y(n_11676)
);

INVx1_ASAP7_75t_L g11677 ( 
.A(n_11550),
.Y(n_11677)
);

OR2x2_ASAP7_75t_L g11678 ( 
.A(n_11400),
.B(n_11417),
.Y(n_11678)
);

INVx2_ASAP7_75t_L g11679 ( 
.A(n_11539),
.Y(n_11679)
);

INVx2_ASAP7_75t_L g11680 ( 
.A(n_11558),
.Y(n_11680)
);

AND2x2_ASAP7_75t_L g11681 ( 
.A(n_11571),
.B(n_2918),
.Y(n_11681)
);

AND2x2_ASAP7_75t_L g11682 ( 
.A(n_11579),
.B(n_2918),
.Y(n_11682)
);

INVx2_ASAP7_75t_L g11683 ( 
.A(n_11561),
.Y(n_11683)
);

HB1xp67_ASAP7_75t_L g11684 ( 
.A(n_11536),
.Y(n_11684)
);

INVx4_ASAP7_75t_L g11685 ( 
.A(n_11563),
.Y(n_11685)
);

AND2x2_ASAP7_75t_L g11686 ( 
.A(n_11580),
.B(n_2919),
.Y(n_11686)
);

NAND2x1_ASAP7_75t_L g11687 ( 
.A(n_11536),
.B(n_1738),
.Y(n_11687)
);

OR2x2_ASAP7_75t_L g11688 ( 
.A(n_11427),
.B(n_1739),
.Y(n_11688)
);

OR2x2_ASAP7_75t_L g11689 ( 
.A(n_11436),
.B(n_1740),
.Y(n_11689)
);

AND2x2_ASAP7_75t_L g11690 ( 
.A(n_11397),
.B(n_1740),
.Y(n_11690)
);

INVxp67_ASAP7_75t_L g11691 ( 
.A(n_11461),
.Y(n_11691)
);

AOI221xp5_ASAP7_75t_L g11692 ( 
.A1(n_11556),
.A2(n_1744),
.B1(n_1741),
.B2(n_1743),
.C(n_1745),
.Y(n_11692)
);

NAND2xp5_ASAP7_75t_L g11693 ( 
.A(n_11408),
.B(n_1741),
.Y(n_11693)
);

NAND2xp33_ASAP7_75t_R g11694 ( 
.A(n_11453),
.B(n_2907),
.Y(n_11694)
);

NAND2xp5_ASAP7_75t_L g11695 ( 
.A(n_11537),
.B(n_11507),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_11551),
.Y(n_11696)
);

OR2x2_ASAP7_75t_L g11697 ( 
.A(n_11459),
.B(n_1744),
.Y(n_11697)
);

AND2x4_ASAP7_75t_L g11698 ( 
.A(n_11445),
.B(n_1745),
.Y(n_11698)
);

INVx2_ASAP7_75t_L g11699 ( 
.A(n_11555),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_11552),
.Y(n_11700)
);

OR2x6_ASAP7_75t_L g11701 ( 
.A(n_11444),
.B(n_1746),
.Y(n_11701)
);

AOI22xp33_ASAP7_75t_L g11702 ( 
.A1(n_11429),
.A2(n_1748),
.B1(n_1746),
.B2(n_1747),
.Y(n_11702)
);

INVx1_ASAP7_75t_L g11703 ( 
.A(n_11546),
.Y(n_11703)
);

AOI22xp33_ASAP7_75t_L g11704 ( 
.A1(n_11438),
.A2(n_1749),
.B1(n_1747),
.B2(n_1748),
.Y(n_11704)
);

INVx2_ASAP7_75t_L g11705 ( 
.A(n_11555),
.Y(n_11705)
);

INVx2_ASAP7_75t_L g11706 ( 
.A(n_11564),
.Y(n_11706)
);

OAI21xp5_ASAP7_75t_L g11707 ( 
.A1(n_11415),
.A2(n_1750),
.B(n_1751),
.Y(n_11707)
);

OAI221xp5_ASAP7_75t_L g11708 ( 
.A1(n_11462),
.A2(n_1754),
.B1(n_1751),
.B2(n_1752),
.C(n_1755),
.Y(n_11708)
);

CKINVDCx16_ASAP7_75t_R g11709 ( 
.A(n_11522),
.Y(n_11709)
);

AOI33xp33_ASAP7_75t_L g11710 ( 
.A1(n_11505),
.A2(n_1756),
.A3(n_1758),
.B1(n_1754),
.B2(n_1755),
.B3(n_1757),
.Y(n_11710)
);

AND2x2_ASAP7_75t_L g11711 ( 
.A(n_11504),
.B(n_2920),
.Y(n_11711)
);

INVx2_ASAP7_75t_L g11712 ( 
.A(n_11560),
.Y(n_11712)
);

OR2x2_ASAP7_75t_L g11713 ( 
.A(n_11439),
.B(n_1756),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_11530),
.B(n_11453),
.Y(n_11714)
);

NOR2x1_ASAP7_75t_SL g11715 ( 
.A(n_11448),
.B(n_1757),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_11457),
.B(n_2905),
.Y(n_11716)
);

INVx3_ASAP7_75t_L g11717 ( 
.A(n_11557),
.Y(n_11717)
);

HB1xp67_ASAP7_75t_L g11718 ( 
.A(n_11575),
.Y(n_11718)
);

NAND2xp5_ASAP7_75t_SL g11719 ( 
.A(n_11500),
.B(n_1759),
.Y(n_11719)
);

NAND2xp5_ASAP7_75t_L g11720 ( 
.A(n_11509),
.B(n_1759),
.Y(n_11720)
);

AND2x2_ASAP7_75t_L g11721 ( 
.A(n_11468),
.B(n_2907),
.Y(n_11721)
);

AND2x4_ASAP7_75t_L g11722 ( 
.A(n_11535),
.B(n_1760),
.Y(n_11722)
);

OR2x2_ASAP7_75t_L g11723 ( 
.A(n_11478),
.B(n_11510),
.Y(n_11723)
);

AND2x2_ASAP7_75t_L g11724 ( 
.A(n_11513),
.B(n_2909),
.Y(n_11724)
);

AOI33xp33_ASAP7_75t_L g11725 ( 
.A1(n_11568),
.A2(n_1763),
.A3(n_1765),
.B1(n_1761),
.B2(n_1762),
.B3(n_1764),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_11534),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11540),
.Y(n_11727)
);

INVxp67_ASAP7_75t_L g11728 ( 
.A(n_11498),
.Y(n_11728)
);

INVx2_ASAP7_75t_L g11729 ( 
.A(n_11554),
.Y(n_11729)
);

NAND2xp5_ASAP7_75t_L g11730 ( 
.A(n_11576),
.B(n_1761),
.Y(n_11730)
);

INVx1_ASAP7_75t_L g11731 ( 
.A(n_11549),
.Y(n_11731)
);

NAND2xp5_ASAP7_75t_L g11732 ( 
.A(n_11477),
.B(n_1763),
.Y(n_11732)
);

NOR3xp33_ASAP7_75t_L g11733 ( 
.A(n_11454),
.B(n_1764),
.C(n_1765),
.Y(n_11733)
);

INVx1_ASAP7_75t_L g11734 ( 
.A(n_11515),
.Y(n_11734)
);

INVx2_ASAP7_75t_L g11735 ( 
.A(n_11442),
.Y(n_11735)
);

AND2x4_ASAP7_75t_L g11736 ( 
.A(n_11499),
.B(n_11516),
.Y(n_11736)
);

OR2x2_ASAP7_75t_L g11737 ( 
.A(n_11588),
.B(n_11520),
.Y(n_11737)
);

INVx1_ASAP7_75t_L g11738 ( 
.A(n_11620),
.Y(n_11738)
);

AND2x2_ASAP7_75t_L g11739 ( 
.A(n_11589),
.B(n_11521),
.Y(n_11739)
);

AND2x2_ASAP7_75t_L g11740 ( 
.A(n_11607),
.B(n_11524),
.Y(n_11740)
);

INVxp67_ASAP7_75t_L g11741 ( 
.A(n_11694),
.Y(n_11741)
);

INVx1_ASAP7_75t_SL g11742 ( 
.A(n_11607),
.Y(n_11742)
);

INVx2_ASAP7_75t_L g11743 ( 
.A(n_11612),
.Y(n_11743)
);

HB1xp67_ASAP7_75t_L g11744 ( 
.A(n_11674),
.Y(n_11744)
);

AND2x2_ASAP7_75t_L g11745 ( 
.A(n_11582),
.B(n_11487),
.Y(n_11745)
);

INVx2_ASAP7_75t_L g11746 ( 
.A(n_11583),
.Y(n_11746)
);

HB1xp67_ASAP7_75t_L g11747 ( 
.A(n_11674),
.Y(n_11747)
);

INVx2_ASAP7_75t_L g11748 ( 
.A(n_11581),
.Y(n_11748)
);

NAND2xp5_ASAP7_75t_L g11749 ( 
.A(n_11618),
.B(n_11497),
.Y(n_11749)
);

HB1xp67_ASAP7_75t_L g11750 ( 
.A(n_11671),
.Y(n_11750)
);

NAND2xp33_ASAP7_75t_SL g11751 ( 
.A(n_11687),
.B(n_11495),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_11642),
.Y(n_11752)
);

AND2x2_ASAP7_75t_L g11753 ( 
.A(n_11593),
.B(n_11464),
.Y(n_11753)
);

OR2x2_ASAP7_75t_L g11754 ( 
.A(n_11613),
.B(n_11490),
.Y(n_11754)
);

INVx1_ASAP7_75t_L g11755 ( 
.A(n_11684),
.Y(n_11755)
);

INVx2_ASAP7_75t_L g11756 ( 
.A(n_11584),
.Y(n_11756)
);

AND2x2_ASAP7_75t_L g11757 ( 
.A(n_11616),
.B(n_11466),
.Y(n_11757)
);

INVx1_ASAP7_75t_L g11758 ( 
.A(n_11672),
.Y(n_11758)
);

AND2x2_ASAP7_75t_L g11759 ( 
.A(n_11599),
.B(n_11472),
.Y(n_11759)
);

INVx1_ASAP7_75t_L g11760 ( 
.A(n_11681),
.Y(n_11760)
);

INVx3_ASAP7_75t_L g11761 ( 
.A(n_11611),
.Y(n_11761)
);

BUFx2_ASAP7_75t_SL g11762 ( 
.A(n_11609),
.Y(n_11762)
);

AND2x4_ASAP7_75t_L g11763 ( 
.A(n_11585),
.B(n_11517),
.Y(n_11763)
);

INVx3_ASAP7_75t_SL g11764 ( 
.A(n_11638),
.Y(n_11764)
);

OR2x2_ASAP7_75t_L g11765 ( 
.A(n_11601),
.B(n_11689),
.Y(n_11765)
);

INVx1_ASAP7_75t_L g11766 ( 
.A(n_11682),
.Y(n_11766)
);

INVx2_ASAP7_75t_L g11767 ( 
.A(n_11657),
.Y(n_11767)
);

NOR2xp33_ASAP7_75t_L g11768 ( 
.A(n_11685),
.B(n_11586),
.Y(n_11768)
);

INVx1_ASAP7_75t_L g11769 ( 
.A(n_11686),
.Y(n_11769)
);

AND2x2_ASAP7_75t_L g11770 ( 
.A(n_11604),
.B(n_11514),
.Y(n_11770)
);

INVx2_ASAP7_75t_L g11771 ( 
.A(n_11628),
.Y(n_11771)
);

INVx2_ASAP7_75t_SL g11772 ( 
.A(n_11590),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_11679),
.Y(n_11773)
);

INVx2_ASAP7_75t_L g11774 ( 
.A(n_11608),
.Y(n_11774)
);

NAND2xp5_ASAP7_75t_L g11775 ( 
.A(n_11661),
.B(n_11528),
.Y(n_11775)
);

NAND2xp5_ASAP7_75t_L g11776 ( 
.A(n_11664),
.B(n_11531),
.Y(n_11776)
);

AND2x2_ASAP7_75t_L g11777 ( 
.A(n_11614),
.B(n_11538),
.Y(n_11777)
);

AND2x2_ASAP7_75t_L g11778 ( 
.A(n_11640),
.B(n_11553),
.Y(n_11778)
);

INVx2_ASAP7_75t_L g11779 ( 
.A(n_11615),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_11680),
.Y(n_11780)
);

INVx2_ASAP7_75t_L g11781 ( 
.A(n_11683),
.Y(n_11781)
);

OAI21xp33_ASAP7_75t_L g11782 ( 
.A1(n_11617),
.A2(n_11440),
.B(n_11469),
.Y(n_11782)
);

HB1xp67_ASAP7_75t_L g11783 ( 
.A(n_11671),
.Y(n_11783)
);

AND2x2_ASAP7_75t_L g11784 ( 
.A(n_11736),
.B(n_11632),
.Y(n_11784)
);

OR2x6_ASAP7_75t_L g11785 ( 
.A(n_11659),
.B(n_11545),
.Y(n_11785)
);

AND2x2_ASAP7_75t_L g11786 ( 
.A(n_11626),
.B(n_11691),
.Y(n_11786)
);

OR2x2_ASAP7_75t_L g11787 ( 
.A(n_11595),
.B(n_11460),
.Y(n_11787)
);

INVx1_ASAP7_75t_L g11788 ( 
.A(n_11591),
.Y(n_11788)
);

INVx1_ASAP7_75t_L g11789 ( 
.A(n_11594),
.Y(n_11789)
);

AND2x2_ASAP7_75t_L g11790 ( 
.A(n_11718),
.B(n_11578),
.Y(n_11790)
);

INVx1_ASAP7_75t_L g11791 ( 
.A(n_11597),
.Y(n_11791)
);

AND2x2_ASAP7_75t_L g11792 ( 
.A(n_11646),
.B(n_11523),
.Y(n_11792)
);

AND2x4_ASAP7_75t_SL g11793 ( 
.A(n_11665),
.B(n_11455),
.Y(n_11793)
);

NAND2xp5_ASAP7_75t_L g11794 ( 
.A(n_11714),
.B(n_11519),
.Y(n_11794)
);

OR2x6_ASAP7_75t_L g11795 ( 
.A(n_11701),
.B(n_11562),
.Y(n_11795)
);

NAND2x1p5_ASAP7_75t_SL g11796 ( 
.A(n_11602),
.B(n_11492),
.Y(n_11796)
);

AND2x2_ASAP7_75t_L g11797 ( 
.A(n_11676),
.B(n_11559),
.Y(n_11797)
);

AND2x2_ASAP7_75t_L g11798 ( 
.A(n_11619),
.B(n_11629),
.Y(n_11798)
);

INVx1_ASAP7_75t_L g11799 ( 
.A(n_11621),
.Y(n_11799)
);

HB1xp67_ASAP7_75t_L g11800 ( 
.A(n_11699),
.Y(n_11800)
);

AND2x2_ASAP7_75t_L g11801 ( 
.A(n_11631),
.B(n_11565),
.Y(n_11801)
);

OR2x6_ASAP7_75t_SL g11802 ( 
.A(n_11600),
.B(n_11541),
.Y(n_11802)
);

AND2x2_ASAP7_75t_L g11803 ( 
.A(n_11690),
.B(n_11474),
.Y(n_11803)
);

OR2x2_ASAP7_75t_L g11804 ( 
.A(n_11622),
.B(n_11470),
.Y(n_11804)
);

NAND2x1p5_ASAP7_75t_L g11805 ( 
.A(n_11722),
.B(n_11542),
.Y(n_11805)
);

NOR2xp33_ASAP7_75t_L g11806 ( 
.A(n_11709),
.B(n_11483),
.Y(n_11806)
);

NAND2xp5_ASAP7_75t_L g11807 ( 
.A(n_11627),
.B(n_11544),
.Y(n_11807)
);

INVxp67_ASAP7_75t_L g11808 ( 
.A(n_11639),
.Y(n_11808)
);

INVx1_ASAP7_75t_L g11809 ( 
.A(n_11623),
.Y(n_11809)
);

NOR2x1_ASAP7_75t_L g11810 ( 
.A(n_11647),
.B(n_11574),
.Y(n_11810)
);

INVxp67_ASAP7_75t_SL g11811 ( 
.A(n_11715),
.Y(n_11811)
);

AND2x2_ASAP7_75t_L g11812 ( 
.A(n_11728),
.B(n_11548),
.Y(n_11812)
);

NAND2xp5_ASAP7_75t_L g11813 ( 
.A(n_11637),
.B(n_11577),
.Y(n_11813)
);

AND2x2_ASAP7_75t_L g11814 ( 
.A(n_11624),
.B(n_11456),
.Y(n_11814)
);

INVx1_ASAP7_75t_SL g11815 ( 
.A(n_11716),
.Y(n_11815)
);

INVx1_ASAP7_75t_L g11816 ( 
.A(n_11625),
.Y(n_11816)
);

INVx1_ASAP7_75t_L g11817 ( 
.A(n_11705),
.Y(n_11817)
);

AND2x2_ASAP7_75t_L g11818 ( 
.A(n_11596),
.B(n_1766),
.Y(n_11818)
);

INVx2_ASAP7_75t_L g11819 ( 
.A(n_11636),
.Y(n_11819)
);

INVx1_ASAP7_75t_L g11820 ( 
.A(n_11713),
.Y(n_11820)
);

INVx2_ASAP7_75t_L g11821 ( 
.A(n_11610),
.Y(n_11821)
);

NAND2xp5_ASAP7_75t_L g11822 ( 
.A(n_11587),
.B(n_1766),
.Y(n_11822)
);

NAND2x1p5_ASAP7_75t_L g11823 ( 
.A(n_11698),
.B(n_11721),
.Y(n_11823)
);

NAND2xp5_ASAP7_75t_SL g11824 ( 
.A(n_11644),
.B(n_1768),
.Y(n_11824)
);

OR2x2_ASAP7_75t_L g11825 ( 
.A(n_11592),
.B(n_1768),
.Y(n_11825)
);

HB1xp67_ASAP7_75t_L g11826 ( 
.A(n_11701),
.Y(n_11826)
);

INVx1_ASAP7_75t_L g11827 ( 
.A(n_11711),
.Y(n_11827)
);

OR2x2_ASAP7_75t_L g11828 ( 
.A(n_11723),
.B(n_11641),
.Y(n_11828)
);

AND2x2_ASAP7_75t_L g11829 ( 
.A(n_11630),
.B(n_1769),
.Y(n_11829)
);

BUFx2_ASAP7_75t_SL g11830 ( 
.A(n_11654),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_11717),
.B(n_1769),
.Y(n_11831)
);

NAND2xp5_ASAP7_75t_L g11832 ( 
.A(n_11645),
.B(n_1770),
.Y(n_11832)
);

AND2x2_ASAP7_75t_L g11833 ( 
.A(n_11735),
.B(n_1770),
.Y(n_11833)
);

INVx2_ASAP7_75t_L g11834 ( 
.A(n_11706),
.Y(n_11834)
);

INVx1_ASAP7_75t_L g11835 ( 
.A(n_11724),
.Y(n_11835)
);

AND2x2_ASAP7_75t_L g11836 ( 
.A(n_11729),
.B(n_1771),
.Y(n_11836)
);

AND2x2_ASAP7_75t_L g11837 ( 
.A(n_11712),
.B(n_1771),
.Y(n_11837)
);

OR2x2_ASAP7_75t_L g11838 ( 
.A(n_11688),
.B(n_1772),
.Y(n_11838)
);

AOI21xp5_ASAP7_75t_L g11839 ( 
.A1(n_11695),
.A2(n_1772),
.B(n_1773),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_11700),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_11697),
.Y(n_11841)
);

NAND2xp5_ASAP7_75t_L g11842 ( 
.A(n_11704),
.B(n_1773),
.Y(n_11842)
);

INVx1_ASAP7_75t_L g11843 ( 
.A(n_11727),
.Y(n_11843)
);

INVx1_ASAP7_75t_L g11844 ( 
.A(n_11731),
.Y(n_11844)
);

AND2x2_ASAP7_75t_L g11845 ( 
.A(n_11649),
.B(n_1774),
.Y(n_11845)
);

OR2x2_ASAP7_75t_L g11846 ( 
.A(n_11678),
.B(n_1774),
.Y(n_11846)
);

AND2x2_ASAP7_75t_L g11847 ( 
.A(n_11677),
.B(n_1775),
.Y(n_11847)
);

INVx1_ASAP7_75t_L g11848 ( 
.A(n_11696),
.Y(n_11848)
);

AND2x2_ASAP7_75t_L g11849 ( 
.A(n_11652),
.B(n_1776),
.Y(n_11849)
);

INVx1_ASAP7_75t_L g11850 ( 
.A(n_11658),
.Y(n_11850)
);

OR2x2_ASAP7_75t_L g11851 ( 
.A(n_11693),
.B(n_1776),
.Y(n_11851)
);

OR2x2_ASAP7_75t_L g11852 ( 
.A(n_11663),
.B(n_1777),
.Y(n_11852)
);

HB1xp67_ASAP7_75t_L g11853 ( 
.A(n_11635),
.Y(n_11853)
);

AND2x2_ASAP7_75t_L g11854 ( 
.A(n_11667),
.B(n_1777),
.Y(n_11854)
);

INVx3_ASAP7_75t_L g11855 ( 
.A(n_11668),
.Y(n_11855)
);

NAND4xp75_ASAP7_75t_L g11856 ( 
.A(n_11633),
.B(n_1781),
.C(n_1778),
.D(n_1780),
.Y(n_11856)
);

AND2x2_ASAP7_75t_L g11857 ( 
.A(n_11669),
.B(n_1778),
.Y(n_11857)
);

OR2x6_ASAP7_75t_L g11858 ( 
.A(n_11707),
.B(n_11653),
.Y(n_11858)
);

NAND2xp5_ASAP7_75t_L g11859 ( 
.A(n_11598),
.B(n_1781),
.Y(n_11859)
);

INVx1_ASAP7_75t_L g11860 ( 
.A(n_11703),
.Y(n_11860)
);

AND2x2_ASAP7_75t_L g11861 ( 
.A(n_11726),
.B(n_1782),
.Y(n_11861)
);

AND2x2_ASAP7_75t_L g11862 ( 
.A(n_11634),
.B(n_1782),
.Y(n_11862)
);

INVx1_ASAP7_75t_L g11863 ( 
.A(n_11675),
.Y(n_11863)
);

OR2x2_ASAP7_75t_L g11864 ( 
.A(n_11603),
.B(n_1785),
.Y(n_11864)
);

INVx1_ASAP7_75t_L g11865 ( 
.A(n_11606),
.Y(n_11865)
);

HB1xp67_ASAP7_75t_L g11866 ( 
.A(n_11655),
.Y(n_11866)
);

AND2x2_ASAP7_75t_L g11867 ( 
.A(n_11643),
.B(n_1785),
.Y(n_11867)
);

AOI22xp5_ASAP7_75t_L g11868 ( 
.A1(n_11650),
.A2(n_1788),
.B1(n_1786),
.B2(n_1787),
.Y(n_11868)
);

AND2x2_ASAP7_75t_L g11869 ( 
.A(n_11648),
.B(n_1786),
.Y(n_11869)
);

AND2x2_ASAP7_75t_L g11870 ( 
.A(n_11830),
.B(n_11734),
.Y(n_11870)
);

OAI31xp33_ASAP7_75t_L g11871 ( 
.A1(n_11751),
.A2(n_11605),
.A3(n_11656),
.B(n_11651),
.Y(n_11871)
);

CKINVDCx16_ASAP7_75t_R g11872 ( 
.A(n_11802),
.Y(n_11872)
);

AND2x2_ASAP7_75t_L g11873 ( 
.A(n_11764),
.B(n_11660),
.Y(n_11873)
);

BUFx2_ASAP7_75t_L g11874 ( 
.A(n_11750),
.Y(n_11874)
);

INVx2_ASAP7_75t_L g11875 ( 
.A(n_11761),
.Y(n_11875)
);

HB1xp67_ASAP7_75t_L g11876 ( 
.A(n_11744),
.Y(n_11876)
);

INVx1_ASAP7_75t_L g11877 ( 
.A(n_11800),
.Y(n_11877)
);

INVx1_ASAP7_75t_L g11878 ( 
.A(n_11826),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11783),
.Y(n_11879)
);

OR2x2_ASAP7_75t_L g11880 ( 
.A(n_11742),
.B(n_11662),
.Y(n_11880)
);

NAND2xp5_ASAP7_75t_L g11881 ( 
.A(n_11741),
.B(n_11702),
.Y(n_11881)
);

NAND2xp5_ASAP7_75t_L g11882 ( 
.A(n_11747),
.B(n_11733),
.Y(n_11882)
);

INVx1_ASAP7_75t_L g11883 ( 
.A(n_11817),
.Y(n_11883)
);

NOR2x1_ASAP7_75t_L g11884 ( 
.A(n_11762),
.B(n_11720),
.Y(n_11884)
);

INVx1_ASAP7_75t_L g11885 ( 
.A(n_11738),
.Y(n_11885)
);

OR2x6_ASAP7_75t_L g11886 ( 
.A(n_11767),
.B(n_11730),
.Y(n_11886)
);

INVx2_ASAP7_75t_L g11887 ( 
.A(n_11746),
.Y(n_11887)
);

AND2x2_ASAP7_75t_SL g11888 ( 
.A(n_11740),
.B(n_11710),
.Y(n_11888)
);

INVx1_ASAP7_75t_L g11889 ( 
.A(n_11752),
.Y(n_11889)
);

INVx1_ASAP7_75t_L g11890 ( 
.A(n_11755),
.Y(n_11890)
);

INVx1_ASAP7_75t_L g11891 ( 
.A(n_11774),
.Y(n_11891)
);

AND2x4_ASAP7_75t_L g11892 ( 
.A(n_11743),
.B(n_11673),
.Y(n_11892)
);

INVx2_ASAP7_75t_L g11893 ( 
.A(n_11771),
.Y(n_11893)
);

INVx1_ASAP7_75t_L g11894 ( 
.A(n_11786),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_11798),
.Y(n_11895)
);

AND2x2_ASAP7_75t_L g11896 ( 
.A(n_11759),
.B(n_11719),
.Y(n_11896)
);

INVx2_ASAP7_75t_L g11897 ( 
.A(n_11772),
.Y(n_11897)
);

INVx2_ASAP7_75t_L g11898 ( 
.A(n_11784),
.Y(n_11898)
);

INVx1_ASAP7_75t_L g11899 ( 
.A(n_11838),
.Y(n_11899)
);

AND2x2_ASAP7_75t_L g11900 ( 
.A(n_11811),
.B(n_11670),
.Y(n_11900)
);

AND2x2_ASAP7_75t_L g11901 ( 
.A(n_11745),
.B(n_11732),
.Y(n_11901)
);

NOR2xp33_ASAP7_75t_SL g11902 ( 
.A(n_11866),
.B(n_11666),
.Y(n_11902)
);

INVxp67_ASAP7_75t_L g11903 ( 
.A(n_11768),
.Y(n_11903)
);

INVx1_ASAP7_75t_L g11904 ( 
.A(n_11818),
.Y(n_11904)
);

INVx1_ASAP7_75t_L g11905 ( 
.A(n_11852),
.Y(n_11905)
);

INVx1_ASAP7_75t_L g11906 ( 
.A(n_11748),
.Y(n_11906)
);

AOI33xp33_ASAP7_75t_L g11907 ( 
.A1(n_11865),
.A2(n_11692),
.A3(n_11725),
.B1(n_11708),
.B2(n_2919),
.B3(n_2916),
.Y(n_11907)
);

OR2x2_ASAP7_75t_L g11908 ( 
.A(n_11796),
.B(n_1787),
.Y(n_11908)
);

AND2x4_ASAP7_75t_L g11909 ( 
.A(n_11756),
.B(n_1788),
.Y(n_11909)
);

OR2x2_ASAP7_75t_L g11910 ( 
.A(n_11804),
.B(n_1789),
.Y(n_11910)
);

INVx2_ASAP7_75t_L g11911 ( 
.A(n_11823),
.Y(n_11911)
);

NAND2xp5_ASAP7_75t_L g11912 ( 
.A(n_11763),
.B(n_1789),
.Y(n_11912)
);

INVx2_ASAP7_75t_SL g11913 ( 
.A(n_11855),
.Y(n_11913)
);

NAND2xp5_ASAP7_75t_L g11914 ( 
.A(n_11808),
.B(n_1790),
.Y(n_11914)
);

INVxp67_ASAP7_75t_SL g11915 ( 
.A(n_11805),
.Y(n_11915)
);

INVx1_ASAP7_75t_L g11916 ( 
.A(n_11758),
.Y(n_11916)
);

AOI22xp5_ASAP7_75t_L g11917 ( 
.A1(n_11775),
.A2(n_2902),
.B1(n_2903),
.B2(n_2901),
.Y(n_11917)
);

INVx2_ASAP7_75t_L g11918 ( 
.A(n_11760),
.Y(n_11918)
);

INVxp67_ASAP7_75t_L g11919 ( 
.A(n_11806),
.Y(n_11919)
);

INVx1_ASAP7_75t_L g11920 ( 
.A(n_11766),
.Y(n_11920)
);

NAND2xp5_ASAP7_75t_L g11921 ( 
.A(n_11753),
.B(n_1790),
.Y(n_11921)
);

NAND2xp5_ASAP7_75t_L g11922 ( 
.A(n_11778),
.B(n_1791),
.Y(n_11922)
);

INVx1_ASAP7_75t_L g11923 ( 
.A(n_11769),
.Y(n_11923)
);

BUFx3_ASAP7_75t_L g11924 ( 
.A(n_11827),
.Y(n_11924)
);

HB1xp67_ASAP7_75t_L g11925 ( 
.A(n_11785),
.Y(n_11925)
);

INVx2_ASAP7_75t_L g11926 ( 
.A(n_11781),
.Y(n_11926)
);

INVx1_ASAP7_75t_L g11927 ( 
.A(n_11829),
.Y(n_11927)
);

AND2x2_ASAP7_75t_L g11928 ( 
.A(n_11757),
.B(n_1793),
.Y(n_11928)
);

INVx1_ASAP7_75t_L g11929 ( 
.A(n_11737),
.Y(n_11929)
);

OR2x2_ASAP7_75t_L g11930 ( 
.A(n_11787),
.B(n_11828),
.Y(n_11930)
);

INVx1_ASAP7_75t_L g11931 ( 
.A(n_11833),
.Y(n_11931)
);

INVx2_ASAP7_75t_L g11932 ( 
.A(n_11821),
.Y(n_11932)
);

AOI321xp33_ASAP7_75t_L g11933 ( 
.A1(n_11807),
.A2(n_2909),
.A3(n_2906),
.B1(n_2910),
.B2(n_2908),
.C(n_2904),
.Y(n_11933)
);

INVx2_ASAP7_75t_SL g11934 ( 
.A(n_11779),
.Y(n_11934)
);

INVx1_ASAP7_75t_SL g11935 ( 
.A(n_11846),
.Y(n_11935)
);

AND2x2_ASAP7_75t_L g11936 ( 
.A(n_11739),
.B(n_1794),
.Y(n_11936)
);

OR2x2_ASAP7_75t_L g11937 ( 
.A(n_11795),
.B(n_1795),
.Y(n_11937)
);

INVx2_ASAP7_75t_SL g11938 ( 
.A(n_11836),
.Y(n_11938)
);

INVx1_ASAP7_75t_L g11939 ( 
.A(n_11837),
.Y(n_11939)
);

INVx1_ASAP7_75t_L g11940 ( 
.A(n_11847),
.Y(n_11940)
);

NAND2x1_ASAP7_75t_L g11941 ( 
.A(n_11785),
.B(n_1795),
.Y(n_11941)
);

INVx2_ASAP7_75t_L g11942 ( 
.A(n_11849),
.Y(n_11942)
);

INVx1_ASAP7_75t_L g11943 ( 
.A(n_11854),
.Y(n_11943)
);

AND2x2_ASAP7_75t_L g11944 ( 
.A(n_11777),
.B(n_1796),
.Y(n_11944)
);

AOI211xp5_ASAP7_75t_L g11945 ( 
.A1(n_11782),
.A2(n_1804),
.B(n_1813),
.C(n_1796),
.Y(n_11945)
);

INVx1_ASAP7_75t_L g11946 ( 
.A(n_11857),
.Y(n_11946)
);

INVx2_ASAP7_75t_SL g11947 ( 
.A(n_11845),
.Y(n_11947)
);

NAND2xp5_ASAP7_75t_L g11948 ( 
.A(n_11770),
.B(n_1797),
.Y(n_11948)
);

NOR3x1_ASAP7_75t_L g11949 ( 
.A(n_11776),
.B(n_11794),
.C(n_11749),
.Y(n_11949)
);

OR2x2_ASAP7_75t_L g11950 ( 
.A(n_11795),
.B(n_1797),
.Y(n_11950)
);

OR2x2_ASAP7_75t_L g11951 ( 
.A(n_11825),
.B(n_1798),
.Y(n_11951)
);

OR2x2_ASAP7_75t_L g11952 ( 
.A(n_11765),
.B(n_1798),
.Y(n_11952)
);

AND2x2_ASAP7_75t_L g11953 ( 
.A(n_11792),
.B(n_1799),
.Y(n_11953)
);

AND2x2_ASAP7_75t_L g11954 ( 
.A(n_11790),
.B(n_1799),
.Y(n_11954)
);

INVx2_ASAP7_75t_L g11955 ( 
.A(n_11861),
.Y(n_11955)
);

HB1xp67_ASAP7_75t_L g11956 ( 
.A(n_11853),
.Y(n_11956)
);

OR2x2_ASAP7_75t_L g11957 ( 
.A(n_11859),
.B(n_1800),
.Y(n_11957)
);

INVx1_ASAP7_75t_L g11958 ( 
.A(n_11862),
.Y(n_11958)
);

INVx2_ASAP7_75t_L g11959 ( 
.A(n_11819),
.Y(n_11959)
);

INVx1_ASAP7_75t_L g11960 ( 
.A(n_11867),
.Y(n_11960)
);

OR2x2_ASAP7_75t_L g11961 ( 
.A(n_11815),
.B(n_11754),
.Y(n_11961)
);

NAND2xp5_ASAP7_75t_L g11962 ( 
.A(n_11801),
.B(n_1801),
.Y(n_11962)
);

INVxp67_ASAP7_75t_SL g11963 ( 
.A(n_11822),
.Y(n_11963)
);

NAND2xp5_ASAP7_75t_L g11964 ( 
.A(n_11814),
.B(n_1802),
.Y(n_11964)
);

OR2x2_ASAP7_75t_L g11965 ( 
.A(n_11813),
.B(n_11864),
.Y(n_11965)
);

INVx1_ASAP7_75t_L g11966 ( 
.A(n_11869),
.Y(n_11966)
);

NAND2xp5_ASAP7_75t_L g11967 ( 
.A(n_11810),
.B(n_1802),
.Y(n_11967)
);

NAND2xp5_ASAP7_75t_L g11968 ( 
.A(n_11803),
.B(n_1803),
.Y(n_11968)
);

NAND2xp5_ASAP7_75t_L g11969 ( 
.A(n_11793),
.B(n_1804),
.Y(n_11969)
);

AOI21xp5_ASAP7_75t_L g11970 ( 
.A1(n_11839),
.A2(n_1805),
.B(n_1806),
.Y(n_11970)
);

INVx1_ASAP7_75t_L g11971 ( 
.A(n_11835),
.Y(n_11971)
);

INVxp67_ASAP7_75t_SL g11972 ( 
.A(n_11831),
.Y(n_11972)
);

INVx1_ASAP7_75t_L g11973 ( 
.A(n_11773),
.Y(n_11973)
);

BUFx3_ASAP7_75t_L g11974 ( 
.A(n_11780),
.Y(n_11974)
);

NAND2xp5_ASAP7_75t_L g11975 ( 
.A(n_11841),
.B(n_1805),
.Y(n_11975)
);

AND2x4_ASAP7_75t_L g11976 ( 
.A(n_11788),
.B(n_1806),
.Y(n_11976)
);

INVx1_ASAP7_75t_L g11977 ( 
.A(n_11789),
.Y(n_11977)
);

AND2x2_ASAP7_75t_L g11978 ( 
.A(n_11797),
.B(n_11820),
.Y(n_11978)
);

NAND3xp33_ASAP7_75t_L g11979 ( 
.A(n_11812),
.B(n_11824),
.C(n_11799),
.Y(n_11979)
);

INVx1_ASAP7_75t_L g11980 ( 
.A(n_11791),
.Y(n_11980)
);

AND2x2_ASAP7_75t_L g11981 ( 
.A(n_11858),
.B(n_1807),
.Y(n_11981)
);

AND2x2_ASAP7_75t_L g11982 ( 
.A(n_11858),
.B(n_1807),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_11809),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11876),
.Y(n_11984)
);

INVx2_ASAP7_75t_L g11985 ( 
.A(n_11941),
.Y(n_11985)
);

INVxp67_ASAP7_75t_SL g11986 ( 
.A(n_11956),
.Y(n_11986)
);

INVx2_ASAP7_75t_L g11987 ( 
.A(n_11874),
.Y(n_11987)
);

OAI33xp33_ASAP7_75t_L g11988 ( 
.A1(n_11879),
.A2(n_11816),
.A3(n_11863),
.B1(n_11840),
.B2(n_11848),
.B3(n_11844),
.Y(n_11988)
);

HB1xp67_ASAP7_75t_L g11989 ( 
.A(n_11925),
.Y(n_11989)
);

NOR2x1_ASAP7_75t_L g11990 ( 
.A(n_11930),
.B(n_11856),
.Y(n_11990)
);

NAND2x1p5_ASAP7_75t_L g11991 ( 
.A(n_11884),
.B(n_11870),
.Y(n_11991)
);

INVx1_ASAP7_75t_L g11992 ( 
.A(n_11937),
.Y(n_11992)
);

OAI22xp33_ASAP7_75t_L g11993 ( 
.A1(n_11872),
.A2(n_11902),
.B1(n_11908),
.B2(n_11967),
.Y(n_11993)
);

OR2x2_ASAP7_75t_L g11994 ( 
.A(n_11950),
.B(n_11834),
.Y(n_11994)
);

BUFx2_ASAP7_75t_L g11995 ( 
.A(n_11915),
.Y(n_11995)
);

INVx1_ASAP7_75t_L g11996 ( 
.A(n_11944),
.Y(n_11996)
);

NOR2xp33_ASAP7_75t_L g11997 ( 
.A(n_11875),
.B(n_11851),
.Y(n_11997)
);

INVx1_ASAP7_75t_L g11998 ( 
.A(n_11953),
.Y(n_11998)
);

BUFx3_ASAP7_75t_L g11999 ( 
.A(n_11924),
.Y(n_11999)
);

INVx2_ASAP7_75t_SL g12000 ( 
.A(n_11873),
.Y(n_12000)
);

NAND2xp5_ASAP7_75t_L g12001 ( 
.A(n_11878),
.B(n_11868),
.Y(n_12001)
);

INVx1_ASAP7_75t_L g12002 ( 
.A(n_11981),
.Y(n_12002)
);

INVx1_ASAP7_75t_L g12003 ( 
.A(n_11982),
.Y(n_12003)
);

NAND2xp5_ASAP7_75t_SL g12004 ( 
.A(n_11871),
.B(n_11843),
.Y(n_12004)
);

OAI22xp33_ASAP7_75t_SL g12005 ( 
.A1(n_11877),
.A2(n_11860),
.B1(n_11850),
.B2(n_11842),
.Y(n_12005)
);

INVx1_ASAP7_75t_L g12006 ( 
.A(n_11928),
.Y(n_12006)
);

INVx2_ASAP7_75t_L g12007 ( 
.A(n_11898),
.Y(n_12007)
);

NOR2x1p5_ASAP7_75t_SL g12008 ( 
.A(n_11961),
.B(n_11832),
.Y(n_12008)
);

INVx1_ASAP7_75t_L g12009 ( 
.A(n_11954),
.Y(n_12009)
);

OR2x2_ASAP7_75t_L g12010 ( 
.A(n_11897),
.B(n_1808),
.Y(n_12010)
);

INVx2_ASAP7_75t_L g12011 ( 
.A(n_11887),
.Y(n_12011)
);

OR2x2_ASAP7_75t_L g12012 ( 
.A(n_11893),
.B(n_1808),
.Y(n_12012)
);

OAI32xp33_ASAP7_75t_L g12013 ( 
.A1(n_11882),
.A2(n_1812),
.A3(n_1814),
.B1(n_1811),
.B2(n_1813),
.Y(n_12013)
);

NAND2xp5_ASAP7_75t_L g12014 ( 
.A(n_11888),
.B(n_1810),
.Y(n_12014)
);

NOR3xp33_ASAP7_75t_L g12015 ( 
.A(n_11979),
.B(n_1810),
.C(n_1811),
.Y(n_12015)
);

AOI32xp33_ASAP7_75t_L g12016 ( 
.A1(n_11900),
.A2(n_1815),
.A3(n_1812),
.B1(n_1814),
.B2(n_1816),
.Y(n_12016)
);

INVx1_ASAP7_75t_L g12017 ( 
.A(n_11936),
.Y(n_12017)
);

INVx2_ASAP7_75t_L g12018 ( 
.A(n_11911),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_11978),
.Y(n_12019)
);

INVx2_ASAP7_75t_SL g12020 ( 
.A(n_11974),
.Y(n_12020)
);

AOI32xp33_ASAP7_75t_L g12021 ( 
.A1(n_11896),
.A2(n_11894),
.A3(n_11895),
.B1(n_11901),
.B2(n_11891),
.Y(n_12021)
);

AOI22xp5_ASAP7_75t_L g12022 ( 
.A1(n_11903),
.A2(n_1817),
.B1(n_1815),
.B2(n_1816),
.Y(n_12022)
);

AND2x4_ASAP7_75t_L g12023 ( 
.A(n_11913),
.B(n_1817),
.Y(n_12023)
);

INVx2_ASAP7_75t_L g12024 ( 
.A(n_11951),
.Y(n_12024)
);

INVx2_ASAP7_75t_L g12025 ( 
.A(n_11880),
.Y(n_12025)
);

INVx1_ASAP7_75t_L g12026 ( 
.A(n_11969),
.Y(n_12026)
);

INVx2_ASAP7_75t_L g12027 ( 
.A(n_11909),
.Y(n_12027)
);

OR2x2_ASAP7_75t_L g12028 ( 
.A(n_11922),
.B(n_1818),
.Y(n_12028)
);

INVx1_ASAP7_75t_L g12029 ( 
.A(n_11952),
.Y(n_12029)
);

INVx1_ASAP7_75t_L g12030 ( 
.A(n_11927),
.Y(n_12030)
);

OR2x2_ASAP7_75t_L g12031 ( 
.A(n_11948),
.B(n_1819),
.Y(n_12031)
);

INVx2_ASAP7_75t_L g12032 ( 
.A(n_11947),
.Y(n_12032)
);

NAND2xp5_ASAP7_75t_L g12033 ( 
.A(n_11934),
.B(n_1820),
.Y(n_12033)
);

OAI22xp33_ASAP7_75t_L g12034 ( 
.A1(n_11881),
.A2(n_1823),
.B1(n_1820),
.B2(n_1822),
.Y(n_12034)
);

INVx1_ASAP7_75t_L g12035 ( 
.A(n_11912),
.Y(n_12035)
);

XNOR2x1_ASAP7_75t_L g12036 ( 
.A(n_11965),
.B(n_1824),
.Y(n_12036)
);

OR2x6_ASAP7_75t_L g12037 ( 
.A(n_11932),
.B(n_1822),
.Y(n_12037)
);

INVx1_ASAP7_75t_L g12038 ( 
.A(n_11910),
.Y(n_12038)
);

OAI322xp33_ASAP7_75t_L g12039 ( 
.A1(n_11889),
.A2(n_1829),
.A3(n_1828),
.B1(n_1826),
.B2(n_1824),
.C1(n_1825),
.C2(n_1827),
.Y(n_12039)
);

OR3x2_ASAP7_75t_L g12040 ( 
.A(n_11929),
.B(n_2914),
.C(n_2901),
.Y(n_12040)
);

OR2x2_ASAP7_75t_L g12041 ( 
.A(n_11964),
.B(n_1826),
.Y(n_12041)
);

A2O1A1Ixp33_ASAP7_75t_L g12042 ( 
.A1(n_11933),
.A2(n_1838),
.B(n_1847),
.C(n_1827),
.Y(n_12042)
);

INVx2_ASAP7_75t_L g12043 ( 
.A(n_11976),
.Y(n_12043)
);

OR2x2_ASAP7_75t_L g12044 ( 
.A(n_11921),
.B(n_1828),
.Y(n_12044)
);

AND2x2_ASAP7_75t_L g12045 ( 
.A(n_11942),
.B(n_11955),
.Y(n_12045)
);

OR2x2_ASAP7_75t_L g12046 ( 
.A(n_11968),
.B(n_1829),
.Y(n_12046)
);

INVx1_ASAP7_75t_L g12047 ( 
.A(n_11914),
.Y(n_12047)
);

INVx1_ASAP7_75t_L g12048 ( 
.A(n_11940),
.Y(n_12048)
);

INVx1_ASAP7_75t_L g12049 ( 
.A(n_11943),
.Y(n_12049)
);

HB1xp67_ASAP7_75t_L g12050 ( 
.A(n_11935),
.Y(n_12050)
);

HB1xp67_ASAP7_75t_L g12051 ( 
.A(n_11938),
.Y(n_12051)
);

INVx1_ASAP7_75t_L g12052 ( 
.A(n_11946),
.Y(n_12052)
);

OAI322xp33_ASAP7_75t_L g12053 ( 
.A1(n_11885),
.A2(n_1838),
.A3(n_1837),
.B1(n_1835),
.B2(n_1830),
.C1(n_1833),
.C2(n_1836),
.Y(n_12053)
);

INVx2_ASAP7_75t_SL g12054 ( 
.A(n_11892),
.Y(n_12054)
);

INVx1_ASAP7_75t_L g12055 ( 
.A(n_11958),
.Y(n_12055)
);

NOR2x1_ASAP7_75t_L g12056 ( 
.A(n_11890),
.B(n_1830),
.Y(n_12056)
);

NAND4xp75_ASAP7_75t_L g12057 ( 
.A(n_11949),
.B(n_11906),
.C(n_11920),
.D(n_11916),
.Y(n_12057)
);

O2A1O1Ixp5_ASAP7_75t_R g12058 ( 
.A1(n_11962),
.A2(n_1836),
.B(n_1833),
.C(n_1835),
.Y(n_12058)
);

NAND2xp33_ASAP7_75t_L g12059 ( 
.A(n_11959),
.B(n_1837),
.Y(n_12059)
);

INVx1_ASAP7_75t_L g12060 ( 
.A(n_11960),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11966),
.Y(n_12061)
);

AOI32xp33_ASAP7_75t_L g12062 ( 
.A1(n_11923),
.A2(n_1841),
.A3(n_1839),
.B1(n_1840),
.B2(n_1843),
.Y(n_12062)
);

OR2x2_ASAP7_75t_L g12063 ( 
.A(n_11886),
.B(n_1839),
.Y(n_12063)
);

INVx1_ASAP7_75t_L g12064 ( 
.A(n_11918),
.Y(n_12064)
);

OAI22xp33_ASAP7_75t_L g12065 ( 
.A1(n_11917),
.A2(n_1844),
.B1(n_1841),
.B2(n_1843),
.Y(n_12065)
);

OR2x2_ASAP7_75t_L g12066 ( 
.A(n_11886),
.B(n_1845),
.Y(n_12066)
);

INVx1_ASAP7_75t_L g12067 ( 
.A(n_11904),
.Y(n_12067)
);

NAND2xp5_ASAP7_75t_L g12068 ( 
.A(n_11931),
.B(n_1845),
.Y(n_12068)
);

HB1xp67_ASAP7_75t_L g12069 ( 
.A(n_11899),
.Y(n_12069)
);

NAND2xp5_ASAP7_75t_L g12070 ( 
.A(n_11939),
.B(n_1846),
.Y(n_12070)
);

INVx2_ASAP7_75t_L g12071 ( 
.A(n_11926),
.Y(n_12071)
);

OAI221xp5_ASAP7_75t_L g12072 ( 
.A1(n_11919),
.A2(n_1848),
.B1(n_1846),
.B2(n_1847),
.C(n_1849),
.Y(n_12072)
);

OAI222xp33_ASAP7_75t_L g12073 ( 
.A1(n_11971),
.A2(n_2912),
.B1(n_2908),
.B2(n_2913),
.C1(n_2911),
.C2(n_2906),
.Y(n_12073)
);

INVx1_ASAP7_75t_L g12074 ( 
.A(n_11975),
.Y(n_12074)
);

AOI22xp5_ASAP7_75t_L g12075 ( 
.A1(n_11963),
.A2(n_1850),
.B1(n_1848),
.B2(n_1849),
.Y(n_12075)
);

INVx1_ASAP7_75t_L g12076 ( 
.A(n_11883),
.Y(n_12076)
);

INVx1_ASAP7_75t_L g12077 ( 
.A(n_11905),
.Y(n_12077)
);

INVx1_ASAP7_75t_L g12078 ( 
.A(n_11973),
.Y(n_12078)
);

AND2x2_ASAP7_75t_L g12079 ( 
.A(n_11972),
.B(n_1851),
.Y(n_12079)
);

NAND2xp5_ASAP7_75t_L g12080 ( 
.A(n_11970),
.B(n_1851),
.Y(n_12080)
);

OAI21xp33_ASAP7_75t_L g12081 ( 
.A1(n_11907),
.A2(n_1852),
.B(n_1853),
.Y(n_12081)
);

INVx1_ASAP7_75t_L g12082 ( 
.A(n_11977),
.Y(n_12082)
);

INVx2_ASAP7_75t_SL g12083 ( 
.A(n_11980),
.Y(n_12083)
);

OR2x2_ASAP7_75t_L g12084 ( 
.A(n_11957),
.B(n_1853),
.Y(n_12084)
);

CKINVDCx16_ASAP7_75t_R g12085 ( 
.A(n_11983),
.Y(n_12085)
);

NAND2xp5_ASAP7_75t_SL g12086 ( 
.A(n_11945),
.B(n_1854),
.Y(n_12086)
);

INVx1_ASAP7_75t_L g12087 ( 
.A(n_11876),
.Y(n_12087)
);

AOI22xp5_ASAP7_75t_L g12088 ( 
.A1(n_11872),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.Y(n_12088)
);

OR2x2_ASAP7_75t_L g12089 ( 
.A(n_11872),
.B(n_1855),
.Y(n_12089)
);

NAND4xp75_ASAP7_75t_SL g12090 ( 
.A(n_11871),
.B(n_1858),
.C(n_1856),
.D(n_1857),
.Y(n_12090)
);

OR2x6_ASAP7_75t_L g12091 ( 
.A(n_11874),
.B(n_1858),
.Y(n_12091)
);

NAND2xp5_ASAP7_75t_L g12092 ( 
.A(n_11872),
.B(n_1859),
.Y(n_12092)
);

HB1xp67_ASAP7_75t_L g12093 ( 
.A(n_11941),
.Y(n_12093)
);

NAND2xp5_ASAP7_75t_L g12094 ( 
.A(n_11872),
.B(n_1860),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_11876),
.Y(n_12095)
);

AND2x2_ASAP7_75t_L g12096 ( 
.A(n_11874),
.B(n_1860),
.Y(n_12096)
);

OAI22xp5_ASAP7_75t_L g12097 ( 
.A1(n_11872),
.A2(n_1863),
.B1(n_1861),
.B2(n_1862),
.Y(n_12097)
);

INVx2_ASAP7_75t_SL g12098 ( 
.A(n_11941),
.Y(n_12098)
);

AOI22xp5_ASAP7_75t_L g12099 ( 
.A1(n_11872),
.A2(n_1865),
.B1(n_1863),
.B2(n_1864),
.Y(n_12099)
);

OR2x2_ASAP7_75t_L g12100 ( 
.A(n_11872),
.B(n_1864),
.Y(n_12100)
);

INVx1_ASAP7_75t_L g12101 ( 
.A(n_11876),
.Y(n_12101)
);

NAND2xp5_ASAP7_75t_L g12102 ( 
.A(n_11872),
.B(n_1865),
.Y(n_12102)
);

INVx1_ASAP7_75t_L g12103 ( 
.A(n_11876),
.Y(n_12103)
);

INVxp67_ASAP7_75t_SL g12104 ( 
.A(n_11956),
.Y(n_12104)
);

NAND2xp5_ASAP7_75t_L g12105 ( 
.A(n_11872),
.B(n_1866),
.Y(n_12105)
);

AND2x2_ASAP7_75t_L g12106 ( 
.A(n_11874),
.B(n_1867),
.Y(n_12106)
);

INVx1_ASAP7_75t_L g12107 ( 
.A(n_11876),
.Y(n_12107)
);

OR2x2_ASAP7_75t_L g12108 ( 
.A(n_11872),
.B(n_1868),
.Y(n_12108)
);

INVx1_ASAP7_75t_L g12109 ( 
.A(n_12093),
.Y(n_12109)
);

INVx1_ASAP7_75t_L g12110 ( 
.A(n_12089),
.Y(n_12110)
);

INVx2_ASAP7_75t_SL g12111 ( 
.A(n_12098),
.Y(n_12111)
);

INVx2_ASAP7_75t_L g12112 ( 
.A(n_11991),
.Y(n_12112)
);

XOR2x2_ASAP7_75t_L g12113 ( 
.A(n_12090),
.B(n_1871),
.Y(n_12113)
);

HB1xp67_ASAP7_75t_L g12114 ( 
.A(n_12091),
.Y(n_12114)
);

XNOR2xp5_ASAP7_75t_L g12115 ( 
.A(n_12036),
.B(n_1873),
.Y(n_12115)
);

BUFx2_ASAP7_75t_SL g12116 ( 
.A(n_11985),
.Y(n_12116)
);

INVx2_ASAP7_75t_L g12117 ( 
.A(n_12091),
.Y(n_12117)
);

XOR2xp5_ASAP7_75t_L g12118 ( 
.A(n_12040),
.B(n_1871),
.Y(n_12118)
);

XOR2x2_ASAP7_75t_L g12119 ( 
.A(n_11990),
.B(n_1874),
.Y(n_12119)
);

NOR2xp33_ASAP7_75t_L g12120 ( 
.A(n_12100),
.B(n_1874),
.Y(n_12120)
);

INVx2_ASAP7_75t_L g12121 ( 
.A(n_11999),
.Y(n_12121)
);

INVx2_ASAP7_75t_L g12122 ( 
.A(n_11987),
.Y(n_12122)
);

INVx2_ASAP7_75t_L g12123 ( 
.A(n_11995),
.Y(n_12123)
);

INVx1_ASAP7_75t_L g12124 ( 
.A(n_12108),
.Y(n_12124)
);

INVx1_ASAP7_75t_SL g12125 ( 
.A(n_12096),
.Y(n_12125)
);

OR2x2_ASAP7_75t_L g12126 ( 
.A(n_12092),
.B(n_1875),
.Y(n_12126)
);

INVx1_ASAP7_75t_SL g12127 ( 
.A(n_12106),
.Y(n_12127)
);

INVx2_ASAP7_75t_L g12128 ( 
.A(n_12000),
.Y(n_12128)
);

INVx2_ASAP7_75t_L g12129 ( 
.A(n_12037),
.Y(n_12129)
);

CKINVDCx14_ASAP7_75t_R g12130 ( 
.A(n_12050),
.Y(n_12130)
);

INVx2_ASAP7_75t_L g12131 ( 
.A(n_12037),
.Y(n_12131)
);

HB1xp67_ASAP7_75t_SL g12132 ( 
.A(n_12054),
.Y(n_12132)
);

INVx1_ASAP7_75t_L g12133 ( 
.A(n_11989),
.Y(n_12133)
);

XOR2x2_ASAP7_75t_L g12134 ( 
.A(n_12004),
.B(n_12057),
.Y(n_12134)
);

XNOR2xp5_ASAP7_75t_L g12135 ( 
.A(n_11993),
.B(n_1877),
.Y(n_12135)
);

INVx1_ASAP7_75t_L g12136 ( 
.A(n_11986),
.Y(n_12136)
);

NOR2xp33_ASAP7_75t_L g12137 ( 
.A(n_11984),
.B(n_12087),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_12104),
.Y(n_12138)
);

XOR2xp5_ASAP7_75t_L g12139 ( 
.A(n_12051),
.B(n_1876),
.Y(n_12139)
);

OR2x2_ASAP7_75t_L g12140 ( 
.A(n_12094),
.B(n_1876),
.Y(n_12140)
);

INVx2_ASAP7_75t_L g12141 ( 
.A(n_12063),
.Y(n_12141)
);

INVx1_ASAP7_75t_L g12142 ( 
.A(n_12102),
.Y(n_12142)
);

OAI22xp5_ASAP7_75t_SL g12143 ( 
.A1(n_12085),
.A2(n_1879),
.B1(n_1877),
.B2(n_1878),
.Y(n_12143)
);

INVx2_ASAP7_75t_L g12144 ( 
.A(n_12066),
.Y(n_12144)
);

NOR2x1_ASAP7_75t_R g12145 ( 
.A(n_12020),
.B(n_1878),
.Y(n_12145)
);

INVxp67_ASAP7_75t_L g12146 ( 
.A(n_12056),
.Y(n_12146)
);

BUFx3_ASAP7_75t_L g12147 ( 
.A(n_12095),
.Y(n_12147)
);

INVx1_ASAP7_75t_L g12148 ( 
.A(n_12105),
.Y(n_12148)
);

XOR2x2_ASAP7_75t_L g12149 ( 
.A(n_12058),
.B(n_1880),
.Y(n_12149)
);

INVx1_ASAP7_75t_L g12150 ( 
.A(n_12069),
.Y(n_12150)
);

XNOR2x1_ASAP7_75t_L g12151 ( 
.A(n_12008),
.B(n_2903),
.Y(n_12151)
);

INVx3_ASAP7_75t_L g12152 ( 
.A(n_12023),
.Y(n_12152)
);

INVx1_ASAP7_75t_L g12153 ( 
.A(n_12101),
.Y(n_12153)
);

XNOR2xp5_ASAP7_75t_L g12154 ( 
.A(n_12019),
.B(n_1881),
.Y(n_12154)
);

INVx2_ASAP7_75t_L g12155 ( 
.A(n_12103),
.Y(n_12155)
);

INVx1_ASAP7_75t_L g12156 ( 
.A(n_12107),
.Y(n_12156)
);

INVx1_ASAP7_75t_SL g12157 ( 
.A(n_11994),
.Y(n_12157)
);

AND2x2_ASAP7_75t_L g12158 ( 
.A(n_12025),
.B(n_1880),
.Y(n_12158)
);

INVx2_ASAP7_75t_L g12159 ( 
.A(n_12084),
.Y(n_12159)
);

AO22x1_ASAP7_75t_L g12160 ( 
.A1(n_12015),
.A2(n_1884),
.B1(n_1881),
.B2(n_1882),
.Y(n_12160)
);

INVxp67_ASAP7_75t_L g12161 ( 
.A(n_12014),
.Y(n_12161)
);

INVx2_ASAP7_75t_L g12162 ( 
.A(n_12028),
.Y(n_12162)
);

INVx1_ASAP7_75t_L g12163 ( 
.A(n_12006),
.Y(n_12163)
);

XNOR2x1_ASAP7_75t_L g12164 ( 
.A(n_12045),
.B(n_2912),
.Y(n_12164)
);

INVx1_ASAP7_75t_SL g12165 ( 
.A(n_12079),
.Y(n_12165)
);

BUFx3_ASAP7_75t_L g12166 ( 
.A(n_12043),
.Y(n_12166)
);

INVx1_ASAP7_75t_L g12167 ( 
.A(n_12009),
.Y(n_12167)
);

INVx1_ASAP7_75t_SL g12168 ( 
.A(n_12010),
.Y(n_12168)
);

INVx1_ASAP7_75t_L g12169 ( 
.A(n_11996),
.Y(n_12169)
);

INVx1_ASAP7_75t_L g12170 ( 
.A(n_11998),
.Y(n_12170)
);

INVx1_ASAP7_75t_L g12171 ( 
.A(n_12017),
.Y(n_12171)
);

INVx1_ASAP7_75t_L g12172 ( 
.A(n_12002),
.Y(n_12172)
);

INVxp67_ASAP7_75t_L g12173 ( 
.A(n_11997),
.Y(n_12173)
);

INVx1_ASAP7_75t_L g12174 ( 
.A(n_12003),
.Y(n_12174)
);

INVx1_ASAP7_75t_L g12175 ( 
.A(n_12012),
.Y(n_12175)
);

INVx2_ASAP7_75t_L g12176 ( 
.A(n_12046),
.Y(n_12176)
);

AND2x2_ASAP7_75t_L g12177 ( 
.A(n_12032),
.B(n_1882),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_12018),
.Y(n_12178)
);

OA22x2_ASAP7_75t_L g12179 ( 
.A1(n_11992),
.A2(n_1886),
.B1(n_1887),
.B2(n_1885),
.Y(n_12179)
);

HB1xp67_ASAP7_75t_L g12180 ( 
.A(n_12097),
.Y(n_12180)
);

NAND2xp5_ASAP7_75t_L g12181 ( 
.A(n_12042),
.B(n_1884),
.Y(n_12181)
);

AOI22xp5_ASAP7_75t_L g12182 ( 
.A1(n_12081),
.A2(n_1890),
.B1(n_1886),
.B2(n_1888),
.Y(n_12182)
);

INVxp67_ASAP7_75t_L g12183 ( 
.A(n_12059),
.Y(n_12183)
);

INVx2_ASAP7_75t_L g12184 ( 
.A(n_12031),
.Y(n_12184)
);

INVx1_ASAP7_75t_L g12185 ( 
.A(n_12033),
.Y(n_12185)
);

INVx1_ASAP7_75t_L g12186 ( 
.A(n_12007),
.Y(n_12186)
);

AO22x2_ASAP7_75t_L g12187 ( 
.A1(n_12030),
.A2(n_1892),
.B1(n_1888),
.B2(n_1891),
.Y(n_12187)
);

INVxp67_ASAP7_75t_L g12188 ( 
.A(n_12080),
.Y(n_12188)
);

INVxp67_ASAP7_75t_L g12189 ( 
.A(n_12001),
.Y(n_12189)
);

INVx2_ASAP7_75t_L g12190 ( 
.A(n_12044),
.Y(n_12190)
);

AOI22xp5_ASAP7_75t_SL g12191 ( 
.A1(n_12005),
.A2(n_12038),
.B1(n_12029),
.B2(n_12077),
.Y(n_12191)
);

INVx2_ASAP7_75t_SL g12192 ( 
.A(n_12027),
.Y(n_12192)
);

INVx1_ASAP7_75t_L g12193 ( 
.A(n_12011),
.Y(n_12193)
);

INVx2_ASAP7_75t_L g12194 ( 
.A(n_12041),
.Y(n_12194)
);

XOR2x2_ASAP7_75t_L g12195 ( 
.A(n_12086),
.B(n_1891),
.Y(n_12195)
);

NOR2xp67_ASAP7_75t_L g12196 ( 
.A(n_12083),
.B(n_1892),
.Y(n_12196)
);

HB1xp67_ASAP7_75t_L g12197 ( 
.A(n_12024),
.Y(n_12197)
);

AO22x2_ASAP7_75t_L g12198 ( 
.A1(n_12048),
.A2(n_12052),
.B1(n_12055),
.B2(n_12049),
.Y(n_12198)
);

INVx1_ASAP7_75t_L g12199 ( 
.A(n_12068),
.Y(n_12199)
);

INVx2_ASAP7_75t_L g12200 ( 
.A(n_12071),
.Y(n_12200)
);

INVx1_ASAP7_75t_L g12201 ( 
.A(n_12070),
.Y(n_12201)
);

AO22x2_ASAP7_75t_L g12202 ( 
.A1(n_12060),
.A2(n_12061),
.B1(n_12067),
.B2(n_12064),
.Y(n_12202)
);

BUFx2_ASAP7_75t_L g12203 ( 
.A(n_12076),
.Y(n_12203)
);

INVx1_ASAP7_75t_L g12204 ( 
.A(n_12088),
.Y(n_12204)
);

INVx1_ASAP7_75t_L g12205 ( 
.A(n_12099),
.Y(n_12205)
);

XNOR2x2_ASAP7_75t_L g12206 ( 
.A(n_12075),
.B(n_1893),
.Y(n_12206)
);

OAI22xp33_ASAP7_75t_SL g12207 ( 
.A1(n_12078),
.A2(n_1896),
.B1(n_1894),
.B2(n_1895),
.Y(n_12207)
);

INVx1_ASAP7_75t_L g12208 ( 
.A(n_12026),
.Y(n_12208)
);

INVx1_ASAP7_75t_L g12209 ( 
.A(n_12082),
.Y(n_12209)
);

XNOR2x1_ASAP7_75t_L g12210 ( 
.A(n_12034),
.B(n_2898),
.Y(n_12210)
);

INVxp67_ASAP7_75t_L g12211 ( 
.A(n_12072),
.Y(n_12211)
);

NOR2xp33_ASAP7_75t_L g12212 ( 
.A(n_11988),
.B(n_1896),
.Y(n_12212)
);

NAND2xp5_ASAP7_75t_L g12213 ( 
.A(n_12021),
.B(n_1897),
.Y(n_12213)
);

AOI22xp33_ASAP7_75t_L g12214 ( 
.A1(n_12035),
.A2(n_1901),
.B1(n_1898),
.B2(n_1900),
.Y(n_12214)
);

INVx1_ASAP7_75t_L g12215 ( 
.A(n_12013),
.Y(n_12215)
);

AND2x2_ASAP7_75t_L g12216 ( 
.A(n_12074),
.B(n_1898),
.Y(n_12216)
);

AND2x2_ASAP7_75t_L g12217 ( 
.A(n_12047),
.B(n_1901),
.Y(n_12217)
);

NOR2xp33_ASAP7_75t_SL g12218 ( 
.A(n_12073),
.B(n_1902),
.Y(n_12218)
);

NOR2xp33_ASAP7_75t_L g12219 ( 
.A(n_12065),
.B(n_1902),
.Y(n_12219)
);

INVx2_ASAP7_75t_L g12220 ( 
.A(n_12022),
.Y(n_12220)
);

NAND2xp33_ASAP7_75t_L g12221 ( 
.A(n_12016),
.B(n_1904),
.Y(n_12221)
);

XOR2x2_ASAP7_75t_L g12222 ( 
.A(n_12062),
.B(n_1906),
.Y(n_12222)
);

INVx2_ASAP7_75t_L g12223 ( 
.A(n_12039),
.Y(n_12223)
);

INVx1_ASAP7_75t_L g12224 ( 
.A(n_12053),
.Y(n_12224)
);

AOI22xp5_ASAP7_75t_SL g12225 ( 
.A1(n_12093),
.A2(n_1908),
.B1(n_1906),
.B2(n_1907),
.Y(n_12225)
);

INVx1_ASAP7_75t_SL g12226 ( 
.A(n_12089),
.Y(n_12226)
);

NOR2x1_ASAP7_75t_R g12227 ( 
.A(n_11995),
.B(n_1907),
.Y(n_12227)
);

INVx2_ASAP7_75t_L g12228 ( 
.A(n_12098),
.Y(n_12228)
);

AND2x2_ASAP7_75t_L g12229 ( 
.A(n_11995),
.B(n_1908),
.Y(n_12229)
);

INVx1_ASAP7_75t_L g12230 ( 
.A(n_12093),
.Y(n_12230)
);

XOR2x2_ASAP7_75t_L g12231 ( 
.A(n_12090),
.B(n_1909),
.Y(n_12231)
);

INVx1_ASAP7_75t_SL g12232 ( 
.A(n_12089),
.Y(n_12232)
);

XOR2x2_ASAP7_75t_L g12233 ( 
.A(n_12090),
.B(n_1909),
.Y(n_12233)
);

INVx2_ASAP7_75t_SL g12234 ( 
.A(n_12098),
.Y(n_12234)
);

INVx2_ASAP7_75t_L g12235 ( 
.A(n_12098),
.Y(n_12235)
);

NAND2xp5_ASAP7_75t_L g12236 ( 
.A(n_12098),
.B(n_1910),
.Y(n_12236)
);

NOR2x1_ASAP7_75t_R g12237 ( 
.A(n_11995),
.B(n_1910),
.Y(n_12237)
);

AND2x2_ASAP7_75t_L g12238 ( 
.A(n_11995),
.B(n_1911),
.Y(n_12238)
);

NOR2xp33_ASAP7_75t_L g12239 ( 
.A(n_12098),
.B(n_1911),
.Y(n_12239)
);

INVx1_ASAP7_75t_L g12240 ( 
.A(n_12093),
.Y(n_12240)
);

INVx2_ASAP7_75t_SL g12241 ( 
.A(n_12098),
.Y(n_12241)
);

XOR2x2_ASAP7_75t_L g12242 ( 
.A(n_12090),
.B(n_1912),
.Y(n_12242)
);

INVx1_ASAP7_75t_L g12243 ( 
.A(n_12093),
.Y(n_12243)
);

XOR2x2_ASAP7_75t_L g12244 ( 
.A(n_12090),
.B(n_1912),
.Y(n_12244)
);

XNOR2x1_ASAP7_75t_L g12245 ( 
.A(n_11990),
.B(n_2897),
.Y(n_12245)
);

INVx2_ASAP7_75t_L g12246 ( 
.A(n_12098),
.Y(n_12246)
);

INVxp67_ASAP7_75t_L g12247 ( 
.A(n_12093),
.Y(n_12247)
);

INVx1_ASAP7_75t_SL g12248 ( 
.A(n_12089),
.Y(n_12248)
);

INVxp67_ASAP7_75t_L g12249 ( 
.A(n_12093),
.Y(n_12249)
);

INVx2_ASAP7_75t_L g12250 ( 
.A(n_12098),
.Y(n_12250)
);

XOR2x2_ASAP7_75t_L g12251 ( 
.A(n_12090),
.B(n_1913),
.Y(n_12251)
);

XNOR2x1_ASAP7_75t_SL g12252 ( 
.A(n_11991),
.B(n_1913),
.Y(n_12252)
);

AND2x2_ASAP7_75t_L g12253 ( 
.A(n_11995),
.B(n_1914),
.Y(n_12253)
);

INVx1_ASAP7_75t_L g12254 ( 
.A(n_12093),
.Y(n_12254)
);

XOR2x2_ASAP7_75t_L g12255 ( 
.A(n_12090),
.B(n_1915),
.Y(n_12255)
);

INVx4_ASAP7_75t_L g12256 ( 
.A(n_11999),
.Y(n_12256)
);

NAND2xp5_ASAP7_75t_L g12257 ( 
.A(n_12098),
.B(n_1916),
.Y(n_12257)
);

NAND2xp5_ASAP7_75t_L g12258 ( 
.A(n_12252),
.B(n_1916),
.Y(n_12258)
);

INVx1_ASAP7_75t_L g12259 ( 
.A(n_12114),
.Y(n_12259)
);

INVx1_ASAP7_75t_L g12260 ( 
.A(n_12139),
.Y(n_12260)
);

OAI21x1_ASAP7_75t_L g12261 ( 
.A1(n_12179),
.A2(n_2904),
.B(n_2899),
.Y(n_12261)
);

INVx1_ASAP7_75t_L g12262 ( 
.A(n_12116),
.Y(n_12262)
);

INVx1_ASAP7_75t_L g12263 ( 
.A(n_12196),
.Y(n_12263)
);

AND2x2_ASAP7_75t_L g12264 ( 
.A(n_12228),
.B(n_1917),
.Y(n_12264)
);

NAND2xp5_ASAP7_75t_L g12265 ( 
.A(n_12111),
.B(n_1918),
.Y(n_12265)
);

CKINVDCx14_ASAP7_75t_R g12266 ( 
.A(n_12130),
.Y(n_12266)
);

NAND2xp5_ASAP7_75t_L g12267 ( 
.A(n_12234),
.B(n_1918),
.Y(n_12267)
);

AOI211x1_ASAP7_75t_L g12268 ( 
.A1(n_12160),
.A2(n_1922),
.B(n_1920),
.C(n_1921),
.Y(n_12268)
);

CKINVDCx16_ASAP7_75t_R g12269 ( 
.A(n_12132),
.Y(n_12269)
);

AOI22xp33_ASAP7_75t_L g12270 ( 
.A1(n_12134),
.A2(n_1922),
.B1(n_1920),
.B2(n_1921),
.Y(n_12270)
);

INVx1_ASAP7_75t_L g12271 ( 
.A(n_12229),
.Y(n_12271)
);

AOI22xp33_ASAP7_75t_L g12272 ( 
.A1(n_12123),
.A2(n_1925),
.B1(n_1923),
.B2(n_1924),
.Y(n_12272)
);

OA21x2_ASAP7_75t_L g12273 ( 
.A1(n_12212),
.A2(n_1923),
.B(n_1924),
.Y(n_12273)
);

BUFx2_ASAP7_75t_L g12274 ( 
.A(n_12146),
.Y(n_12274)
);

INVx1_ASAP7_75t_L g12275 ( 
.A(n_12238),
.Y(n_12275)
);

OR2x2_ASAP7_75t_L g12276 ( 
.A(n_12241),
.B(n_1925),
.Y(n_12276)
);

HB1xp67_ASAP7_75t_L g12277 ( 
.A(n_12151),
.Y(n_12277)
);

INVxp67_ASAP7_75t_L g12278 ( 
.A(n_12227),
.Y(n_12278)
);

AND2x2_ASAP7_75t_L g12279 ( 
.A(n_12235),
.B(n_1926),
.Y(n_12279)
);

INVx1_ASAP7_75t_L g12280 ( 
.A(n_12253),
.Y(n_12280)
);

NAND2xp5_ASAP7_75t_SL g12281 ( 
.A(n_12112),
.B(n_1926),
.Y(n_12281)
);

INVx2_ASAP7_75t_L g12282 ( 
.A(n_12166),
.Y(n_12282)
);

HB1xp67_ASAP7_75t_L g12283 ( 
.A(n_12245),
.Y(n_12283)
);

NAND2xp5_ASAP7_75t_L g12284 ( 
.A(n_12152),
.B(n_1927),
.Y(n_12284)
);

INVx1_ASAP7_75t_SL g12285 ( 
.A(n_12226),
.Y(n_12285)
);

INVxp67_ASAP7_75t_SL g12286 ( 
.A(n_12237),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_12145),
.Y(n_12287)
);

INVx1_ASAP7_75t_L g12288 ( 
.A(n_12143),
.Y(n_12288)
);

INVx1_ASAP7_75t_SL g12289 ( 
.A(n_12232),
.Y(n_12289)
);

HB1xp67_ASAP7_75t_L g12290 ( 
.A(n_12197),
.Y(n_12290)
);

INVx2_ASAP7_75t_SL g12291 ( 
.A(n_12246),
.Y(n_12291)
);

OR2x2_ASAP7_75t_L g12292 ( 
.A(n_12250),
.B(n_1927),
.Y(n_12292)
);

INVx2_ASAP7_75t_L g12293 ( 
.A(n_12256),
.Y(n_12293)
);

AOI222xp33_ASAP7_75t_L g12294 ( 
.A1(n_12213),
.A2(n_1930),
.B1(n_1932),
.B2(n_1928),
.C1(n_1929),
.C2(n_1931),
.Y(n_12294)
);

INVx1_ASAP7_75t_L g12295 ( 
.A(n_12154),
.Y(n_12295)
);

INVx3_ASAP7_75t_SL g12296 ( 
.A(n_12191),
.Y(n_12296)
);

AND2x2_ASAP7_75t_L g12297 ( 
.A(n_12248),
.B(n_1929),
.Y(n_12297)
);

AND2x2_ASAP7_75t_L g12298 ( 
.A(n_12128),
.B(n_1930),
.Y(n_12298)
);

AND2x2_ASAP7_75t_L g12299 ( 
.A(n_12125),
.B(n_12127),
.Y(n_12299)
);

NAND2xp5_ASAP7_75t_L g12300 ( 
.A(n_12225),
.B(n_1931),
.Y(n_12300)
);

INVxp67_ASAP7_75t_SL g12301 ( 
.A(n_12164),
.Y(n_12301)
);

AOI22xp33_ASAP7_75t_L g12302 ( 
.A1(n_12147),
.A2(n_1934),
.B1(n_1932),
.B2(n_1933),
.Y(n_12302)
);

NOR2x1_ASAP7_75t_L g12303 ( 
.A(n_12150),
.B(n_1933),
.Y(n_12303)
);

INVx1_ASAP7_75t_L g12304 ( 
.A(n_12187),
.Y(n_12304)
);

NAND2xp5_ASAP7_75t_L g12305 ( 
.A(n_12109),
.B(n_1934),
.Y(n_12305)
);

NOR2xp33_ASAP7_75t_L g12306 ( 
.A(n_12247),
.B(n_1935),
.Y(n_12306)
);

INVx1_ASAP7_75t_SL g12307 ( 
.A(n_12157),
.Y(n_12307)
);

INVx1_ASAP7_75t_L g12308 ( 
.A(n_12187),
.Y(n_12308)
);

INVx4_ASAP7_75t_L g12309 ( 
.A(n_12203),
.Y(n_12309)
);

NAND2xp5_ASAP7_75t_L g12310 ( 
.A(n_12230),
.B(n_1936),
.Y(n_12310)
);

INVx1_ASAP7_75t_L g12311 ( 
.A(n_12198),
.Y(n_12311)
);

NAND2xp5_ASAP7_75t_L g12312 ( 
.A(n_12240),
.B(n_1936),
.Y(n_12312)
);

NAND2xp5_ASAP7_75t_L g12313 ( 
.A(n_12243),
.B(n_1937),
.Y(n_12313)
);

OAI21xp5_ASAP7_75t_L g12314 ( 
.A1(n_12249),
.A2(n_12137),
.B(n_12133),
.Y(n_12314)
);

AND2x2_ASAP7_75t_L g12315 ( 
.A(n_12165),
.B(n_1937),
.Y(n_12315)
);

NAND2xp5_ASAP7_75t_L g12316 ( 
.A(n_12254),
.B(n_1938),
.Y(n_12316)
);

OR2x2_ASAP7_75t_L g12317 ( 
.A(n_12117),
.B(n_1939),
.Y(n_12317)
);

AND2x2_ASAP7_75t_L g12318 ( 
.A(n_12122),
.B(n_1939),
.Y(n_12318)
);

NAND2x1_ASAP7_75t_L g12319 ( 
.A(n_12136),
.B(n_1940),
.Y(n_12319)
);

OR2x2_ASAP7_75t_L g12320 ( 
.A(n_12138),
.B(n_1940),
.Y(n_12320)
);

INVx2_ASAP7_75t_L g12321 ( 
.A(n_12129),
.Y(n_12321)
);

AND2x2_ASAP7_75t_L g12322 ( 
.A(n_12110),
.B(n_1941),
.Y(n_12322)
);

INVx1_ASAP7_75t_L g12323 ( 
.A(n_12198),
.Y(n_12323)
);

NAND2xp5_ASAP7_75t_L g12324 ( 
.A(n_12192),
.B(n_1941),
.Y(n_12324)
);

INVx1_ASAP7_75t_L g12325 ( 
.A(n_12202),
.Y(n_12325)
);

INVx1_ASAP7_75t_L g12326 ( 
.A(n_12202),
.Y(n_12326)
);

INVx1_ASAP7_75t_L g12327 ( 
.A(n_12236),
.Y(n_12327)
);

NOR2x1_ASAP7_75t_R g12328 ( 
.A(n_12124),
.B(n_1942),
.Y(n_12328)
);

INVx1_ASAP7_75t_SL g12329 ( 
.A(n_12119),
.Y(n_12329)
);

INVx1_ASAP7_75t_L g12330 ( 
.A(n_12257),
.Y(n_12330)
);

AND2x2_ASAP7_75t_L g12331 ( 
.A(n_12121),
.B(n_1943),
.Y(n_12331)
);

INVxp33_ASAP7_75t_L g12332 ( 
.A(n_12118),
.Y(n_12332)
);

INVx1_ASAP7_75t_SL g12333 ( 
.A(n_12158),
.Y(n_12333)
);

INVx1_ASAP7_75t_L g12334 ( 
.A(n_12135),
.Y(n_12334)
);

AOI22xp33_ASAP7_75t_L g12335 ( 
.A1(n_12223),
.A2(n_1945),
.B1(n_1943),
.B2(n_1944),
.Y(n_12335)
);

INVx1_ASAP7_75t_L g12336 ( 
.A(n_12177),
.Y(n_12336)
);

INVx1_ASAP7_75t_L g12337 ( 
.A(n_12180),
.Y(n_12337)
);

NOR2xp33_ASAP7_75t_L g12338 ( 
.A(n_12218),
.B(n_1944),
.Y(n_12338)
);

NOR2x1_ASAP7_75t_L g12339 ( 
.A(n_12131),
.B(n_12115),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_L g12340 ( 
.A(n_12239),
.B(n_1945),
.Y(n_12340)
);

AND3x2_ASAP7_75t_L g12341 ( 
.A(n_12183),
.B(n_1948),
.C(n_1947),
.Y(n_12341)
);

AND2x2_ASAP7_75t_L g12342 ( 
.A(n_12215),
.B(n_1946),
.Y(n_12342)
);

INVx3_ASAP7_75t_L g12343 ( 
.A(n_12155),
.Y(n_12343)
);

AND2x2_ASAP7_75t_L g12344 ( 
.A(n_12159),
.B(n_1946),
.Y(n_12344)
);

INVx1_ASAP7_75t_L g12345 ( 
.A(n_12126),
.Y(n_12345)
);

INVx1_ASAP7_75t_L g12346 ( 
.A(n_12140),
.Y(n_12346)
);

OR2x2_ASAP7_75t_L g12347 ( 
.A(n_12181),
.B(n_1948),
.Y(n_12347)
);

AND2x2_ASAP7_75t_L g12348 ( 
.A(n_12141),
.B(n_1949),
.Y(n_12348)
);

INVx2_ASAP7_75t_L g12349 ( 
.A(n_12144),
.Y(n_12349)
);

NAND2xp5_ASAP7_75t_L g12350 ( 
.A(n_12224),
.B(n_1950),
.Y(n_12350)
);

INVx2_ASAP7_75t_L g12351 ( 
.A(n_12216),
.Y(n_12351)
);

INVx2_ASAP7_75t_L g12352 ( 
.A(n_12217),
.Y(n_12352)
);

INVx1_ASAP7_75t_L g12353 ( 
.A(n_12113),
.Y(n_12353)
);

AOI22xp33_ASAP7_75t_L g12354 ( 
.A1(n_12178),
.A2(n_1952),
.B1(n_1950),
.B2(n_1951),
.Y(n_12354)
);

AND2x2_ASAP7_75t_L g12355 ( 
.A(n_12163),
.B(n_1951),
.Y(n_12355)
);

NOR2xp33_ASAP7_75t_L g12356 ( 
.A(n_12168),
.B(n_1952),
.Y(n_12356)
);

INVx1_ASAP7_75t_L g12357 ( 
.A(n_12231),
.Y(n_12357)
);

NAND2xp5_ASAP7_75t_SL g12358 ( 
.A(n_12207),
.B(n_1953),
.Y(n_12358)
);

INVx2_ASAP7_75t_L g12359 ( 
.A(n_12233),
.Y(n_12359)
);

AND2x2_ASAP7_75t_L g12360 ( 
.A(n_12167),
.B(n_12169),
.Y(n_12360)
);

HB1xp67_ASAP7_75t_L g12361 ( 
.A(n_12242),
.Y(n_12361)
);

INVx1_ASAP7_75t_SL g12362 ( 
.A(n_12244),
.Y(n_12362)
);

INVx4_ASAP7_75t_L g12363 ( 
.A(n_12200),
.Y(n_12363)
);

CKINVDCx16_ASAP7_75t_R g12364 ( 
.A(n_12182),
.Y(n_12364)
);

INVxp67_ASAP7_75t_L g12365 ( 
.A(n_12120),
.Y(n_12365)
);

OR2x2_ASAP7_75t_L g12366 ( 
.A(n_12170),
.B(n_1953),
.Y(n_12366)
);

NAND2xp5_ASAP7_75t_L g12367 ( 
.A(n_12171),
.B(n_1954),
.Y(n_12367)
);

INVx1_ASAP7_75t_L g12368 ( 
.A(n_12251),
.Y(n_12368)
);

OR2x2_ASAP7_75t_L g12369 ( 
.A(n_12172),
.B(n_1954),
.Y(n_12369)
);

NAND2xp5_ASAP7_75t_L g12370 ( 
.A(n_12174),
.B(n_1955),
.Y(n_12370)
);

INVx1_ASAP7_75t_L g12371 ( 
.A(n_12255),
.Y(n_12371)
);

AND2x2_ASAP7_75t_L g12372 ( 
.A(n_12204),
.B(n_1956),
.Y(n_12372)
);

INVx1_ASAP7_75t_L g12373 ( 
.A(n_12153),
.Y(n_12373)
);

INVx1_ASAP7_75t_L g12374 ( 
.A(n_12156),
.Y(n_12374)
);

INVx4_ASAP7_75t_L g12375 ( 
.A(n_12162),
.Y(n_12375)
);

BUFx3_ASAP7_75t_L g12376 ( 
.A(n_12186),
.Y(n_12376)
);

INVx1_ASAP7_75t_L g12377 ( 
.A(n_12195),
.Y(n_12377)
);

OAI21xp5_ASAP7_75t_L g12378 ( 
.A1(n_12173),
.A2(n_1957),
.B(n_1958),
.Y(n_12378)
);

OR2x2_ASAP7_75t_L g12379 ( 
.A(n_12205),
.B(n_1957),
.Y(n_12379)
);

INVx1_ASAP7_75t_SL g12380 ( 
.A(n_12210),
.Y(n_12380)
);

NAND2xp5_ASAP7_75t_L g12381 ( 
.A(n_12175),
.B(n_1958),
.Y(n_12381)
);

INVx1_ASAP7_75t_L g12382 ( 
.A(n_12222),
.Y(n_12382)
);

BUFx3_ASAP7_75t_L g12383 ( 
.A(n_12193),
.Y(n_12383)
);

AOI22xp33_ASAP7_75t_L g12384 ( 
.A1(n_12220),
.A2(n_1961),
.B1(n_1959),
.B2(n_1960),
.Y(n_12384)
);

CKINVDCx16_ASAP7_75t_R g12385 ( 
.A(n_12142),
.Y(n_12385)
);

INVx2_ASAP7_75t_L g12386 ( 
.A(n_12176),
.Y(n_12386)
);

INVx1_ASAP7_75t_L g12387 ( 
.A(n_12206),
.Y(n_12387)
);

AND2x2_ASAP7_75t_L g12388 ( 
.A(n_12148),
.B(n_1959),
.Y(n_12388)
);

INVx1_ASAP7_75t_L g12389 ( 
.A(n_12149),
.Y(n_12389)
);

NAND2xp5_ASAP7_75t_L g12390 ( 
.A(n_12219),
.B(n_12188),
.Y(n_12390)
);

OR2x2_ASAP7_75t_L g12391 ( 
.A(n_12184),
.B(n_1960),
.Y(n_12391)
);

INVx1_ASAP7_75t_L g12392 ( 
.A(n_12221),
.Y(n_12392)
);

INVx3_ASAP7_75t_L g12393 ( 
.A(n_12190),
.Y(n_12393)
);

NOR2xp33_ASAP7_75t_L g12394 ( 
.A(n_12189),
.B(n_1961),
.Y(n_12394)
);

AND2x2_ASAP7_75t_L g12395 ( 
.A(n_12194),
.B(n_12161),
.Y(n_12395)
);

HB1xp67_ASAP7_75t_L g12396 ( 
.A(n_12209),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_12208),
.Y(n_12397)
);

INVx1_ASAP7_75t_L g12398 ( 
.A(n_12290),
.Y(n_12398)
);

AOI22xp5_ASAP7_75t_L g12399 ( 
.A1(n_12266),
.A2(n_12211),
.B1(n_12185),
.B2(n_12201),
.Y(n_12399)
);

OAI21xp33_ASAP7_75t_L g12400 ( 
.A1(n_12332),
.A2(n_12199),
.B(n_12214),
.Y(n_12400)
);

NAND2xp5_ASAP7_75t_L g12401 ( 
.A(n_12269),
.B(n_1962),
.Y(n_12401)
);

OAI21xp5_ASAP7_75t_L g12402 ( 
.A1(n_12278),
.A2(n_1964),
.B(n_1963),
.Y(n_12402)
);

AOI21xp33_ASAP7_75t_L g12403 ( 
.A1(n_12307),
.A2(n_1962),
.B(n_1963),
.Y(n_12403)
);

OR2x2_ASAP7_75t_L g12404 ( 
.A(n_12296),
.B(n_1964),
.Y(n_12404)
);

OR2x2_ASAP7_75t_L g12405 ( 
.A(n_12309),
.B(n_12258),
.Y(n_12405)
);

AOI211x1_ASAP7_75t_L g12406 ( 
.A1(n_12314),
.A2(n_1967),
.B(n_1965),
.C(n_1966),
.Y(n_12406)
);

INVx1_ASAP7_75t_L g12407 ( 
.A(n_12319),
.Y(n_12407)
);

AOI22xp5_ASAP7_75t_L g12408 ( 
.A1(n_12291),
.A2(n_1969),
.B1(n_1966),
.B2(n_1968),
.Y(n_12408)
);

AND2x2_ASAP7_75t_L g12409 ( 
.A(n_12342),
.B(n_1970),
.Y(n_12409)
);

AOI21xp5_ASAP7_75t_L g12410 ( 
.A1(n_12311),
.A2(n_1970),
.B(n_1971),
.Y(n_12410)
);

INVx1_ASAP7_75t_L g12411 ( 
.A(n_12325),
.Y(n_12411)
);

AOI221xp5_ASAP7_75t_L g12412 ( 
.A1(n_12326),
.A2(n_1973),
.B1(n_1971),
.B2(n_1972),
.C(n_1974),
.Y(n_12412)
);

INVx1_ASAP7_75t_SL g12413 ( 
.A(n_12341),
.Y(n_12413)
);

AND2x2_ASAP7_75t_L g12414 ( 
.A(n_12362),
.B(n_1972),
.Y(n_12414)
);

INVx1_ASAP7_75t_L g12415 ( 
.A(n_12323),
.Y(n_12415)
);

INVx1_ASAP7_75t_L g12416 ( 
.A(n_12303),
.Y(n_12416)
);

NOR2x1_ASAP7_75t_L g12417 ( 
.A(n_12263),
.B(n_1973),
.Y(n_12417)
);

OAI22xp5_ASAP7_75t_L g12418 ( 
.A1(n_12335),
.A2(n_1980),
.B1(n_1977),
.B2(n_1979),
.Y(n_12418)
);

INVx2_ASAP7_75t_L g12419 ( 
.A(n_12276),
.Y(n_12419)
);

AND2x4_ASAP7_75t_L g12420 ( 
.A(n_12262),
.B(n_1979),
.Y(n_12420)
);

AND2x2_ASAP7_75t_L g12421 ( 
.A(n_12359),
.B(n_1977),
.Y(n_12421)
);

BUFx2_ASAP7_75t_L g12422 ( 
.A(n_12328),
.Y(n_12422)
);

INVx1_ASAP7_75t_L g12423 ( 
.A(n_12361),
.Y(n_12423)
);

NAND2xp5_ASAP7_75t_L g12424 ( 
.A(n_12304),
.B(n_1980),
.Y(n_12424)
);

INVx2_ASAP7_75t_L g12425 ( 
.A(n_12282),
.Y(n_12425)
);

AOI221xp5_ASAP7_75t_L g12426 ( 
.A1(n_12387),
.A2(n_1983),
.B1(n_1981),
.B2(n_1982),
.C(n_1984),
.Y(n_12426)
);

AOI322xp5_ASAP7_75t_L g12427 ( 
.A1(n_12337),
.A2(n_1988),
.A3(n_1987),
.B1(n_1984),
.B2(n_1982),
.C1(n_1983),
.C2(n_1985),
.Y(n_12427)
);

AOI22xp5_ASAP7_75t_L g12428 ( 
.A1(n_12259),
.A2(n_1990),
.B1(n_1985),
.B2(n_1989),
.Y(n_12428)
);

INVx2_ASAP7_75t_L g12429 ( 
.A(n_12317),
.Y(n_12429)
);

NAND2xp5_ASAP7_75t_L g12430 ( 
.A(n_12308),
.B(n_1989),
.Y(n_12430)
);

AOI22xp5_ASAP7_75t_L g12431 ( 
.A1(n_12285),
.A2(n_1993),
.B1(n_1990),
.B2(n_1992),
.Y(n_12431)
);

AND2x2_ASAP7_75t_L g12432 ( 
.A(n_12277),
.B(n_1992),
.Y(n_12432)
);

NAND2xp5_ASAP7_75t_L g12433 ( 
.A(n_12389),
.B(n_1994),
.Y(n_12433)
);

NAND2xp5_ASAP7_75t_L g12434 ( 
.A(n_12353),
.B(n_1994),
.Y(n_12434)
);

NOR2x1_ASAP7_75t_L g12435 ( 
.A(n_12375),
.B(n_1995),
.Y(n_12435)
);

AOI22xp33_ASAP7_75t_L g12436 ( 
.A1(n_12274),
.A2(n_1997),
.B1(n_1995),
.B2(n_1996),
.Y(n_12436)
);

AOI22xp5_ASAP7_75t_L g12437 ( 
.A1(n_12289),
.A2(n_1999),
.B1(n_1996),
.B2(n_1998),
.Y(n_12437)
);

NOR2x1p5_ASAP7_75t_L g12438 ( 
.A(n_12286),
.B(n_1998),
.Y(n_12438)
);

AOI32xp33_ASAP7_75t_L g12439 ( 
.A1(n_12339),
.A2(n_2001),
.A3(n_1999),
.B1(n_2000),
.B2(n_2003),
.Y(n_12439)
);

AOI221xp5_ASAP7_75t_SL g12440 ( 
.A1(n_12329),
.A2(n_2003),
.B1(n_2000),
.B2(n_2001),
.C(n_2004),
.Y(n_12440)
);

INVxp67_ASAP7_75t_L g12441 ( 
.A(n_12338),
.Y(n_12441)
);

INVx1_ASAP7_75t_L g12442 ( 
.A(n_12283),
.Y(n_12442)
);

AOI22xp33_ASAP7_75t_L g12443 ( 
.A1(n_12321),
.A2(n_2006),
.B1(n_2004),
.B2(n_2005),
.Y(n_12443)
);

INVx1_ASAP7_75t_L g12444 ( 
.A(n_12300),
.Y(n_12444)
);

INVx1_ASAP7_75t_L g12445 ( 
.A(n_12264),
.Y(n_12445)
);

OR2x2_ASAP7_75t_L g12446 ( 
.A(n_12357),
.B(n_2005),
.Y(n_12446)
);

INVx1_ASAP7_75t_L g12447 ( 
.A(n_12279),
.Y(n_12447)
);

AOI21xp33_ASAP7_75t_L g12448 ( 
.A1(n_12368),
.A2(n_2006),
.B(n_2008),
.Y(n_12448)
);

NAND2xp5_ASAP7_75t_L g12449 ( 
.A(n_12371),
.B(n_2009),
.Y(n_12449)
);

NAND2xp5_ASAP7_75t_L g12450 ( 
.A(n_12268),
.B(n_12297),
.Y(n_12450)
);

OAI22xp33_ASAP7_75t_L g12451 ( 
.A1(n_12385),
.A2(n_2011),
.B1(n_2009),
.B2(n_2010),
.Y(n_12451)
);

INVx1_ASAP7_75t_L g12452 ( 
.A(n_12315),
.Y(n_12452)
);

NOR2xp33_ASAP7_75t_L g12453 ( 
.A(n_12363),
.B(n_2010),
.Y(n_12453)
);

NAND2xp5_ASAP7_75t_L g12454 ( 
.A(n_12318),
.B(n_2012),
.Y(n_12454)
);

OAI21xp33_ASAP7_75t_L g12455 ( 
.A1(n_12287),
.A2(n_2013),
.B(n_2014),
.Y(n_12455)
);

INVx1_ASAP7_75t_L g12456 ( 
.A(n_12320),
.Y(n_12456)
);

NAND2xp5_ASAP7_75t_L g12457 ( 
.A(n_12322),
.B(n_12288),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_12261),
.Y(n_12458)
);

AND2x2_ASAP7_75t_L g12459 ( 
.A(n_12299),
.B(n_12293),
.Y(n_12459)
);

OR2x2_ASAP7_75t_L g12460 ( 
.A(n_12265),
.B(n_2013),
.Y(n_12460)
);

AOI21xp5_ASAP7_75t_L g12461 ( 
.A1(n_12358),
.A2(n_12301),
.B(n_12281),
.Y(n_12461)
);

OAI22xp33_ASAP7_75t_L g12462 ( 
.A1(n_12364),
.A2(n_2016),
.B1(n_2014),
.B2(n_2015),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_12292),
.Y(n_12463)
);

AOI22xp5_ASAP7_75t_L g12464 ( 
.A1(n_12380),
.A2(n_2018),
.B1(n_2015),
.B2(n_2017),
.Y(n_12464)
);

NAND2xp5_ASAP7_75t_L g12465 ( 
.A(n_12298),
.B(n_2017),
.Y(n_12465)
);

INVx1_ASAP7_75t_L g12466 ( 
.A(n_12366),
.Y(n_12466)
);

AND2x2_ASAP7_75t_L g12467 ( 
.A(n_12372),
.B(n_2018),
.Y(n_12467)
);

OAI32xp33_ASAP7_75t_L g12468 ( 
.A1(n_12350),
.A2(n_2021),
.A3(n_2019),
.B1(n_2020),
.B2(n_2022),
.Y(n_12468)
);

INVx1_ASAP7_75t_L g12469 ( 
.A(n_12369),
.Y(n_12469)
);

AO21x1_ASAP7_75t_L g12470 ( 
.A1(n_12306),
.A2(n_2019),
.B(n_2020),
.Y(n_12470)
);

AOI21xp33_ASAP7_75t_SL g12471 ( 
.A1(n_12273),
.A2(n_2021),
.B(n_2022),
.Y(n_12471)
);

INVx1_ASAP7_75t_SL g12472 ( 
.A(n_12344),
.Y(n_12472)
);

NOR2xp33_ASAP7_75t_L g12473 ( 
.A(n_12343),
.B(n_2023),
.Y(n_12473)
);

AND2x4_ASAP7_75t_L g12474 ( 
.A(n_12349),
.B(n_2913),
.Y(n_12474)
);

INVx2_ASAP7_75t_SL g12475 ( 
.A(n_12331),
.Y(n_12475)
);

OAI31xp33_ASAP7_75t_L g12476 ( 
.A1(n_12396),
.A2(n_2025),
.A3(n_2023),
.B(n_2024),
.Y(n_12476)
);

NAND2xp5_ASAP7_75t_L g12477 ( 
.A(n_12348),
.B(n_2024),
.Y(n_12477)
);

AND2x2_ASAP7_75t_L g12478 ( 
.A(n_12271),
.B(n_2025),
.Y(n_12478)
);

NAND2xp5_ASAP7_75t_L g12479 ( 
.A(n_12355),
.B(n_2026),
.Y(n_12479)
);

INVx1_ASAP7_75t_L g12480 ( 
.A(n_12267),
.Y(n_12480)
);

INVxp33_ASAP7_75t_L g12481 ( 
.A(n_12356),
.Y(n_12481)
);

OAI22xp5_ASAP7_75t_L g12482 ( 
.A1(n_12270),
.A2(n_2029),
.B1(n_2027),
.B2(n_2028),
.Y(n_12482)
);

AND2x2_ASAP7_75t_L g12483 ( 
.A(n_12275),
.B(n_2027),
.Y(n_12483)
);

INVx2_ASAP7_75t_L g12484 ( 
.A(n_12391),
.Y(n_12484)
);

INVx2_ASAP7_75t_L g12485 ( 
.A(n_12379),
.Y(n_12485)
);

INVx1_ASAP7_75t_L g12486 ( 
.A(n_12284),
.Y(n_12486)
);

XOR2x2_ASAP7_75t_L g12487 ( 
.A(n_12260),
.B(n_2028),
.Y(n_12487)
);

NAND2xp5_ASAP7_75t_L g12488 ( 
.A(n_12280),
.B(n_2030),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_12324),
.Y(n_12489)
);

AO21x1_ASAP7_75t_L g12490 ( 
.A1(n_12305),
.A2(n_12312),
.B(n_12310),
.Y(n_12490)
);

NAND2xp5_ASAP7_75t_L g12491 ( 
.A(n_12393),
.B(n_2030),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_12313),
.Y(n_12492)
);

AND2x2_ASAP7_75t_L g12493 ( 
.A(n_12351),
.B(n_2031),
.Y(n_12493)
);

NAND2xp5_ASAP7_75t_L g12494 ( 
.A(n_12333),
.B(n_2031),
.Y(n_12494)
);

AND2x2_ASAP7_75t_L g12495 ( 
.A(n_12352),
.B(n_2032),
.Y(n_12495)
);

AOI22xp5_ASAP7_75t_L g12496 ( 
.A1(n_12392),
.A2(n_2036),
.B1(n_2032),
.B2(n_2034),
.Y(n_12496)
);

AOI22xp5_ASAP7_75t_L g12497 ( 
.A1(n_12382),
.A2(n_12386),
.B1(n_12295),
.B2(n_12334),
.Y(n_12497)
);

AOI321xp33_ASAP7_75t_L g12498 ( 
.A1(n_12377),
.A2(n_12395),
.A3(n_12336),
.B1(n_12360),
.B2(n_12374),
.C(n_12373),
.Y(n_12498)
);

NAND2xp5_ASAP7_75t_L g12499 ( 
.A(n_12272),
.B(n_2034),
.Y(n_12499)
);

AOI22xp5_ASAP7_75t_L g12500 ( 
.A1(n_12394),
.A2(n_2039),
.B1(n_2036),
.B2(n_2037),
.Y(n_12500)
);

AOI22xp5_ASAP7_75t_L g12501 ( 
.A1(n_12376),
.A2(n_12383),
.B1(n_12273),
.B2(n_12365),
.Y(n_12501)
);

INVx2_ASAP7_75t_L g12502 ( 
.A(n_12347),
.Y(n_12502)
);

OR2x2_ASAP7_75t_L g12503 ( 
.A(n_12316),
.B(n_2037),
.Y(n_12503)
);

INVx2_ASAP7_75t_L g12504 ( 
.A(n_12388),
.Y(n_12504)
);

AOI21xp33_ASAP7_75t_L g12505 ( 
.A1(n_12390),
.A2(n_2040),
.B(n_2041),
.Y(n_12505)
);

INVx1_ASAP7_75t_SL g12506 ( 
.A(n_12381),
.Y(n_12506)
);

INVx2_ASAP7_75t_L g12507 ( 
.A(n_12345),
.Y(n_12507)
);

AND2x2_ASAP7_75t_L g12508 ( 
.A(n_12346),
.B(n_2041),
.Y(n_12508)
);

INVx2_ASAP7_75t_SL g12509 ( 
.A(n_12397),
.Y(n_12509)
);

AOI21xp5_ASAP7_75t_L g12510 ( 
.A1(n_12340),
.A2(n_2042),
.B(n_2043),
.Y(n_12510)
);

NOR4xp25_ASAP7_75t_SL g12511 ( 
.A(n_12327),
.B(n_2047),
.C(n_2044),
.D(n_2045),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_12367),
.Y(n_12512)
);

O2A1O1Ixp33_ASAP7_75t_L g12513 ( 
.A1(n_12370),
.A2(n_2050),
.B(n_2048),
.C(n_2049),
.Y(n_12513)
);

AOI222xp33_ASAP7_75t_L g12514 ( 
.A1(n_12330),
.A2(n_2052),
.B1(n_2054),
.B2(n_2048),
.C1(n_2049),
.C2(n_2053),
.Y(n_12514)
);

AOI22xp5_ASAP7_75t_L g12515 ( 
.A1(n_12294),
.A2(n_2056),
.B1(n_2052),
.B2(n_2055),
.Y(n_12515)
);

INVx1_ASAP7_75t_SL g12516 ( 
.A(n_12378),
.Y(n_12516)
);

INVx2_ASAP7_75t_SL g12517 ( 
.A(n_12354),
.Y(n_12517)
);

NAND2xp5_ASAP7_75t_L g12518 ( 
.A(n_12384),
.B(n_2056),
.Y(n_12518)
);

INVx1_ASAP7_75t_L g12519 ( 
.A(n_12302),
.Y(n_12519)
);

INVx1_ASAP7_75t_L g12520 ( 
.A(n_12290),
.Y(n_12520)
);

NAND2xp5_ASAP7_75t_L g12521 ( 
.A(n_12266),
.B(n_2057),
.Y(n_12521)
);

AND2x2_ASAP7_75t_L g12522 ( 
.A(n_12266),
.B(n_2058),
.Y(n_12522)
);

INVx1_ASAP7_75t_L g12523 ( 
.A(n_12290),
.Y(n_12523)
);

NAND2xp5_ASAP7_75t_L g12524 ( 
.A(n_12266),
.B(n_2058),
.Y(n_12524)
);

NOR2xp33_ASAP7_75t_L g12525 ( 
.A(n_12266),
.B(n_2059),
.Y(n_12525)
);

AOI211xp5_ASAP7_75t_SL g12526 ( 
.A1(n_12290),
.A2(n_2061),
.B(n_2059),
.C(n_2060),
.Y(n_12526)
);

INVx1_ASAP7_75t_L g12527 ( 
.A(n_12290),
.Y(n_12527)
);

INVx1_ASAP7_75t_L g12528 ( 
.A(n_12290),
.Y(n_12528)
);

AOI22xp5_ASAP7_75t_L g12529 ( 
.A1(n_12266),
.A2(n_2063),
.B1(n_2061),
.B2(n_2062),
.Y(n_12529)
);

INVx1_ASAP7_75t_L g12530 ( 
.A(n_12522),
.Y(n_12530)
);

INVx1_ASAP7_75t_L g12531 ( 
.A(n_12404),
.Y(n_12531)
);

NAND2xp5_ASAP7_75t_L g12532 ( 
.A(n_12526),
.B(n_2064),
.Y(n_12532)
);

AOI221x1_ASAP7_75t_L g12533 ( 
.A1(n_12471),
.A2(n_12415),
.B1(n_12411),
.B2(n_12400),
.C(n_12461),
.Y(n_12533)
);

AOI21xp33_ASAP7_75t_L g12534 ( 
.A1(n_12407),
.A2(n_2065),
.B(n_2066),
.Y(n_12534)
);

OAI21xp5_ASAP7_75t_SL g12535 ( 
.A1(n_12501),
.A2(n_2067),
.B(n_2066),
.Y(n_12535)
);

INVxp67_ASAP7_75t_SL g12536 ( 
.A(n_12435),
.Y(n_12536)
);

INVx1_ASAP7_75t_L g12537 ( 
.A(n_12521),
.Y(n_12537)
);

OAI32xp33_ASAP7_75t_L g12538 ( 
.A1(n_12413),
.A2(n_2068),
.A3(n_2065),
.B1(n_2067),
.B2(n_2069),
.Y(n_12538)
);

INVx1_ASAP7_75t_L g12539 ( 
.A(n_12524),
.Y(n_12539)
);

AOI22xp5_ASAP7_75t_L g12540 ( 
.A1(n_12423),
.A2(n_2070),
.B1(n_2068),
.B2(n_2069),
.Y(n_12540)
);

NAND2xp5_ASAP7_75t_L g12541 ( 
.A(n_12414),
.B(n_2070),
.Y(n_12541)
);

AOI22xp33_ASAP7_75t_L g12542 ( 
.A1(n_12398),
.A2(n_2073),
.B1(n_2071),
.B2(n_2072),
.Y(n_12542)
);

AOI22xp5_ASAP7_75t_L g12543 ( 
.A1(n_12442),
.A2(n_2074),
.B1(n_2071),
.B2(n_2073),
.Y(n_12543)
);

AOI22xp5_ASAP7_75t_L g12544 ( 
.A1(n_12525),
.A2(n_2076),
.B1(n_2074),
.B2(n_2075),
.Y(n_12544)
);

AND2x2_ASAP7_75t_L g12545 ( 
.A(n_12421),
.B(n_2076),
.Y(n_12545)
);

OAI22xp5_ASAP7_75t_L g12546 ( 
.A1(n_12520),
.A2(n_2079),
.B1(n_2077),
.B2(n_2078),
.Y(n_12546)
);

OAI21xp33_ASAP7_75t_L g12547 ( 
.A1(n_12497),
.A2(n_2917),
.B(n_2915),
.Y(n_12547)
);

AOI22xp33_ASAP7_75t_L g12548 ( 
.A1(n_12523),
.A2(n_2079),
.B1(n_2077),
.B2(n_2078),
.Y(n_12548)
);

NAND2xp5_ASAP7_75t_L g12549 ( 
.A(n_12432),
.B(n_2080),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_12459),
.B(n_2080),
.Y(n_12550)
);

NOR3xp33_ASAP7_75t_L g12551 ( 
.A(n_12434),
.B(n_12449),
.C(n_12433),
.Y(n_12551)
);

NAND2xp5_ASAP7_75t_L g12552 ( 
.A(n_12409),
.B(n_2081),
.Y(n_12552)
);

INVx1_ASAP7_75t_L g12553 ( 
.A(n_12401),
.Y(n_12553)
);

OAI22xp33_ASAP7_75t_SL g12554 ( 
.A1(n_12416),
.A2(n_2083),
.B1(n_2081),
.B2(n_2082),
.Y(n_12554)
);

OAI22xp33_ASAP7_75t_SL g12555 ( 
.A1(n_12527),
.A2(n_2084),
.B1(n_2082),
.B2(n_2083),
.Y(n_12555)
);

NAND2xp33_ASAP7_75t_L g12556 ( 
.A(n_12417),
.B(n_2084),
.Y(n_12556)
);

OR2x2_ASAP7_75t_L g12557 ( 
.A(n_12446),
.B(n_2085),
.Y(n_12557)
);

INVx1_ASAP7_75t_L g12558 ( 
.A(n_12470),
.Y(n_12558)
);

AOI22x1_ASAP7_75t_SL g12559 ( 
.A1(n_12452),
.A2(n_2088),
.B1(n_2086),
.B2(n_2087),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_12474),
.B(n_2086),
.Y(n_12560)
);

O2A1O1Ixp33_ASAP7_75t_L g12561 ( 
.A1(n_12528),
.A2(n_2091),
.B(n_2088),
.C(n_2090),
.Y(n_12561)
);

INVx1_ASAP7_75t_L g12562 ( 
.A(n_12420),
.Y(n_12562)
);

INVxp67_ASAP7_75t_SL g12563 ( 
.A(n_12438),
.Y(n_12563)
);

AND2x2_ASAP7_75t_L g12564 ( 
.A(n_12422),
.B(n_2090),
.Y(n_12564)
);

INVx2_ASAP7_75t_L g12565 ( 
.A(n_12420),
.Y(n_12565)
);

NAND4xp75_ASAP7_75t_L g12566 ( 
.A(n_12406),
.B(n_2093),
.C(n_2091),
.D(n_2092),
.Y(n_12566)
);

AOI22xp5_ASAP7_75t_L g12567 ( 
.A1(n_12425),
.A2(n_2094),
.B1(n_2092),
.B2(n_2093),
.Y(n_12567)
);

INVx1_ASAP7_75t_L g12568 ( 
.A(n_12478),
.Y(n_12568)
);

OR2x2_ASAP7_75t_L g12569 ( 
.A(n_12405),
.B(n_2094),
.Y(n_12569)
);

NOR2xp33_ASAP7_75t_L g12570 ( 
.A(n_12455),
.B(n_2095),
.Y(n_12570)
);

AOI22xp5_ASAP7_75t_L g12571 ( 
.A1(n_12517),
.A2(n_2097),
.B1(n_2095),
.B2(n_2096),
.Y(n_12571)
);

INVx1_ASAP7_75t_L g12572 ( 
.A(n_12483),
.Y(n_12572)
);

OAI21xp33_ASAP7_75t_SL g12573 ( 
.A1(n_12458),
.A2(n_2098),
.B(n_2100),
.Y(n_12573)
);

AND2x2_ASAP7_75t_L g12574 ( 
.A(n_12467),
.B(n_12493),
.Y(n_12574)
);

INVx1_ASAP7_75t_L g12575 ( 
.A(n_12487),
.Y(n_12575)
);

INVx1_ASAP7_75t_L g12576 ( 
.A(n_12508),
.Y(n_12576)
);

OAI221xp5_ASAP7_75t_L g12577 ( 
.A1(n_12439),
.A2(n_2102),
.B1(n_2098),
.B2(n_2101),
.C(n_2103),
.Y(n_12577)
);

OAI21xp5_ASAP7_75t_L g12578 ( 
.A1(n_12399),
.A2(n_2101),
.B(n_2102),
.Y(n_12578)
);

OAI21xp5_ASAP7_75t_SL g12579 ( 
.A1(n_12515),
.A2(n_2106),
.B(n_2105),
.Y(n_12579)
);

INVx2_ASAP7_75t_L g12580 ( 
.A(n_12460),
.Y(n_12580)
);

INVx1_ASAP7_75t_L g12581 ( 
.A(n_12424),
.Y(n_12581)
);

OAI22xp5_ASAP7_75t_L g12582 ( 
.A1(n_12431),
.A2(n_2106),
.B1(n_2104),
.B2(n_2105),
.Y(n_12582)
);

OR2x2_ASAP7_75t_L g12583 ( 
.A(n_12450),
.B(n_2107),
.Y(n_12583)
);

OAI22xp33_ASAP7_75t_L g12584 ( 
.A1(n_12481),
.A2(n_2110),
.B1(n_2107),
.B2(n_2108),
.Y(n_12584)
);

OR2x2_ASAP7_75t_L g12585 ( 
.A(n_12491),
.B(n_2108),
.Y(n_12585)
);

AOI22xp33_ASAP7_75t_L g12586 ( 
.A1(n_12507),
.A2(n_2113),
.B1(n_2110),
.B2(n_2111),
.Y(n_12586)
);

NAND2xp5_ASAP7_75t_L g12587 ( 
.A(n_12440),
.B(n_2114),
.Y(n_12587)
);

NAND3xp33_ASAP7_75t_L g12588 ( 
.A(n_12498),
.B(n_2114),
.C(n_2115),
.Y(n_12588)
);

OR2x2_ASAP7_75t_L g12589 ( 
.A(n_12494),
.B(n_2115),
.Y(n_12589)
);

OA21x2_ASAP7_75t_L g12590 ( 
.A1(n_12457),
.A2(n_2116),
.B(n_2117),
.Y(n_12590)
);

NAND4xp25_ASAP7_75t_L g12591 ( 
.A(n_12519),
.B(n_12516),
.C(n_12472),
.D(n_12445),
.Y(n_12591)
);

OAI22xp5_ASAP7_75t_L g12592 ( 
.A1(n_12437),
.A2(n_2119),
.B1(n_2117),
.B2(n_2118),
.Y(n_12592)
);

NAND2xp5_ASAP7_75t_SL g12593 ( 
.A(n_12462),
.B(n_2118),
.Y(n_12593)
);

INVx1_ASAP7_75t_SL g12594 ( 
.A(n_12495),
.Y(n_12594)
);

INVx1_ASAP7_75t_L g12595 ( 
.A(n_12430),
.Y(n_12595)
);

AND2x2_ASAP7_75t_L g12596 ( 
.A(n_12419),
.B(n_12504),
.Y(n_12596)
);

AOI31xp33_ASAP7_75t_L g12597 ( 
.A1(n_12447),
.A2(n_2121),
.A3(n_2119),
.B(n_2120),
.Y(n_12597)
);

AOI22xp5_ASAP7_75t_L g12598 ( 
.A1(n_12475),
.A2(n_2122),
.B1(n_2120),
.B2(n_2121),
.Y(n_12598)
);

INVx1_ASAP7_75t_L g12599 ( 
.A(n_12479),
.Y(n_12599)
);

A2O1A1Ixp33_ASAP7_75t_L g12600 ( 
.A1(n_12473),
.A2(n_2125),
.B(n_2123),
.C(n_2124),
.Y(n_12600)
);

AOI22xp5_ASAP7_75t_L g12601 ( 
.A1(n_12509),
.A2(n_2128),
.B1(n_2125),
.B2(n_2127),
.Y(n_12601)
);

INVx1_ASAP7_75t_L g12602 ( 
.A(n_12465),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_12477),
.Y(n_12603)
);

INVx1_ASAP7_75t_L g12604 ( 
.A(n_12454),
.Y(n_12604)
);

INVx1_ASAP7_75t_L g12605 ( 
.A(n_12488),
.Y(n_12605)
);

NAND2xp5_ASAP7_75t_L g12606 ( 
.A(n_12410),
.B(n_2127),
.Y(n_12606)
);

AOI22xp5_ASAP7_75t_L g12607 ( 
.A1(n_12441),
.A2(n_2130),
.B1(n_2128),
.B2(n_2129),
.Y(n_12607)
);

OAI21xp5_ASAP7_75t_SL g12608 ( 
.A1(n_12506),
.A2(n_2131),
.B(n_2130),
.Y(n_12608)
);

INVx1_ASAP7_75t_L g12609 ( 
.A(n_12529),
.Y(n_12609)
);

AOI21xp5_ASAP7_75t_L g12610 ( 
.A1(n_12513),
.A2(n_2129),
.B(n_2133),
.Y(n_12610)
);

XNOR2x1_ASAP7_75t_L g12611 ( 
.A(n_12482),
.B(n_2133),
.Y(n_12611)
);

OAI221xp5_ASAP7_75t_L g12612 ( 
.A1(n_12476),
.A2(n_2138),
.B1(n_2134),
.B2(n_2136),
.C(n_2141),
.Y(n_12612)
);

AOI321xp33_ASAP7_75t_L g12613 ( 
.A1(n_12444),
.A2(n_2141),
.A3(n_2143),
.B1(n_2134),
.B2(n_2138),
.C(n_2142),
.Y(n_12613)
);

AND2x2_ASAP7_75t_L g12614 ( 
.A(n_12429),
.B(n_2144),
.Y(n_12614)
);

AND2x2_ASAP7_75t_L g12615 ( 
.A(n_12485),
.B(n_2144),
.Y(n_12615)
);

AO22x1_ASAP7_75t_L g12616 ( 
.A1(n_12453),
.A2(n_2147),
.B1(n_2145),
.B2(n_2146),
.Y(n_12616)
);

NOR2xp33_ASAP7_75t_L g12617 ( 
.A(n_12448),
.B(n_12403),
.Y(n_12617)
);

AOI221xp5_ASAP7_75t_L g12618 ( 
.A1(n_12456),
.A2(n_2147),
.B1(n_2145),
.B2(n_2146),
.C(n_2149),
.Y(n_12618)
);

OAI22xp5_ASAP7_75t_L g12619 ( 
.A1(n_12464),
.A2(n_2152),
.B1(n_2150),
.B2(n_2151),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_12499),
.Y(n_12620)
);

INVx2_ASAP7_75t_L g12621 ( 
.A(n_12503),
.Y(n_12621)
);

AOI22xp5_ASAP7_75t_L g12622 ( 
.A1(n_12418),
.A2(n_2153),
.B1(n_2150),
.B2(n_2152),
.Y(n_12622)
);

AOI22xp5_ASAP7_75t_L g12623 ( 
.A1(n_12463),
.A2(n_2155),
.B1(n_2153),
.B2(n_2154),
.Y(n_12623)
);

INVx1_ASAP7_75t_L g12624 ( 
.A(n_12518),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12466),
.Y(n_12625)
);

AOI21xp5_ASAP7_75t_L g12626 ( 
.A1(n_12510),
.A2(n_2154),
.B(n_2156),
.Y(n_12626)
);

NOR2x1_ASAP7_75t_L g12627 ( 
.A(n_12451),
.B(n_2156),
.Y(n_12627)
);

OAI22xp33_ASAP7_75t_SL g12628 ( 
.A1(n_12469),
.A2(n_2159),
.B1(n_2157),
.B2(n_2158),
.Y(n_12628)
);

OAI21xp5_ASAP7_75t_SL g12629 ( 
.A1(n_12426),
.A2(n_2159),
.B(n_2158),
.Y(n_12629)
);

XNOR2xp5_ASAP7_75t_L g12630 ( 
.A(n_12496),
.B(n_2157),
.Y(n_12630)
);

AOI21xp33_ASAP7_75t_SL g12631 ( 
.A1(n_12505),
.A2(n_2160),
.B(n_2162),
.Y(n_12631)
);

INVxp67_ASAP7_75t_L g12632 ( 
.A(n_12514),
.Y(n_12632)
);

INVxp33_ASAP7_75t_L g12633 ( 
.A(n_12484),
.Y(n_12633)
);

AND2x2_ASAP7_75t_L g12634 ( 
.A(n_12511),
.B(n_2160),
.Y(n_12634)
);

OAI22xp5_ASAP7_75t_L g12635 ( 
.A1(n_12436),
.A2(n_2164),
.B1(n_2162),
.B2(n_2163),
.Y(n_12635)
);

NAND2xp5_ASAP7_75t_L g12636 ( 
.A(n_12428),
.B(n_2163),
.Y(n_12636)
);

INVx1_ASAP7_75t_L g12637 ( 
.A(n_12402),
.Y(n_12637)
);

NOR2xp33_ASAP7_75t_L g12638 ( 
.A(n_12468),
.B(n_2165),
.Y(n_12638)
);

NAND2xp5_ASAP7_75t_L g12639 ( 
.A(n_12412),
.B(n_12427),
.Y(n_12639)
);

NAND2xp5_ASAP7_75t_L g12640 ( 
.A(n_12443),
.B(n_2165),
.Y(n_12640)
);

INVx2_ASAP7_75t_L g12641 ( 
.A(n_12502),
.Y(n_12641)
);

AND2x2_ASAP7_75t_L g12642 ( 
.A(n_12486),
.B(n_2166),
.Y(n_12642)
);

OAI211xp5_ASAP7_75t_L g12643 ( 
.A1(n_12480),
.A2(n_2168),
.B(n_2166),
.C(n_2167),
.Y(n_12643)
);

INVx1_ASAP7_75t_L g12644 ( 
.A(n_12490),
.Y(n_12644)
);

NOR2xp33_ASAP7_75t_L g12645 ( 
.A(n_12489),
.B(n_2167),
.Y(n_12645)
);

AND2x2_ASAP7_75t_L g12646 ( 
.A(n_12492),
.B(n_2168),
.Y(n_12646)
);

NAND2xp5_ASAP7_75t_L g12647 ( 
.A(n_12408),
.B(n_2170),
.Y(n_12647)
);

AOI21xp5_ASAP7_75t_L g12648 ( 
.A1(n_12512),
.A2(n_2171),
.B(n_2173),
.Y(n_12648)
);

AOI21xp33_ASAP7_75t_SL g12649 ( 
.A1(n_12500),
.A2(n_2171),
.B(n_2174),
.Y(n_12649)
);

NOR2xp33_ASAP7_75t_L g12650 ( 
.A(n_12562),
.B(n_2174),
.Y(n_12650)
);

NOR2xp33_ASAP7_75t_L g12651 ( 
.A(n_12565),
.B(n_2175),
.Y(n_12651)
);

AND2x2_ASAP7_75t_L g12652 ( 
.A(n_12564),
.B(n_2175),
.Y(n_12652)
);

NAND2xp33_ASAP7_75t_L g12653 ( 
.A(n_12634),
.B(n_2176),
.Y(n_12653)
);

NAND2xp5_ASAP7_75t_SL g12654 ( 
.A(n_12554),
.B(n_2176),
.Y(n_12654)
);

NAND2xp5_ASAP7_75t_L g12655 ( 
.A(n_12616),
.B(n_12550),
.Y(n_12655)
);

NAND2xp5_ASAP7_75t_L g12656 ( 
.A(n_12615),
.B(n_2177),
.Y(n_12656)
);

INVx2_ASAP7_75t_L g12657 ( 
.A(n_12590),
.Y(n_12657)
);

INVx2_ASAP7_75t_L g12658 ( 
.A(n_12590),
.Y(n_12658)
);

OAI222xp33_ASAP7_75t_L g12659 ( 
.A1(n_12558),
.A2(n_2180),
.B1(n_2183),
.B2(n_2178),
.C1(n_2179),
.C2(n_2182),
.Y(n_12659)
);

NAND2xp5_ASAP7_75t_L g12660 ( 
.A(n_12545),
.B(n_2178),
.Y(n_12660)
);

NAND2xp5_ASAP7_75t_L g12661 ( 
.A(n_12614),
.B(n_2179),
.Y(n_12661)
);

AOI22xp33_ASAP7_75t_L g12662 ( 
.A1(n_12588),
.A2(n_2183),
.B1(n_2180),
.B2(n_2182),
.Y(n_12662)
);

INVx1_ASAP7_75t_L g12663 ( 
.A(n_12559),
.Y(n_12663)
);

CKINVDCx20_ASAP7_75t_R g12664 ( 
.A(n_12575),
.Y(n_12664)
);

NOR2xp33_ASAP7_75t_L g12665 ( 
.A(n_12633),
.B(n_2184),
.Y(n_12665)
);

AND2x4_ASAP7_75t_L g12666 ( 
.A(n_12536),
.B(n_2184),
.Y(n_12666)
);

AND2x2_ASAP7_75t_L g12667 ( 
.A(n_12574),
.B(n_2185),
.Y(n_12667)
);

AOI22xp33_ASAP7_75t_L g12668 ( 
.A1(n_12641),
.A2(n_2188),
.B1(n_2185),
.B2(n_2186),
.Y(n_12668)
);

BUFx2_ASAP7_75t_L g12669 ( 
.A(n_12573),
.Y(n_12669)
);

NOR2xp67_ASAP7_75t_L g12670 ( 
.A(n_12643),
.B(n_2189),
.Y(n_12670)
);

INVx1_ASAP7_75t_SL g12671 ( 
.A(n_12557),
.Y(n_12671)
);

NAND2xp5_ASAP7_75t_L g12672 ( 
.A(n_12597),
.B(n_2188),
.Y(n_12672)
);

INVx1_ASAP7_75t_L g12673 ( 
.A(n_12532),
.Y(n_12673)
);

OAI21xp5_ASAP7_75t_SL g12674 ( 
.A1(n_12535),
.A2(n_2189),
.B(n_2190),
.Y(n_12674)
);

OR2x2_ASAP7_75t_L g12675 ( 
.A(n_12583),
.B(n_2190),
.Y(n_12675)
);

INVxp67_ASAP7_75t_L g12676 ( 
.A(n_12645),
.Y(n_12676)
);

INVx1_ASAP7_75t_L g12677 ( 
.A(n_12569),
.Y(n_12677)
);

NAND2xp5_ASAP7_75t_L g12678 ( 
.A(n_12563),
.B(n_2191),
.Y(n_12678)
);

NAND2xp5_ASAP7_75t_L g12679 ( 
.A(n_12530),
.B(n_2191),
.Y(n_12679)
);

NAND2xp5_ASAP7_75t_L g12680 ( 
.A(n_12642),
.B(n_2192),
.Y(n_12680)
);

HB1xp67_ASAP7_75t_L g12681 ( 
.A(n_12566),
.Y(n_12681)
);

INVx1_ASAP7_75t_L g12682 ( 
.A(n_12549),
.Y(n_12682)
);

NAND2xp5_ASAP7_75t_L g12683 ( 
.A(n_12646),
.B(n_2192),
.Y(n_12683)
);

INVx1_ASAP7_75t_L g12684 ( 
.A(n_12552),
.Y(n_12684)
);

OR2x2_ASAP7_75t_L g12685 ( 
.A(n_12587),
.B(n_2193),
.Y(n_12685)
);

INVx1_ASAP7_75t_L g12686 ( 
.A(n_12556),
.Y(n_12686)
);

NAND2xp5_ASAP7_75t_L g12687 ( 
.A(n_12555),
.B(n_2195),
.Y(n_12687)
);

NAND3xp33_ASAP7_75t_SL g12688 ( 
.A(n_12608),
.B(n_2196),
.C(n_2197),
.Y(n_12688)
);

INVx2_ASAP7_75t_L g12689 ( 
.A(n_12589),
.Y(n_12689)
);

NAND2xp5_ASAP7_75t_SL g12690 ( 
.A(n_12628),
.B(n_2196),
.Y(n_12690)
);

NAND2xp5_ASAP7_75t_L g12691 ( 
.A(n_12531),
.B(n_2197),
.Y(n_12691)
);

OAI21xp33_ASAP7_75t_L g12692 ( 
.A1(n_12591),
.A2(n_2198),
.B(n_2199),
.Y(n_12692)
);

INVx1_ASAP7_75t_L g12693 ( 
.A(n_12541),
.Y(n_12693)
);

NAND2xp5_ASAP7_75t_L g12694 ( 
.A(n_12648),
.B(n_2198),
.Y(n_12694)
);

NAND2xp5_ASAP7_75t_L g12695 ( 
.A(n_12540),
.B(n_2200),
.Y(n_12695)
);

HB1xp67_ASAP7_75t_L g12696 ( 
.A(n_12627),
.Y(n_12696)
);

OAI22xp5_ASAP7_75t_L g12697 ( 
.A1(n_12571),
.A2(n_12632),
.B1(n_12622),
.B2(n_12577),
.Y(n_12697)
);

INVx2_ASAP7_75t_L g12698 ( 
.A(n_12585),
.Y(n_12698)
);

INVxp67_ASAP7_75t_L g12699 ( 
.A(n_12638),
.Y(n_12699)
);

NAND2xp5_ASAP7_75t_L g12700 ( 
.A(n_12543),
.B(n_2200),
.Y(n_12700)
);

INVx1_ASAP7_75t_L g12701 ( 
.A(n_12560),
.Y(n_12701)
);

AND2x2_ASAP7_75t_L g12702 ( 
.A(n_12596),
.B(n_2201),
.Y(n_12702)
);

AOI22xp33_ASAP7_75t_L g12703 ( 
.A1(n_12625),
.A2(n_2204),
.B1(n_2201),
.B2(n_2202),
.Y(n_12703)
);

INVx2_ASAP7_75t_L g12704 ( 
.A(n_12611),
.Y(n_12704)
);

INVx1_ASAP7_75t_L g12705 ( 
.A(n_12606),
.Y(n_12705)
);

NAND2xp5_ASAP7_75t_L g12706 ( 
.A(n_12542),
.B(n_2202),
.Y(n_12706)
);

AND2x2_ASAP7_75t_L g12707 ( 
.A(n_12568),
.B(n_2204),
.Y(n_12707)
);

INVx3_ASAP7_75t_L g12708 ( 
.A(n_12580),
.Y(n_12708)
);

NAND2xp5_ASAP7_75t_L g12709 ( 
.A(n_12548),
.B(n_2205),
.Y(n_12709)
);

OR2x2_ASAP7_75t_L g12710 ( 
.A(n_12594),
.B(n_12572),
.Y(n_12710)
);

AND2x2_ASAP7_75t_L g12711 ( 
.A(n_12576),
.B(n_2205),
.Y(n_12711)
);

INVx2_ASAP7_75t_L g12712 ( 
.A(n_12621),
.Y(n_12712)
);

AND2x2_ASAP7_75t_L g12713 ( 
.A(n_12609),
.B(n_2206),
.Y(n_12713)
);

NOR2xp33_ASAP7_75t_L g12714 ( 
.A(n_12547),
.B(n_2206),
.Y(n_12714)
);

NAND2xp5_ASAP7_75t_L g12715 ( 
.A(n_12601),
.B(n_2207),
.Y(n_12715)
);

AND2x2_ASAP7_75t_L g12716 ( 
.A(n_12578),
.B(n_2208),
.Y(n_12716)
);

NOR2xp33_ASAP7_75t_L g12717 ( 
.A(n_12612),
.B(n_2208),
.Y(n_12717)
);

NOR2xp33_ASAP7_75t_L g12718 ( 
.A(n_12579),
.B(n_2210),
.Y(n_12718)
);

NOR2xp33_ASAP7_75t_L g12719 ( 
.A(n_12649),
.B(n_2210),
.Y(n_12719)
);

NAND2xp5_ASAP7_75t_L g12720 ( 
.A(n_12644),
.B(n_2211),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_12598),
.B(n_2211),
.Y(n_12721)
);

NOR2xp33_ASAP7_75t_L g12722 ( 
.A(n_12534),
.B(n_2212),
.Y(n_12722)
);

NOR2xp33_ASAP7_75t_L g12723 ( 
.A(n_12631),
.B(n_2213),
.Y(n_12723)
);

NAND2xp5_ASAP7_75t_L g12724 ( 
.A(n_12584),
.B(n_2213),
.Y(n_12724)
);

INVx1_ASAP7_75t_L g12725 ( 
.A(n_12640),
.Y(n_12725)
);

AND2x4_ASAP7_75t_SL g12726 ( 
.A(n_12537),
.B(n_2214),
.Y(n_12726)
);

NOR2x1_ASAP7_75t_L g12727 ( 
.A(n_12600),
.B(n_2215),
.Y(n_12727)
);

AOI22xp33_ASAP7_75t_R g12728 ( 
.A1(n_12637),
.A2(n_2218),
.B1(n_2216),
.B2(n_2217),
.Y(n_12728)
);

AND2x2_ASAP7_75t_L g12729 ( 
.A(n_12539),
.B(n_2217),
.Y(n_12729)
);

AND2x2_ASAP7_75t_L g12730 ( 
.A(n_12570),
.B(n_2219),
.Y(n_12730)
);

AOI22x1_ASAP7_75t_L g12731 ( 
.A1(n_12630),
.A2(n_2222),
.B1(n_2220),
.B2(n_2221),
.Y(n_12731)
);

AOI21xp5_ASAP7_75t_L g12732 ( 
.A1(n_12626),
.A2(n_2220),
.B(n_2221),
.Y(n_12732)
);

INVx2_ASAP7_75t_L g12733 ( 
.A(n_12553),
.Y(n_12733)
);

NAND2xp5_ASAP7_75t_L g12734 ( 
.A(n_12544),
.B(n_2222),
.Y(n_12734)
);

OR2x2_ASAP7_75t_L g12735 ( 
.A(n_12647),
.B(n_2223),
.Y(n_12735)
);

CKINVDCx20_ASAP7_75t_R g12736 ( 
.A(n_12639),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_12586),
.B(n_2223),
.Y(n_12737)
);

INVx2_ASAP7_75t_L g12738 ( 
.A(n_12602),
.Y(n_12738)
);

NAND2xp5_ASAP7_75t_L g12739 ( 
.A(n_12533),
.B(n_2225),
.Y(n_12739)
);

HB1xp67_ASAP7_75t_L g12740 ( 
.A(n_12546),
.Y(n_12740)
);

OR2x2_ASAP7_75t_L g12741 ( 
.A(n_12636),
.B(n_2225),
.Y(n_12741)
);

INVx1_ASAP7_75t_L g12742 ( 
.A(n_12561),
.Y(n_12742)
);

INVx2_ASAP7_75t_L g12743 ( 
.A(n_12603),
.Y(n_12743)
);

OR2x2_ASAP7_75t_L g12744 ( 
.A(n_12619),
.B(n_2226),
.Y(n_12744)
);

INVx1_ASAP7_75t_L g12745 ( 
.A(n_12613),
.Y(n_12745)
);

NAND2xp5_ASAP7_75t_L g12746 ( 
.A(n_12610),
.B(n_2226),
.Y(n_12746)
);

NAND2xp5_ASAP7_75t_SL g12747 ( 
.A(n_12582),
.B(n_2227),
.Y(n_12747)
);

NAND2xp5_ASAP7_75t_L g12748 ( 
.A(n_12623),
.B(n_2228),
.Y(n_12748)
);

INVx1_ASAP7_75t_L g12749 ( 
.A(n_12538),
.Y(n_12749)
);

NAND2xp5_ASAP7_75t_L g12750 ( 
.A(n_12635),
.B(n_2228),
.Y(n_12750)
);

AOI22xp33_ASAP7_75t_SL g12751 ( 
.A1(n_12617),
.A2(n_2231),
.B1(n_2229),
.B2(n_2230),
.Y(n_12751)
);

OR2x2_ASAP7_75t_L g12752 ( 
.A(n_12592),
.B(n_2231),
.Y(n_12752)
);

INVx2_ASAP7_75t_L g12753 ( 
.A(n_12604),
.Y(n_12753)
);

NAND2xp5_ASAP7_75t_SL g12754 ( 
.A(n_12618),
.B(n_2232),
.Y(n_12754)
);

OR2x2_ASAP7_75t_L g12755 ( 
.A(n_12593),
.B(n_2233),
.Y(n_12755)
);

AND2x2_ASAP7_75t_L g12756 ( 
.A(n_12581),
.B(n_2233),
.Y(n_12756)
);

NAND2xp5_ASAP7_75t_L g12757 ( 
.A(n_12567),
.B(n_12607),
.Y(n_12757)
);

NOR2x1_ASAP7_75t_L g12758 ( 
.A(n_12629),
.B(n_2234),
.Y(n_12758)
);

NAND2xp5_ASAP7_75t_L g12759 ( 
.A(n_12599),
.B(n_2234),
.Y(n_12759)
);

NOR2xp33_ASAP7_75t_L g12760 ( 
.A(n_12595),
.B(n_2236),
.Y(n_12760)
);

NOR2xp33_ASAP7_75t_L g12761 ( 
.A(n_12620),
.B(n_2236),
.Y(n_12761)
);

AOI221xp5_ASAP7_75t_L g12762 ( 
.A1(n_12551),
.A2(n_2240),
.B1(n_2237),
.B2(n_2238),
.C(n_2241),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_12624),
.B(n_2237),
.Y(n_12763)
);

INVx1_ASAP7_75t_L g12764 ( 
.A(n_12605),
.Y(n_12764)
);

INVx1_ASAP7_75t_L g12765 ( 
.A(n_12634),
.Y(n_12765)
);

INVx1_ASAP7_75t_L g12766 ( 
.A(n_12634),
.Y(n_12766)
);

INVx1_ASAP7_75t_L g12767 ( 
.A(n_12634),
.Y(n_12767)
);

AOI22xp33_ASAP7_75t_L g12768 ( 
.A1(n_12588),
.A2(n_2241),
.B1(n_2238),
.B2(n_2240),
.Y(n_12768)
);

INVx1_ASAP7_75t_L g12769 ( 
.A(n_12657),
.Y(n_12769)
);

OA22x2_ASAP7_75t_L g12770 ( 
.A1(n_12674),
.A2(n_2245),
.B1(n_2243),
.B2(n_2244),
.Y(n_12770)
);

AOI221xp5_ASAP7_75t_L g12771 ( 
.A1(n_12692),
.A2(n_2245),
.B1(n_2243),
.B2(n_2244),
.C(n_2246),
.Y(n_12771)
);

OAI322xp33_ASAP7_75t_L g12772 ( 
.A1(n_12739),
.A2(n_2270),
.A3(n_2254),
.B1(n_2278),
.B2(n_2286),
.C1(n_2262),
.C2(n_2246),
.Y(n_12772)
);

AOI22xp5_ASAP7_75t_L g12773 ( 
.A1(n_12664),
.A2(n_2249),
.B1(n_2247),
.B2(n_2248),
.Y(n_12773)
);

OAI322xp33_ASAP7_75t_L g12774 ( 
.A1(n_12765),
.A2(n_12766),
.A3(n_12767),
.B1(n_12663),
.B2(n_12720),
.C1(n_12749),
.C2(n_12699),
.Y(n_12774)
);

AOI22xp5_ASAP7_75t_L g12775 ( 
.A1(n_12736),
.A2(n_2249),
.B1(n_2247),
.B2(n_2248),
.Y(n_12775)
);

OAI22xp5_ASAP7_75t_L g12776 ( 
.A1(n_12662),
.A2(n_2252),
.B1(n_2250),
.B2(n_2251),
.Y(n_12776)
);

NAND4xp75_ASAP7_75t_L g12777 ( 
.A(n_12713),
.B(n_2253),
.C(n_2250),
.D(n_2251),
.Y(n_12777)
);

OAI22x1_ASAP7_75t_L g12778 ( 
.A1(n_12731),
.A2(n_2255),
.B1(n_2253),
.B2(n_2254),
.Y(n_12778)
);

INVx2_ASAP7_75t_L g12779 ( 
.A(n_12658),
.Y(n_12779)
);

AOI22xp33_ASAP7_75t_L g12780 ( 
.A1(n_12708),
.A2(n_2257),
.B1(n_2258),
.B2(n_2256),
.Y(n_12780)
);

INVx2_ASAP7_75t_SL g12781 ( 
.A(n_12726),
.Y(n_12781)
);

INVx2_ASAP7_75t_L g12782 ( 
.A(n_12666),
.Y(n_12782)
);

AOI22xp5_ASAP7_75t_L g12783 ( 
.A1(n_12745),
.A2(n_2257),
.B1(n_2255),
.B2(n_2256),
.Y(n_12783)
);

INVx1_ASAP7_75t_L g12784 ( 
.A(n_12702),
.Y(n_12784)
);

INVx2_ASAP7_75t_L g12785 ( 
.A(n_12666),
.Y(n_12785)
);

INVx1_ASAP7_75t_L g12786 ( 
.A(n_12667),
.Y(n_12786)
);

A2O1A1Ixp33_ASAP7_75t_L g12787 ( 
.A1(n_12665),
.A2(n_2260),
.B(n_2258),
.C(n_2259),
.Y(n_12787)
);

NAND4xp75_ASAP7_75t_L g12788 ( 
.A(n_12678),
.B(n_2263),
.C(n_2260),
.D(n_2261),
.Y(n_12788)
);

INVx2_ASAP7_75t_SL g12789 ( 
.A(n_12652),
.Y(n_12789)
);

INVx1_ASAP7_75t_L g12790 ( 
.A(n_12669),
.Y(n_12790)
);

AOI22xp5_ASAP7_75t_L g12791 ( 
.A1(n_12653),
.A2(n_2265),
.B1(n_2261),
.B2(n_2264),
.Y(n_12791)
);

AOI22xp5_ASAP7_75t_L g12792 ( 
.A1(n_12712),
.A2(n_2267),
.B1(n_2265),
.B2(n_2266),
.Y(n_12792)
);

INVx1_ASAP7_75t_L g12793 ( 
.A(n_12707),
.Y(n_12793)
);

OA22x2_ASAP7_75t_L g12794 ( 
.A1(n_12681),
.A2(n_2268),
.B1(n_2266),
.B2(n_2267),
.Y(n_12794)
);

AOI221xp5_ASAP7_75t_L g12795 ( 
.A1(n_12697),
.A2(n_2272),
.B1(n_2269),
.B2(n_2271),
.C(n_2273),
.Y(n_12795)
);

AO22x2_ASAP7_75t_L g12796 ( 
.A1(n_12686),
.A2(n_2273),
.B1(n_2271),
.B2(n_2272),
.Y(n_12796)
);

INVx1_ASAP7_75t_L g12797 ( 
.A(n_12711),
.Y(n_12797)
);

NAND4xp75_ASAP7_75t_SL g12798 ( 
.A(n_12670),
.B(n_2276),
.C(n_2274),
.D(n_2275),
.Y(n_12798)
);

OAI322xp33_ASAP7_75t_L g12799 ( 
.A1(n_12710),
.A2(n_2302),
.A3(n_2284),
.B1(n_2310),
.B2(n_2319),
.C1(n_2293),
.C2(n_2276),
.Y(n_12799)
);

INVx2_ASAP7_75t_L g12800 ( 
.A(n_12675),
.Y(n_12800)
);

AOI22xp5_ASAP7_75t_L g12801 ( 
.A1(n_12708),
.A2(n_2279),
.B1(n_2277),
.B2(n_2278),
.Y(n_12801)
);

INVx1_ASAP7_75t_L g12802 ( 
.A(n_12729),
.Y(n_12802)
);

NOR4xp25_ASAP7_75t_L g12803 ( 
.A(n_12654),
.B(n_2280),
.C(n_2277),
.D(n_2279),
.Y(n_12803)
);

AOI22xp5_ASAP7_75t_L g12804 ( 
.A1(n_12671),
.A2(n_2283),
.B1(n_2281),
.B2(n_2282),
.Y(n_12804)
);

INVx2_ASAP7_75t_L g12805 ( 
.A(n_12763),
.Y(n_12805)
);

INVx1_ASAP7_75t_L g12806 ( 
.A(n_12756),
.Y(n_12806)
);

AND4x1_ASAP7_75t_L g12807 ( 
.A(n_12722),
.B(n_2283),
.C(n_2281),
.D(n_2282),
.Y(n_12807)
);

AOI22xp5_ASAP7_75t_L g12808 ( 
.A1(n_12718),
.A2(n_2288),
.B1(n_2285),
.B2(n_2287),
.Y(n_12808)
);

HB1xp67_ASAP7_75t_L g12809 ( 
.A(n_12696),
.Y(n_12809)
);

INVx1_ASAP7_75t_L g12810 ( 
.A(n_12672),
.Y(n_12810)
);

AOI221xp5_ASAP7_75t_L g12811 ( 
.A1(n_12688),
.A2(n_2290),
.B1(n_2288),
.B2(n_2289),
.C(n_2291),
.Y(n_12811)
);

OA22x2_ASAP7_75t_L g12812 ( 
.A1(n_12687),
.A2(n_2292),
.B1(n_2289),
.B2(n_2290),
.Y(n_12812)
);

INVx1_ASAP7_75t_L g12813 ( 
.A(n_12655),
.Y(n_12813)
);

INVx1_ASAP7_75t_L g12814 ( 
.A(n_12660),
.Y(n_12814)
);

INVx1_ASAP7_75t_L g12815 ( 
.A(n_12691),
.Y(n_12815)
);

HB1xp67_ASAP7_75t_L g12816 ( 
.A(n_12659),
.Y(n_12816)
);

AOI31xp33_ASAP7_75t_L g12817 ( 
.A1(n_12755),
.A2(n_2294),
.A3(n_2292),
.B(n_2293),
.Y(n_12817)
);

AOI221xp5_ASAP7_75t_L g12818 ( 
.A1(n_12742),
.A2(n_2296),
.B1(n_2294),
.B2(n_2295),
.C(n_2297),
.Y(n_12818)
);

INVx1_ASAP7_75t_L g12819 ( 
.A(n_12679),
.Y(n_12819)
);

INVx1_ASAP7_75t_L g12820 ( 
.A(n_12650),
.Y(n_12820)
);

INVx1_ASAP7_75t_SL g12821 ( 
.A(n_12685),
.Y(n_12821)
);

INVx1_ASAP7_75t_L g12822 ( 
.A(n_12680),
.Y(n_12822)
);

INVx2_ASAP7_75t_L g12823 ( 
.A(n_12735),
.Y(n_12823)
);

INVx1_ASAP7_75t_L g12824 ( 
.A(n_12683),
.Y(n_12824)
);

INVx1_ASAP7_75t_L g12825 ( 
.A(n_12656),
.Y(n_12825)
);

INVx1_ASAP7_75t_SL g12826 ( 
.A(n_12661),
.Y(n_12826)
);

AOI22xp33_ASAP7_75t_SL g12827 ( 
.A1(n_12740),
.A2(n_2298),
.B1(n_2295),
.B2(n_2296),
.Y(n_12827)
);

INVx1_ASAP7_75t_L g12828 ( 
.A(n_12651),
.Y(n_12828)
);

OA22x2_ASAP7_75t_L g12829 ( 
.A1(n_12690),
.A2(n_2302),
.B1(n_2299),
.B2(n_2300),
.Y(n_12829)
);

INVx1_ASAP7_75t_SL g12830 ( 
.A(n_12716),
.Y(n_12830)
);

AOI22xp5_ASAP7_75t_L g12831 ( 
.A1(n_12714),
.A2(n_2304),
.B1(n_2300),
.B2(n_2303),
.Y(n_12831)
);

HB1xp67_ASAP7_75t_L g12832 ( 
.A(n_12727),
.Y(n_12832)
);

AO22x1_ASAP7_75t_L g12833 ( 
.A1(n_12758),
.A2(n_2305),
.B1(n_2303),
.B2(n_2304),
.Y(n_12833)
);

OAI322xp33_ASAP7_75t_L g12834 ( 
.A1(n_12754),
.A2(n_2331),
.A3(n_2314),
.B1(n_2339),
.B2(n_2347),
.C1(n_2323),
.C2(n_2306),
.Y(n_12834)
);

AOI22xp5_ASAP7_75t_L g12835 ( 
.A1(n_12717),
.A2(n_12719),
.B1(n_12723),
.B2(n_12677),
.Y(n_12835)
);

INVx3_ASAP7_75t_L g12836 ( 
.A(n_12733),
.Y(n_12836)
);

INVx1_ASAP7_75t_L g12837 ( 
.A(n_12724),
.Y(n_12837)
);

INVx1_ASAP7_75t_L g12838 ( 
.A(n_12694),
.Y(n_12838)
);

OAI322xp33_ASAP7_75t_L g12839 ( 
.A1(n_12764),
.A2(n_2332),
.A3(n_2314),
.B1(n_2340),
.B2(n_2348),
.C1(n_2323),
.C2(n_2306),
.Y(n_12839)
);

OAI22xp5_ASAP7_75t_L g12840 ( 
.A1(n_12768),
.A2(n_2309),
.B1(n_2307),
.B2(n_2308),
.Y(n_12840)
);

AOI22xp5_ASAP7_75t_L g12841 ( 
.A1(n_12738),
.A2(n_2310),
.B1(n_2307),
.B2(n_2308),
.Y(n_12841)
);

AOI22xp5_ASAP7_75t_L g12842 ( 
.A1(n_12743),
.A2(n_2313),
.B1(n_2311),
.B2(n_2312),
.Y(n_12842)
);

INVx1_ASAP7_75t_L g12843 ( 
.A(n_12761),
.Y(n_12843)
);

AOI22xp5_ASAP7_75t_L g12844 ( 
.A1(n_12753),
.A2(n_2313),
.B1(n_2311),
.B2(n_2312),
.Y(n_12844)
);

INVx2_ASAP7_75t_L g12845 ( 
.A(n_12741),
.Y(n_12845)
);

OA22x2_ASAP7_75t_L g12846 ( 
.A1(n_12746),
.A2(n_2318),
.B1(n_2316),
.B2(n_2317),
.Y(n_12846)
);

AOI22xp5_ASAP7_75t_L g12847 ( 
.A1(n_12704),
.A2(n_2319),
.B1(n_2317),
.B2(n_2318),
.Y(n_12847)
);

OAI22xp5_ASAP7_75t_L g12848 ( 
.A1(n_12706),
.A2(n_2322),
.B1(n_2320),
.B2(n_2321),
.Y(n_12848)
);

AOI22xp5_ASAP7_75t_L g12849 ( 
.A1(n_12730),
.A2(n_2324),
.B1(n_2320),
.B2(n_2321),
.Y(n_12849)
);

AND4x1_ASAP7_75t_L g12850 ( 
.A(n_12673),
.B(n_2326),
.C(n_2324),
.D(n_2325),
.Y(n_12850)
);

NAND4xp25_ASAP7_75t_L g12851 ( 
.A(n_12757),
.B(n_2328),
.C(n_2326),
.D(n_2327),
.Y(n_12851)
);

INVx1_ASAP7_75t_L g12852 ( 
.A(n_12760),
.Y(n_12852)
);

AOI22xp5_ASAP7_75t_L g12853 ( 
.A1(n_12676),
.A2(n_2330),
.B1(n_2327),
.B2(n_2329),
.Y(n_12853)
);

AOI22xp5_ASAP7_75t_L g12854 ( 
.A1(n_12725),
.A2(n_2335),
.B1(n_2333),
.B2(n_2334),
.Y(n_12854)
);

AOI22x1_ASAP7_75t_L g12855 ( 
.A1(n_12732),
.A2(n_2336),
.B1(n_2333),
.B2(n_2334),
.Y(n_12855)
);

INVx2_ASAP7_75t_SL g12856 ( 
.A(n_12689),
.Y(n_12856)
);

OA22x2_ASAP7_75t_L g12857 ( 
.A1(n_12750),
.A2(n_2338),
.B1(n_2336),
.B2(n_2337),
.Y(n_12857)
);

INVx1_ASAP7_75t_L g12858 ( 
.A(n_12759),
.Y(n_12858)
);

NOR3xp33_ASAP7_75t_L g12859 ( 
.A(n_12774),
.B(n_12684),
.C(n_12682),
.Y(n_12859)
);

INVx1_ASAP7_75t_L g12860 ( 
.A(n_12794),
.Y(n_12860)
);

AOI21xp5_ASAP7_75t_L g12861 ( 
.A1(n_12809),
.A2(n_12747),
.B(n_12700),
.Y(n_12861)
);

NAND3xp33_ASAP7_75t_L g12862 ( 
.A(n_12811),
.B(n_12728),
.C(n_12715),
.Y(n_12862)
);

OAI211xp5_ASAP7_75t_SL g12863 ( 
.A1(n_12790),
.A2(n_12701),
.B(n_12705),
.C(n_12693),
.Y(n_12863)
);

NAND2xp5_ASAP7_75t_L g12864 ( 
.A(n_12833),
.B(n_12751),
.Y(n_12864)
);

NOR3xp33_ASAP7_75t_L g12865 ( 
.A(n_12813),
.B(n_12698),
.C(n_12734),
.Y(n_12865)
);

AOI21xp5_ASAP7_75t_SL g12866 ( 
.A1(n_12778),
.A2(n_12787),
.B(n_12817),
.Y(n_12866)
);

NOR2x1_ASAP7_75t_L g12867 ( 
.A(n_12777),
.B(n_12721),
.Y(n_12867)
);

NOR2xp33_ASAP7_75t_L g12868 ( 
.A(n_12834),
.B(n_12709),
.Y(n_12868)
);

INVx1_ASAP7_75t_L g12869 ( 
.A(n_12846),
.Y(n_12869)
);

AOI211x1_ASAP7_75t_L g12870 ( 
.A1(n_12769),
.A2(n_12737),
.B(n_12695),
.C(n_12748),
.Y(n_12870)
);

AOI22xp5_ASAP7_75t_L g12871 ( 
.A1(n_12856),
.A2(n_12744),
.B1(n_12752),
.B2(n_12762),
.Y(n_12871)
);

NOR3xp33_ASAP7_75t_L g12872 ( 
.A(n_12836),
.B(n_12668),
.C(n_12703),
.Y(n_12872)
);

NAND2xp5_ASAP7_75t_SL g12873 ( 
.A(n_12803),
.B(n_2337),
.Y(n_12873)
);

NAND2xp5_ASAP7_75t_L g12874 ( 
.A(n_12827),
.B(n_2338),
.Y(n_12874)
);

AOI21xp5_ASAP7_75t_L g12875 ( 
.A1(n_12779),
.A2(n_12781),
.B(n_12782),
.Y(n_12875)
);

AO22x2_ASAP7_75t_L g12876 ( 
.A1(n_12786),
.A2(n_12785),
.B1(n_12784),
.B2(n_12789),
.Y(n_12876)
);

AO21x1_ASAP7_75t_L g12877 ( 
.A1(n_12776),
.A2(n_2339),
.B(n_2340),
.Y(n_12877)
);

NOR3x1_ASAP7_75t_L g12878 ( 
.A(n_12840),
.B(n_12788),
.C(n_12851),
.Y(n_12878)
);

AOI21xp5_ASAP7_75t_L g12879 ( 
.A1(n_12832),
.A2(n_2349),
.B(n_2341),
.Y(n_12879)
);

AOI211x1_ASAP7_75t_L g12880 ( 
.A1(n_12807),
.A2(n_2344),
.B(n_2342),
.C(n_2343),
.Y(n_12880)
);

INVx1_ASAP7_75t_L g12881 ( 
.A(n_12812),
.Y(n_12881)
);

OR2x2_ASAP7_75t_L g12882 ( 
.A(n_12816),
.B(n_2342),
.Y(n_12882)
);

OA22x2_ASAP7_75t_L g12883 ( 
.A1(n_12791),
.A2(n_2345),
.B1(n_2343),
.B2(n_2344),
.Y(n_12883)
);

OAI22xp5_ASAP7_75t_L g12884 ( 
.A1(n_12831),
.A2(n_2347),
.B1(n_2345),
.B2(n_2346),
.Y(n_12884)
);

OAI21xp33_ASAP7_75t_SL g12885 ( 
.A1(n_12798),
.A2(n_2356),
.B(n_2346),
.Y(n_12885)
);

NOR4xp25_ASAP7_75t_L g12886 ( 
.A(n_12830),
.B(n_2350),
.C(n_2348),
.D(n_2349),
.Y(n_12886)
);

NOR4xp25_ASAP7_75t_L g12887 ( 
.A(n_12821),
.B(n_2353),
.C(n_2350),
.D(n_2351),
.Y(n_12887)
);

AOI22x1_ASAP7_75t_L g12888 ( 
.A1(n_12805),
.A2(n_2354),
.B1(n_2351),
.B2(n_2353),
.Y(n_12888)
);

AND4x1_ASAP7_75t_L g12889 ( 
.A(n_12835),
.B(n_2356),
.C(n_2354),
.D(n_2355),
.Y(n_12889)
);

AO22x2_ASAP7_75t_L g12890 ( 
.A1(n_12793),
.A2(n_2360),
.B1(n_2361),
.B2(n_2358),
.Y(n_12890)
);

INVx1_ASAP7_75t_L g12891 ( 
.A(n_12857),
.Y(n_12891)
);

AOI21xp5_ASAP7_75t_L g12892 ( 
.A1(n_12848),
.A2(n_2367),
.B(n_2357),
.Y(n_12892)
);

NAND2xp5_ASAP7_75t_L g12893 ( 
.A(n_12850),
.B(n_2358),
.Y(n_12893)
);

AOI21xp5_ASAP7_75t_L g12894 ( 
.A1(n_12800),
.A2(n_2369),
.B(n_2360),
.Y(n_12894)
);

INVxp67_ASAP7_75t_SL g12895 ( 
.A(n_12796),
.Y(n_12895)
);

OAI21xp33_ASAP7_75t_L g12896 ( 
.A1(n_12797),
.A2(n_2361),
.B(n_2362),
.Y(n_12896)
);

NAND3xp33_ASAP7_75t_L g12897 ( 
.A(n_12771),
.B(n_2362),
.C(n_2363),
.Y(n_12897)
);

NOR4xp25_ASAP7_75t_L g12898 ( 
.A(n_12826),
.B(n_2365),
.C(n_2363),
.D(n_2364),
.Y(n_12898)
);

AOI22xp5_ASAP7_75t_L g12899 ( 
.A1(n_12802),
.A2(n_2376),
.B1(n_2384),
.B2(n_2365),
.Y(n_12899)
);

AOI22xp5_ASAP7_75t_L g12900 ( 
.A1(n_12806),
.A2(n_2377),
.B1(n_2386),
.B2(n_2367),
.Y(n_12900)
);

NOR2xp33_ASAP7_75t_L g12901 ( 
.A(n_12772),
.B(n_12770),
.Y(n_12901)
);

AOI21xp5_ASAP7_75t_L g12902 ( 
.A1(n_12829),
.A2(n_12795),
.B(n_12820),
.Y(n_12902)
);

AOI22xp5_ASAP7_75t_L g12903 ( 
.A1(n_12828),
.A2(n_12810),
.B1(n_12852),
.B2(n_12843),
.Y(n_12903)
);

NOR3xp33_ASAP7_75t_L g12904 ( 
.A(n_12837),
.B(n_2371),
.C(n_2370),
.Y(n_12904)
);

AOI21xp5_ASAP7_75t_L g12905 ( 
.A1(n_12823),
.A2(n_2378),
.B(n_2368),
.Y(n_12905)
);

AOI211xp5_ASAP7_75t_L g12906 ( 
.A1(n_12799),
.A2(n_2371),
.B(n_2368),
.C(n_2370),
.Y(n_12906)
);

INVx1_ASAP7_75t_L g12907 ( 
.A(n_12855),
.Y(n_12907)
);

OAI21xp5_ASAP7_75t_L g12908 ( 
.A1(n_12819),
.A2(n_2382),
.B(n_2373),
.Y(n_12908)
);

XNOR2xp5_ASAP7_75t_L g12909 ( 
.A(n_12808),
.B(n_2373),
.Y(n_12909)
);

NOR3x1_ASAP7_75t_L g12910 ( 
.A(n_12814),
.B(n_12838),
.C(n_12825),
.Y(n_12910)
);

NAND2xp5_ASAP7_75t_L g12911 ( 
.A(n_12775),
.B(n_2374),
.Y(n_12911)
);

OAI21xp5_ASAP7_75t_SL g12912 ( 
.A1(n_12822),
.A2(n_2376),
.B(n_2375),
.Y(n_12912)
);

INVx1_ASAP7_75t_L g12913 ( 
.A(n_12796),
.Y(n_12913)
);

NAND4xp75_ASAP7_75t_SL g12914 ( 
.A(n_12845),
.B(n_2377),
.C(n_2374),
.D(n_2375),
.Y(n_12914)
);

AO22x2_ASAP7_75t_L g12915 ( 
.A1(n_12815),
.A2(n_2381),
.B1(n_2382),
.B2(n_2380),
.Y(n_12915)
);

NOR3xp33_ASAP7_75t_L g12916 ( 
.A(n_12824),
.B(n_12858),
.C(n_12818),
.Y(n_12916)
);

NAND2xp5_ASAP7_75t_L g12917 ( 
.A(n_12783),
.B(n_2379),
.Y(n_12917)
);

OAI22xp5_ASAP7_75t_SL g12918 ( 
.A1(n_12780),
.A2(n_2383),
.B1(n_2379),
.B2(n_2380),
.Y(n_12918)
);

XOR2xp5_ASAP7_75t_L g12919 ( 
.A(n_12849),
.B(n_2385),
.Y(n_12919)
);

AOI22x1_ASAP7_75t_SL g12920 ( 
.A1(n_12839),
.A2(n_2896),
.B1(n_2897),
.B2(n_2895),
.Y(n_12920)
);

INVx1_ASAP7_75t_L g12921 ( 
.A(n_12804),
.Y(n_12921)
);

NOR3xp33_ASAP7_75t_L g12922 ( 
.A(n_12773),
.B(n_2388),
.C(n_2387),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12847),
.Y(n_12923)
);

NOR3x1_ASAP7_75t_L g12924 ( 
.A(n_12841),
.B(n_2386),
.C(n_2387),
.Y(n_12924)
);

NOR2xp33_ASAP7_75t_L g12925 ( 
.A(n_12842),
.B(n_2389),
.Y(n_12925)
);

AOI21xp5_ASAP7_75t_L g12926 ( 
.A1(n_12844),
.A2(n_2399),
.B(n_2390),
.Y(n_12926)
);

INVx2_ASAP7_75t_L g12927 ( 
.A(n_12890),
.Y(n_12927)
);

NOR2x1_ASAP7_75t_L g12928 ( 
.A(n_12913),
.B(n_12792),
.Y(n_12928)
);

NAND2xp5_ASAP7_75t_L g12929 ( 
.A(n_12895),
.B(n_12854),
.Y(n_12929)
);

AND5x1_ASAP7_75t_L g12930 ( 
.A(n_12901),
.B(n_12853),
.C(n_12801),
.D(n_2393),
.E(n_2391),
.Y(n_12930)
);

NAND4xp75_ASAP7_75t_L g12931 ( 
.A(n_12910),
.B(n_2917),
.C(n_2915),
.D(n_2393),
.Y(n_12931)
);

INVx1_ASAP7_75t_L g12932 ( 
.A(n_12882),
.Y(n_12932)
);

OAI21xp5_ASAP7_75t_L g12933 ( 
.A1(n_12875),
.A2(n_2391),
.B(n_2392),
.Y(n_12933)
);

AND2x2_ASAP7_75t_L g12934 ( 
.A(n_12876),
.B(n_2394),
.Y(n_12934)
);

NAND3xp33_ASAP7_75t_L g12935 ( 
.A(n_12859),
.B(n_2392),
.C(n_2396),
.Y(n_12935)
);

AND2x2_ASAP7_75t_L g12936 ( 
.A(n_12876),
.B(n_2397),
.Y(n_12936)
);

NAND3xp33_ASAP7_75t_L g12937 ( 
.A(n_12872),
.B(n_2396),
.C(n_2397),
.Y(n_12937)
);

INVx2_ASAP7_75t_L g12938 ( 
.A(n_12890),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12893),
.Y(n_12939)
);

NAND2xp5_ASAP7_75t_L g12940 ( 
.A(n_12880),
.B(n_2398),
.Y(n_12940)
);

INVx1_ASAP7_75t_L g12941 ( 
.A(n_12883),
.Y(n_12941)
);

NAND2xp5_ASAP7_75t_L g12942 ( 
.A(n_12889),
.B(n_2399),
.Y(n_12942)
);

INVx1_ASAP7_75t_L g12943 ( 
.A(n_12920),
.Y(n_12943)
);

INVx1_ASAP7_75t_L g12944 ( 
.A(n_12877),
.Y(n_12944)
);

NOR2x1_ASAP7_75t_L g12945 ( 
.A(n_12914),
.B(n_2402),
.Y(n_12945)
);

NOR3xp33_ASAP7_75t_L g12946 ( 
.A(n_12863),
.B(n_2401),
.C(n_2403),
.Y(n_12946)
);

NOR2x1_ASAP7_75t_L g12947 ( 
.A(n_12912),
.B(n_2403),
.Y(n_12947)
);

NAND2xp5_ASAP7_75t_L g12948 ( 
.A(n_12879),
.B(n_2401),
.Y(n_12948)
);

NAND4xp25_ASAP7_75t_L g12949 ( 
.A(n_12878),
.B(n_2406),
.C(n_2404),
.D(n_2405),
.Y(n_12949)
);

NOR3xp33_ASAP7_75t_L g12950 ( 
.A(n_12865),
.B(n_2406),
.C(n_2408),
.Y(n_12950)
);

NOR2xp33_ASAP7_75t_SL g12951 ( 
.A(n_12896),
.B(n_12881),
.Y(n_12951)
);

NAND4xp25_ASAP7_75t_L g12952 ( 
.A(n_12906),
.B(n_2410),
.C(n_2408),
.D(n_2409),
.Y(n_12952)
);

NOR2x1_ASAP7_75t_L g12953 ( 
.A(n_12869),
.B(n_2411),
.Y(n_12953)
);

INVx1_ASAP7_75t_L g12954 ( 
.A(n_12874),
.Y(n_12954)
);

AOI22xp5_ASAP7_75t_L g12955 ( 
.A1(n_12860),
.A2(n_2413),
.B1(n_2410),
.B2(n_2411),
.Y(n_12955)
);

INVxp67_ASAP7_75t_L g12956 ( 
.A(n_12888),
.Y(n_12956)
);

NOR2x1_ASAP7_75t_L g12957 ( 
.A(n_12891),
.B(n_2414),
.Y(n_12957)
);

NOR2x1_ASAP7_75t_L g12958 ( 
.A(n_12908),
.B(n_2414),
.Y(n_12958)
);

NOR3x1_ASAP7_75t_L g12959 ( 
.A(n_12897),
.B(n_2413),
.C(n_2415),
.Y(n_12959)
);

NAND2xp5_ASAP7_75t_L g12960 ( 
.A(n_12904),
.B(n_2416),
.Y(n_12960)
);

INVx1_ASAP7_75t_L g12961 ( 
.A(n_12864),
.Y(n_12961)
);

NOR3xp33_ASAP7_75t_L g12962 ( 
.A(n_12861),
.B(n_2417),
.C(n_2418),
.Y(n_12962)
);

INVx1_ASAP7_75t_L g12963 ( 
.A(n_12919),
.Y(n_12963)
);

AOI22xp5_ASAP7_75t_L g12964 ( 
.A1(n_12885),
.A2(n_2420),
.B1(n_2418),
.B2(n_2419),
.Y(n_12964)
);

NAND5xp2_ASAP7_75t_L g12965 ( 
.A(n_12903),
.B(n_2421),
.C(n_2423),
.D(n_2420),
.E(n_2422),
.Y(n_12965)
);

NOR3xp33_ASAP7_75t_L g12966 ( 
.A(n_12916),
.B(n_2419),
.C(n_2421),
.Y(n_12966)
);

AOI21xp5_ASAP7_75t_L g12967 ( 
.A1(n_12866),
.A2(n_2422),
.B(n_2423),
.Y(n_12967)
);

NAND2xp5_ASAP7_75t_L g12968 ( 
.A(n_12894),
.B(n_2424),
.Y(n_12968)
);

NOR3x1_ASAP7_75t_L g12969 ( 
.A(n_12862),
.B(n_2424),
.C(n_2425),
.Y(n_12969)
);

NAND2xp5_ASAP7_75t_SL g12970 ( 
.A(n_12887),
.B(n_2425),
.Y(n_12970)
);

NAND3xp33_ASAP7_75t_L g12971 ( 
.A(n_12922),
.B(n_2426),
.C(n_2427),
.Y(n_12971)
);

NAND5xp2_ASAP7_75t_L g12972 ( 
.A(n_12868),
.B(n_2430),
.C(n_2432),
.D(n_2428),
.E(n_2431),
.Y(n_12972)
);

NAND3xp33_ASAP7_75t_L g12973 ( 
.A(n_12870),
.B(n_2426),
.C(n_2428),
.Y(n_12973)
);

NAND3xp33_ASAP7_75t_L g12974 ( 
.A(n_12946),
.B(n_12871),
.C(n_12907),
.Y(n_12974)
);

NAND4xp25_ASAP7_75t_L g12975 ( 
.A(n_12951),
.B(n_12964),
.C(n_12969),
.D(n_12902),
.Y(n_12975)
);

AOI21xp5_ASAP7_75t_L g12976 ( 
.A1(n_12970),
.A2(n_12873),
.B(n_12911),
.Y(n_12976)
);

AND4x2_ASAP7_75t_L g12977 ( 
.A(n_12928),
.B(n_12867),
.C(n_12892),
.D(n_12926),
.Y(n_12977)
);

INVx1_ASAP7_75t_SL g12978 ( 
.A(n_12934),
.Y(n_12978)
);

NAND3xp33_ASAP7_75t_L g12979 ( 
.A(n_12966),
.B(n_12962),
.C(n_12935),
.Y(n_12979)
);

NAND2xp5_ASAP7_75t_L g12980 ( 
.A(n_12936),
.B(n_12905),
.Y(n_12980)
);

NOR3xp33_ASAP7_75t_L g12981 ( 
.A(n_12929),
.B(n_12961),
.C(n_12943),
.Y(n_12981)
);

NOR3x1_ASAP7_75t_L g12982 ( 
.A(n_12931),
.B(n_12917),
.C(n_12921),
.Y(n_12982)
);

NOR3xp33_ASAP7_75t_L g12983 ( 
.A(n_12932),
.B(n_12973),
.C(n_12944),
.Y(n_12983)
);

INVx2_ASAP7_75t_L g12984 ( 
.A(n_12927),
.Y(n_12984)
);

AOI211xp5_ASAP7_75t_SL g12985 ( 
.A1(n_12956),
.A2(n_12923),
.B(n_12925),
.C(n_12884),
.Y(n_12985)
);

NOR4xp25_ASAP7_75t_L g12986 ( 
.A(n_12941),
.B(n_12909),
.C(n_12924),
.D(n_12886),
.Y(n_12986)
);

NAND3xp33_ASAP7_75t_L g12987 ( 
.A(n_12937),
.B(n_12898),
.C(n_12899),
.Y(n_12987)
);

NOR3xp33_ASAP7_75t_SL g12988 ( 
.A(n_12952),
.B(n_12918),
.C(n_12900),
.Y(n_12988)
);

NAND3xp33_ASAP7_75t_SL g12989 ( 
.A(n_12967),
.B(n_12915),
.C(n_2431),
.Y(n_12989)
);

NAND4xp75_ASAP7_75t_SL g12990 ( 
.A(n_12930),
.B(n_12915),
.C(n_2435),
.D(n_2432),
.Y(n_12990)
);

NOR3xp33_ASAP7_75t_L g12991 ( 
.A(n_12963),
.B(n_2892),
.C(n_2891),
.Y(n_12991)
);

NOR2xp67_ASAP7_75t_L g12992 ( 
.A(n_12965),
.B(n_2435),
.Y(n_12992)
);

INVx1_ASAP7_75t_L g12993 ( 
.A(n_12953),
.Y(n_12993)
);

NOR2xp33_ASAP7_75t_L g12994 ( 
.A(n_12972),
.B(n_2433),
.Y(n_12994)
);

NAND2xp5_ASAP7_75t_L g12995 ( 
.A(n_12957),
.B(n_2436),
.Y(n_12995)
);

NAND3xp33_ASAP7_75t_L g12996 ( 
.A(n_12933),
.B(n_2436),
.C(n_2437),
.Y(n_12996)
);

NAND4xp75_ASAP7_75t_L g12997 ( 
.A(n_12959),
.B(n_2439),
.C(n_2437),
.D(n_2438),
.Y(n_12997)
);

INVx3_ASAP7_75t_L g12998 ( 
.A(n_12938),
.Y(n_12998)
);

OR2x2_ASAP7_75t_L g12999 ( 
.A(n_12942),
.B(n_2438),
.Y(n_12999)
);

NOR3xp33_ASAP7_75t_SL g13000 ( 
.A(n_12940),
.B(n_2439),
.C(n_2440),
.Y(n_13000)
);

INVx1_ASAP7_75t_L g13001 ( 
.A(n_12945),
.Y(n_13001)
);

NOR3xp33_ASAP7_75t_L g13002 ( 
.A(n_12939),
.B(n_2911),
.C(n_2899),
.Y(n_13002)
);

AND2x2_ASAP7_75t_L g13003 ( 
.A(n_12947),
.B(n_2441),
.Y(n_13003)
);

NOR2x1_ASAP7_75t_L g13004 ( 
.A(n_12949),
.B(n_2443),
.Y(n_13004)
);

NAND4xp25_ASAP7_75t_L g13005 ( 
.A(n_12971),
.B(n_2445),
.C(n_2443),
.D(n_2444),
.Y(n_13005)
);

NOR3xp33_ASAP7_75t_L g13006 ( 
.A(n_12954),
.B(n_2444),
.C(n_2445),
.Y(n_13006)
);

NOR3xp33_ASAP7_75t_L g13007 ( 
.A(n_12960),
.B(n_2887),
.C(n_2886),
.Y(n_13007)
);

NOR2xp67_ASAP7_75t_L g13008 ( 
.A(n_12955),
.B(n_12948),
.Y(n_13008)
);

NAND2xp5_ASAP7_75t_L g13009 ( 
.A(n_12950),
.B(n_2446),
.Y(n_13009)
);

NOR3xp33_ASAP7_75t_L g13010 ( 
.A(n_12968),
.B(n_2887),
.C(n_2886),
.Y(n_13010)
);

NAND3xp33_ASAP7_75t_L g13011 ( 
.A(n_12958),
.B(n_2446),
.C(n_2447),
.Y(n_13011)
);

NOR3xp33_ASAP7_75t_L g13012 ( 
.A(n_12929),
.B(n_2890),
.C(n_2889),
.Y(n_13012)
);

NAND2xp5_ASAP7_75t_L g13013 ( 
.A(n_12934),
.B(n_2447),
.Y(n_13013)
);

NOR3xp33_ASAP7_75t_L g13014 ( 
.A(n_12929),
.B(n_2892),
.C(n_2890),
.Y(n_13014)
);

INVx2_ASAP7_75t_L g13015 ( 
.A(n_12934),
.Y(n_13015)
);

NOR2xp67_ASAP7_75t_SL g13016 ( 
.A(n_12944),
.B(n_2448),
.Y(n_13016)
);

NOR3x1_ASAP7_75t_L g13017 ( 
.A(n_12931),
.B(n_2448),
.C(n_2449),
.Y(n_13017)
);

AOI211x1_ASAP7_75t_L g13018 ( 
.A1(n_12935),
.A2(n_2452),
.B(n_2450),
.C(n_2451),
.Y(n_13018)
);

INVx2_ASAP7_75t_L g13019 ( 
.A(n_12934),
.Y(n_13019)
);

NAND3xp33_ASAP7_75t_L g13020 ( 
.A(n_12946),
.B(n_2450),
.C(n_2451),
.Y(n_13020)
);

NAND2xp5_ASAP7_75t_L g13021 ( 
.A(n_12934),
.B(n_2452),
.Y(n_13021)
);

NOR2xp33_ASAP7_75t_L g13022 ( 
.A(n_12972),
.B(n_2453),
.Y(n_13022)
);

INVx1_ASAP7_75t_L g13023 ( 
.A(n_13013),
.Y(n_13023)
);

OAI22xp5_ASAP7_75t_L g13024 ( 
.A1(n_13001),
.A2(n_12984),
.B1(n_12974),
.B2(n_13020),
.Y(n_13024)
);

AOI221xp5_ASAP7_75t_L g13025 ( 
.A1(n_12986),
.A2(n_2455),
.B1(n_2453),
.B2(n_2454),
.C(n_2456),
.Y(n_13025)
);

NOR3xp33_ASAP7_75t_L g13026 ( 
.A(n_12975),
.B(n_2454),
.C(n_2455),
.Y(n_13026)
);

AND2x2_ASAP7_75t_L g13027 ( 
.A(n_13000),
.B(n_12994),
.Y(n_13027)
);

NAND2xp5_ASAP7_75t_L g13028 ( 
.A(n_13016),
.B(n_2457),
.Y(n_13028)
);

INVx1_ASAP7_75t_SL g13029 ( 
.A(n_12990),
.Y(n_13029)
);

AOI221xp5_ASAP7_75t_L g13030 ( 
.A1(n_12981),
.A2(n_2460),
.B1(n_2457),
.B2(n_2459),
.C(n_2461),
.Y(n_13030)
);

AOI222xp33_ASAP7_75t_L g13031 ( 
.A1(n_12989),
.A2(n_2461),
.B1(n_2463),
.B2(n_2459),
.C1(n_2460),
.C2(n_2462),
.Y(n_13031)
);

OAI221xp5_ASAP7_75t_SL g13032 ( 
.A1(n_12978),
.A2(n_2889),
.B1(n_2893),
.B2(n_2888),
.C(n_2885),
.Y(n_13032)
);

AOI22xp5_ASAP7_75t_L g13033 ( 
.A1(n_13022),
.A2(n_12992),
.B1(n_12983),
.B2(n_13010),
.Y(n_13033)
);

INVx1_ASAP7_75t_L g13034 ( 
.A(n_13021),
.Y(n_13034)
);

AOI22xp33_ASAP7_75t_L g13035 ( 
.A1(n_12998),
.A2(n_2465),
.B1(n_2462),
.B2(n_2464),
.Y(n_13035)
);

NAND2xp5_ASAP7_75t_L g13036 ( 
.A(n_13002),
.B(n_2465),
.Y(n_13036)
);

NAND3x1_ASAP7_75t_SL g13037 ( 
.A(n_13004),
.B(n_2466),
.C(n_2467),
.Y(n_13037)
);

AOI222xp33_ASAP7_75t_L g13038 ( 
.A1(n_13003),
.A2(n_2468),
.B1(n_2470),
.B2(n_2466),
.C1(n_2467),
.C2(n_2469),
.Y(n_13038)
);

O2A1O1Ixp33_ASAP7_75t_L g13039 ( 
.A1(n_12995),
.A2(n_12993),
.B(n_12998),
.C(n_13009),
.Y(n_13039)
);

INVx1_ASAP7_75t_SL g13040 ( 
.A(n_12997),
.Y(n_13040)
);

AOI221xp5_ASAP7_75t_L g13041 ( 
.A1(n_13018),
.A2(n_13011),
.B1(n_12987),
.B2(n_12996),
.C(n_12976),
.Y(n_13041)
);

AOI221xp5_ASAP7_75t_L g13042 ( 
.A1(n_12979),
.A2(n_2470),
.B1(n_2468),
.B2(n_2469),
.C(n_2471),
.Y(n_13042)
);

AOI221xp5_ASAP7_75t_L g13043 ( 
.A1(n_13015),
.A2(n_2475),
.B1(n_2473),
.B2(n_2474),
.C(n_2476),
.Y(n_13043)
);

OAI211xp5_ASAP7_75t_L g13044 ( 
.A1(n_13005),
.A2(n_2888),
.B(n_2879),
.C(n_2475),
.Y(n_13044)
);

INVx6_ASAP7_75t_L g13045 ( 
.A(n_12999),
.Y(n_13045)
);

AOI221xp5_ASAP7_75t_L g13046 ( 
.A1(n_13019),
.A2(n_12980),
.B1(n_13007),
.B2(n_12988),
.C(n_13012),
.Y(n_13046)
);

INVx1_ASAP7_75t_L g13047 ( 
.A(n_13017),
.Y(n_13047)
);

OAI21xp33_ASAP7_75t_L g13048 ( 
.A1(n_12985),
.A2(n_2473),
.B(n_2474),
.Y(n_13048)
);

INVx1_ASAP7_75t_L g13049 ( 
.A(n_12977),
.Y(n_13049)
);

OAI311xp33_ASAP7_75t_L g13050 ( 
.A1(n_12982),
.A2(n_2478),
.A3(n_2476),
.B1(n_2477),
.C1(n_2479),
.Y(n_13050)
);

AOI22xp5_ASAP7_75t_L g13051 ( 
.A1(n_13014),
.A2(n_13008),
.B1(n_12991),
.B2(n_13006),
.Y(n_13051)
);

A2O1A1Ixp33_ASAP7_75t_L g13052 ( 
.A1(n_12994),
.A2(n_2479),
.B(n_2477),
.C(n_2478),
.Y(n_13052)
);

INVx1_ASAP7_75t_L g13053 ( 
.A(n_13013),
.Y(n_13053)
);

OAI211xp5_ASAP7_75t_SL g13054 ( 
.A1(n_12985),
.A2(n_2483),
.B(n_2481),
.C(n_2482),
.Y(n_13054)
);

AOI22xp5_ASAP7_75t_L g13055 ( 
.A1(n_12994),
.A2(n_2483),
.B1(n_2481),
.B2(n_2482),
.Y(n_13055)
);

AOI21xp5_ASAP7_75t_L g13056 ( 
.A1(n_12994),
.A2(n_2484),
.B(n_2485),
.Y(n_13056)
);

INVx1_ASAP7_75t_L g13057 ( 
.A(n_13037),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_13028),
.Y(n_13058)
);

INVx1_ASAP7_75t_L g13059 ( 
.A(n_13048),
.Y(n_13059)
);

AOI22xp5_ASAP7_75t_L g13060 ( 
.A1(n_13026),
.A2(n_2488),
.B1(n_2484),
.B2(n_2486),
.Y(n_13060)
);

AO22x1_ASAP7_75t_L g13061 ( 
.A1(n_13029),
.A2(n_2490),
.B1(n_2488),
.B2(n_2489),
.Y(n_13061)
);

NAND3xp33_ASAP7_75t_SL g13062 ( 
.A(n_13031),
.B(n_2497),
.C(n_2489),
.Y(n_13062)
);

AOI22xp5_ASAP7_75t_L g13063 ( 
.A1(n_13024),
.A2(n_2492),
.B1(n_2490),
.B2(n_2491),
.Y(n_13063)
);

INVx1_ASAP7_75t_L g13064 ( 
.A(n_13055),
.Y(n_13064)
);

AOI22xp5_ASAP7_75t_L g13065 ( 
.A1(n_13054),
.A2(n_2494),
.B1(n_2492),
.B2(n_2493),
.Y(n_13065)
);

AOI22xp5_ASAP7_75t_L g13066 ( 
.A1(n_13040),
.A2(n_2496),
.B1(n_2493),
.B2(n_2495),
.Y(n_13066)
);

HB1xp67_ASAP7_75t_L g13067 ( 
.A(n_13036),
.Y(n_13067)
);

CKINVDCx20_ASAP7_75t_R g13068 ( 
.A(n_13033),
.Y(n_13068)
);

AOI22xp5_ASAP7_75t_L g13069 ( 
.A1(n_13049),
.A2(n_2498),
.B1(n_2495),
.B2(n_2496),
.Y(n_13069)
);

INVx1_ASAP7_75t_L g13070 ( 
.A(n_13052),
.Y(n_13070)
);

INVxp67_ASAP7_75t_SL g13071 ( 
.A(n_13032),
.Y(n_13071)
);

INVxp67_ASAP7_75t_L g13072 ( 
.A(n_13038),
.Y(n_13072)
);

INVx2_ASAP7_75t_L g13073 ( 
.A(n_13045),
.Y(n_13073)
);

INVx1_ASAP7_75t_L g13074 ( 
.A(n_13044),
.Y(n_13074)
);

HB1xp67_ASAP7_75t_L g13075 ( 
.A(n_13027),
.Y(n_13075)
);

AOI22xp5_ASAP7_75t_L g13076 ( 
.A1(n_13047),
.A2(n_2500),
.B1(n_2498),
.B2(n_2499),
.Y(n_13076)
);

INVx2_ASAP7_75t_L g13077 ( 
.A(n_13045),
.Y(n_13077)
);

OR2x6_ASAP7_75t_L g13078 ( 
.A(n_13056),
.B(n_2499),
.Y(n_13078)
);

NOR2xp67_ASAP7_75t_L g13079 ( 
.A(n_13035),
.B(n_2500),
.Y(n_13079)
);

INVxp67_ASAP7_75t_SL g13080 ( 
.A(n_13025),
.Y(n_13080)
);

NAND2xp5_ASAP7_75t_SL g13081 ( 
.A(n_13030),
.B(n_2502),
.Y(n_13081)
);

NAND2xp5_ASAP7_75t_L g13082 ( 
.A(n_13042),
.B(n_2895),
.Y(n_13082)
);

INVxp67_ASAP7_75t_SL g13083 ( 
.A(n_13039),
.Y(n_13083)
);

INVx1_ASAP7_75t_L g13084 ( 
.A(n_13051),
.Y(n_13084)
);

INVx1_ASAP7_75t_L g13085 ( 
.A(n_13023),
.Y(n_13085)
);

NAND2xp5_ASAP7_75t_SL g13086 ( 
.A(n_13041),
.B(n_2502),
.Y(n_13086)
);

INVx1_ASAP7_75t_L g13087 ( 
.A(n_13034),
.Y(n_13087)
);

NAND2xp5_ASAP7_75t_SL g13088 ( 
.A(n_13046),
.B(n_2503),
.Y(n_13088)
);

INVx1_ASAP7_75t_L g13089 ( 
.A(n_13053),
.Y(n_13089)
);

INVx1_ASAP7_75t_L g13090 ( 
.A(n_13043),
.Y(n_13090)
);

AOI22xp5_ASAP7_75t_L g13091 ( 
.A1(n_13068),
.A2(n_13050),
.B1(n_2506),
.B2(n_2504),
.Y(n_13091)
);

NOR4xp75_ASAP7_75t_SL g13092 ( 
.A(n_13082),
.B(n_2507),
.C(n_2504),
.D(n_2505),
.Y(n_13092)
);

AND2x2_ASAP7_75t_L g13093 ( 
.A(n_13065),
.B(n_2505),
.Y(n_13093)
);

AND2x2_ASAP7_75t_L g13094 ( 
.A(n_13057),
.B(n_2508),
.Y(n_13094)
);

HB1xp67_ASAP7_75t_L g13095 ( 
.A(n_13061),
.Y(n_13095)
);

CKINVDCx5p33_ASAP7_75t_R g13096 ( 
.A(n_13075),
.Y(n_13096)
);

AOI211xp5_ASAP7_75t_SL g13097 ( 
.A1(n_13072),
.A2(n_2511),
.B(n_2509),
.C(n_2510),
.Y(n_13097)
);

AO22x2_ASAP7_75t_L g13098 ( 
.A1(n_13059),
.A2(n_13074),
.B1(n_13077),
.B2(n_13073),
.Y(n_13098)
);

INVx1_ASAP7_75t_SL g13099 ( 
.A(n_13086),
.Y(n_13099)
);

NAND5xp2_ASAP7_75t_L g13100 ( 
.A(n_13084),
.B(n_2512),
.C(n_2509),
.D(n_2510),
.E(n_2513),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_13078),
.Y(n_13101)
);

NOR2xp33_ASAP7_75t_R g13102 ( 
.A(n_13062),
.B(n_2512),
.Y(n_13102)
);

INVx1_ASAP7_75t_L g13103 ( 
.A(n_13078),
.Y(n_13103)
);

INVx1_ASAP7_75t_L g13104 ( 
.A(n_13088),
.Y(n_13104)
);

NAND4xp25_ASAP7_75t_L g13105 ( 
.A(n_13079),
.B(n_2515),
.C(n_2513),
.D(n_2514),
.Y(n_13105)
);

NOR3xp33_ASAP7_75t_L g13106 ( 
.A(n_13083),
.B(n_2514),
.C(n_2515),
.Y(n_13106)
);

AOI221xp5_ASAP7_75t_L g13107 ( 
.A1(n_13071),
.A2(n_2518),
.B1(n_2516),
.B2(n_2517),
.C(n_2519),
.Y(n_13107)
);

BUFx2_ASAP7_75t_L g13108 ( 
.A(n_13060),
.Y(n_13108)
);

CKINVDCx5p33_ASAP7_75t_R g13109 ( 
.A(n_13067),
.Y(n_13109)
);

INVx2_ASAP7_75t_L g13110 ( 
.A(n_13066),
.Y(n_13110)
);

NAND3x1_ASAP7_75t_SL g13111 ( 
.A(n_13063),
.B(n_13080),
.C(n_13070),
.Y(n_13111)
);

INVxp33_ASAP7_75t_SL g13112 ( 
.A(n_13064),
.Y(n_13112)
);

NAND3xp33_ASAP7_75t_L g13113 ( 
.A(n_13085),
.B(n_2516),
.C(n_2517),
.Y(n_13113)
);

NOR3xp33_ASAP7_75t_L g13114 ( 
.A(n_13087),
.B(n_2518),
.C(n_2519),
.Y(n_13114)
);

NOR2xp33_ASAP7_75t_L g13115 ( 
.A(n_13081),
.B(n_13089),
.Y(n_13115)
);

AND2x4_ASAP7_75t_L g13116 ( 
.A(n_13058),
.B(n_2520),
.Y(n_13116)
);

NAND3xp33_ASAP7_75t_SL g13117 ( 
.A(n_13090),
.B(n_2520),
.C(n_2521),
.Y(n_13117)
);

AND2x4_ASAP7_75t_L g13118 ( 
.A(n_13076),
.B(n_2522),
.Y(n_13118)
);

OAI21xp5_ASAP7_75t_L g13119 ( 
.A1(n_13069),
.A2(n_2522),
.B(n_2524),
.Y(n_13119)
);

OAI22xp5_ASAP7_75t_L g13120 ( 
.A1(n_13065),
.A2(n_2881),
.B1(n_2882),
.B2(n_2880),
.Y(n_13120)
);

XNOR2xp5_ASAP7_75t_L g13121 ( 
.A(n_13068),
.B(n_2525),
.Y(n_13121)
);

CKINVDCx6p67_ASAP7_75t_R g13122 ( 
.A(n_13075),
.Y(n_13122)
);

BUFx6f_ASAP7_75t_L g13123 ( 
.A(n_13073),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_13094),
.Y(n_13124)
);

XNOR2xp5_ASAP7_75t_L g13125 ( 
.A(n_13098),
.B(n_2525),
.Y(n_13125)
);

OAI211xp5_ASAP7_75t_SL g13126 ( 
.A1(n_13099),
.A2(n_2528),
.B(n_2526),
.C(n_2527),
.Y(n_13126)
);

AOI221xp5_ASAP7_75t_L g13127 ( 
.A1(n_13098),
.A2(n_2529),
.B1(n_2526),
.B2(n_2527),
.C(n_2530),
.Y(n_13127)
);

OAI221xp5_ASAP7_75t_L g13128 ( 
.A1(n_13091),
.A2(n_2532),
.B1(n_2529),
.B2(n_2530),
.C(n_2533),
.Y(n_13128)
);

OAI322xp33_ASAP7_75t_L g13129 ( 
.A1(n_13115),
.A2(n_2537),
.A3(n_2536),
.B1(n_2534),
.B2(n_2532),
.C1(n_2533),
.C2(n_2535),
.Y(n_13129)
);

INVx1_ASAP7_75t_L g13130 ( 
.A(n_13121),
.Y(n_13130)
);

AOI221xp5_ASAP7_75t_L g13131 ( 
.A1(n_13120),
.A2(n_2538),
.B1(n_2534),
.B2(n_2536),
.C(n_2539),
.Y(n_13131)
);

NOR2xp33_ASAP7_75t_L g13132 ( 
.A(n_13105),
.B(n_2539),
.Y(n_13132)
);

XNOR2xp5_ASAP7_75t_L g13133 ( 
.A(n_13111),
.B(n_2540),
.Y(n_13133)
);

NAND3xp33_ASAP7_75t_SL g13134 ( 
.A(n_13096),
.B(n_2541),
.C(n_2543),
.Y(n_13134)
);

A2O1A1Ixp33_ASAP7_75t_L g13135 ( 
.A1(n_13097),
.A2(n_2894),
.B(n_2879),
.C(n_2545),
.Y(n_13135)
);

AOI22xp5_ASAP7_75t_L g13136 ( 
.A1(n_13122),
.A2(n_13112),
.B1(n_13123),
.B2(n_13117),
.Y(n_13136)
);

AOI221x1_ASAP7_75t_L g13137 ( 
.A1(n_13104),
.A2(n_2546),
.B1(n_2543),
.B2(n_2544),
.C(n_2547),
.Y(n_13137)
);

AOI22xp5_ASAP7_75t_L g13138 ( 
.A1(n_13123),
.A2(n_2548),
.B1(n_2544),
.B2(n_2547),
.Y(n_13138)
);

A2O1A1Ixp33_ASAP7_75t_L g13139 ( 
.A1(n_13119),
.A2(n_2884),
.B(n_2550),
.C(n_2548),
.Y(n_13139)
);

AOI22xp5_ASAP7_75t_L g13140 ( 
.A1(n_13109),
.A2(n_2551),
.B1(n_2549),
.B2(n_2550),
.Y(n_13140)
);

OAI221xp5_ASAP7_75t_L g13141 ( 
.A1(n_13106),
.A2(n_2553),
.B1(n_2549),
.B2(n_2551),
.C(n_2554),
.Y(n_13141)
);

INVx1_ASAP7_75t_L g13142 ( 
.A(n_13095),
.Y(n_13142)
);

AND2x4_ASAP7_75t_L g13143 ( 
.A(n_13118),
.B(n_2553),
.Y(n_13143)
);

NAND3xp33_ASAP7_75t_SL g13144 ( 
.A(n_13102),
.B(n_2554),
.C(n_2555),
.Y(n_13144)
);

AND3x4_ASAP7_75t_L g13145 ( 
.A(n_13110),
.B(n_2555),
.C(n_2557),
.Y(n_13145)
);

OA21x2_ASAP7_75t_L g13146 ( 
.A1(n_13101),
.A2(n_2568),
.B(n_2557),
.Y(n_13146)
);

AOI22xp5_ASAP7_75t_L g13147 ( 
.A1(n_13093),
.A2(n_2561),
.B1(n_2558),
.B2(n_2560),
.Y(n_13147)
);

OR2x2_ASAP7_75t_L g13148 ( 
.A(n_13100),
.B(n_2560),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_13113),
.Y(n_13149)
);

NOR3xp33_ASAP7_75t_L g13150 ( 
.A(n_13103),
.B(n_2558),
.C(n_2561),
.Y(n_13150)
);

AOI322xp5_ASAP7_75t_L g13151 ( 
.A1(n_13108),
.A2(n_2569),
.A3(n_2568),
.B1(n_2566),
.B2(n_2564),
.C1(n_2565),
.C2(n_2567),
.Y(n_13151)
);

NOR2x1p5_ASAP7_75t_L g13152 ( 
.A(n_13092),
.B(n_2564),
.Y(n_13152)
);

AOI21xp5_ASAP7_75t_L g13153 ( 
.A1(n_13107),
.A2(n_2565),
.B(n_2570),
.Y(n_13153)
);

NAND2xp5_ASAP7_75t_L g13154 ( 
.A(n_13125),
.B(n_13114),
.Y(n_13154)
);

NAND2x1_ASAP7_75t_L g13155 ( 
.A(n_13143),
.B(n_13116),
.Y(n_13155)
);

OR2x2_ASAP7_75t_L g13156 ( 
.A(n_13134),
.B(n_2571),
.Y(n_13156)
);

INVx1_ASAP7_75t_L g13157 ( 
.A(n_13152),
.Y(n_13157)
);

AND2x4_ASAP7_75t_L g13158 ( 
.A(n_13142),
.B(n_2571),
.Y(n_13158)
);

INVx1_ASAP7_75t_L g13159 ( 
.A(n_13133),
.Y(n_13159)
);

NAND2xp33_ASAP7_75t_L g13160 ( 
.A(n_13150),
.B(n_2572),
.Y(n_13160)
);

INVx2_ASAP7_75t_L g13161 ( 
.A(n_13146),
.Y(n_13161)
);

OR2x6_ASAP7_75t_L g13162 ( 
.A(n_13124),
.B(n_2572),
.Y(n_13162)
);

INVx2_ASAP7_75t_L g13163 ( 
.A(n_13146),
.Y(n_13163)
);

INVxp33_ASAP7_75t_L g13164 ( 
.A(n_13132),
.Y(n_13164)
);

AOI21xp5_ASAP7_75t_L g13165 ( 
.A1(n_13144),
.A2(n_2573),
.B(n_2574),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_13148),
.Y(n_13166)
);

INVx2_ASAP7_75t_L g13167 ( 
.A(n_13145),
.Y(n_13167)
);

INVx2_ASAP7_75t_L g13168 ( 
.A(n_13143),
.Y(n_13168)
);

INVx2_ASAP7_75t_L g13169 ( 
.A(n_13138),
.Y(n_13169)
);

NOR2x1p5_ASAP7_75t_L g13170 ( 
.A(n_13130),
.B(n_2573),
.Y(n_13170)
);

NAND2xp5_ASAP7_75t_L g13171 ( 
.A(n_13135),
.B(n_2574),
.Y(n_13171)
);

INVx1_ASAP7_75t_L g13172 ( 
.A(n_13128),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_13140),
.Y(n_13173)
);

OAI22xp5_ASAP7_75t_L g13174 ( 
.A1(n_13157),
.A2(n_13136),
.B1(n_13147),
.B2(n_13139),
.Y(n_13174)
);

INVx1_ASAP7_75t_L g13175 ( 
.A(n_13161),
.Y(n_13175)
);

AND2x2_ASAP7_75t_L g13176 ( 
.A(n_13168),
.B(n_13149),
.Y(n_13176)
);

NOR2xp33_ASAP7_75t_SL g13177 ( 
.A(n_13167),
.B(n_13129),
.Y(n_13177)
);

INVx1_ASAP7_75t_L g13178 ( 
.A(n_13163),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_13170),
.Y(n_13179)
);

INVx1_ASAP7_75t_L g13180 ( 
.A(n_13156),
.Y(n_13180)
);

OAI22x1_ASAP7_75t_L g13181 ( 
.A1(n_13159),
.A2(n_13141),
.B1(n_13126),
.B2(n_13131),
.Y(n_13181)
);

INVx1_ASAP7_75t_L g13182 ( 
.A(n_13171),
.Y(n_13182)
);

OAI22xp5_ASAP7_75t_L g13183 ( 
.A1(n_13154),
.A2(n_13153),
.B1(n_13127),
.B2(n_13137),
.Y(n_13183)
);

NAND2xp5_ASAP7_75t_L g13184 ( 
.A(n_13165),
.B(n_13151),
.Y(n_13184)
);

AOI211xp5_ASAP7_75t_SL g13185 ( 
.A1(n_13166),
.A2(n_2577),
.B(n_2575),
.C(n_2576),
.Y(n_13185)
);

AND3x1_ASAP7_75t_L g13186 ( 
.A(n_13173),
.B(n_2575),
.C(n_2576),
.Y(n_13186)
);

INVx2_ASAP7_75t_L g13187 ( 
.A(n_13162),
.Y(n_13187)
);

OAI22x1_ASAP7_75t_L g13188 ( 
.A1(n_13169),
.A2(n_2579),
.B1(n_2577),
.B2(n_2578),
.Y(n_13188)
);

INVx2_ASAP7_75t_L g13189 ( 
.A(n_13162),
.Y(n_13189)
);

INVx2_ASAP7_75t_L g13190 ( 
.A(n_13158),
.Y(n_13190)
);

INVx1_ASAP7_75t_L g13191 ( 
.A(n_13160),
.Y(n_13191)
);

HB1xp67_ASAP7_75t_L g13192 ( 
.A(n_13155),
.Y(n_13192)
);

NAND2xp5_ASAP7_75t_L g13193 ( 
.A(n_13172),
.B(n_2578),
.Y(n_13193)
);

NAND2xp5_ASAP7_75t_L g13194 ( 
.A(n_13164),
.B(n_2579),
.Y(n_13194)
);

AOI22xp5_ASAP7_75t_L g13195 ( 
.A1(n_13192),
.A2(n_2589),
.B1(n_2597),
.B2(n_2580),
.Y(n_13195)
);

AOI22xp5_ASAP7_75t_L g13196 ( 
.A1(n_13177),
.A2(n_2590),
.B1(n_2598),
.B2(n_2580),
.Y(n_13196)
);

OAI22x1_ASAP7_75t_L g13197 ( 
.A1(n_13187),
.A2(n_2584),
.B1(n_2581),
.B2(n_2583),
.Y(n_13197)
);

OAI22x1_ASAP7_75t_L g13198 ( 
.A1(n_13189),
.A2(n_2585),
.B1(n_2583),
.B2(n_2584),
.Y(n_13198)
);

INVx2_ASAP7_75t_L g13199 ( 
.A(n_13188),
.Y(n_13199)
);

AOI22xp5_ASAP7_75t_L g13200 ( 
.A1(n_13176),
.A2(n_2595),
.B1(n_2603),
.B2(n_2585),
.Y(n_13200)
);

AO22x2_ASAP7_75t_L g13201 ( 
.A1(n_13174),
.A2(n_2588),
.B1(n_2586),
.B2(n_2587),
.Y(n_13201)
);

AOI22xp5_ASAP7_75t_L g13202 ( 
.A1(n_13186),
.A2(n_2597),
.B1(n_2606),
.B2(n_2586),
.Y(n_13202)
);

AOI22xp5_ASAP7_75t_L g13203 ( 
.A1(n_13183),
.A2(n_2599),
.B1(n_2609),
.B2(n_2587),
.Y(n_13203)
);

INVx1_ASAP7_75t_L g13204 ( 
.A(n_13175),
.Y(n_13204)
);

AO22x2_ASAP7_75t_L g13205 ( 
.A1(n_13178),
.A2(n_2592),
.B1(n_2588),
.B2(n_2591),
.Y(n_13205)
);

AOI22xp5_ASAP7_75t_L g13206 ( 
.A1(n_13179),
.A2(n_2602),
.B1(n_2613),
.B2(n_2591),
.Y(n_13206)
);

AOI22xp5_ASAP7_75t_L g13207 ( 
.A1(n_13190),
.A2(n_2603),
.B1(n_2614),
.B2(n_2592),
.Y(n_13207)
);

INVx1_ASAP7_75t_L g13208 ( 
.A(n_13184),
.Y(n_13208)
);

INVx1_ASAP7_75t_L g13209 ( 
.A(n_13193),
.Y(n_13209)
);

OAI22x1_ASAP7_75t_L g13210 ( 
.A1(n_13191),
.A2(n_2596),
.B1(n_2593),
.B2(n_2594),
.Y(n_13210)
);

OAI22x1_ASAP7_75t_L g13211 ( 
.A1(n_13180),
.A2(n_13182),
.B1(n_13194),
.B2(n_13181),
.Y(n_13211)
);

INVx1_ASAP7_75t_L g13212 ( 
.A(n_13185),
.Y(n_13212)
);

OAI22xp5_ASAP7_75t_L g13213 ( 
.A1(n_13192),
.A2(n_2598),
.B1(n_2593),
.B2(n_2596),
.Y(n_13213)
);

OAI22xp5_ASAP7_75t_SL g13214 ( 
.A1(n_13192),
.A2(n_2602),
.B1(n_2600),
.B2(n_2601),
.Y(n_13214)
);

OAI22xp5_ASAP7_75t_L g13215 ( 
.A1(n_13202),
.A2(n_2605),
.B1(n_2600),
.B2(n_2601),
.Y(n_13215)
);

NAND3xp33_ASAP7_75t_SL g13216 ( 
.A(n_13204),
.B(n_2605),
.C(n_2606),
.Y(n_13216)
);

INVx1_ASAP7_75t_L g13217 ( 
.A(n_13212),
.Y(n_13217)
);

INVx2_ASAP7_75t_L g13218 ( 
.A(n_13197),
.Y(n_13218)
);

INVx1_ASAP7_75t_L g13219 ( 
.A(n_13199),
.Y(n_13219)
);

OR3x1_ASAP7_75t_L g13220 ( 
.A(n_13208),
.B(n_2611),
.C(n_2610),
.Y(n_13220)
);

NAND2xp5_ASAP7_75t_SL g13221 ( 
.A(n_13209),
.B(n_2607),
.Y(n_13221)
);

AOI221xp5_ASAP7_75t_L g13222 ( 
.A1(n_13211),
.A2(n_2612),
.B1(n_2610),
.B2(n_2611),
.C(n_2613),
.Y(n_13222)
);

NAND3xp33_ASAP7_75t_SL g13223 ( 
.A(n_13196),
.B(n_2612),
.C(n_2614),
.Y(n_13223)
);

AOI22xp5_ASAP7_75t_L g13224 ( 
.A1(n_13214),
.A2(n_2618),
.B1(n_2615),
.B2(n_2616),
.Y(n_13224)
);

NAND3xp33_ASAP7_75t_L g13225 ( 
.A(n_13203),
.B(n_2615),
.C(n_2616),
.Y(n_13225)
);

OR3x1_ASAP7_75t_L g13226 ( 
.A(n_13198),
.B(n_2620),
.C(n_2619),
.Y(n_13226)
);

NAND3xp33_ASAP7_75t_L g13227 ( 
.A(n_13213),
.B(n_2618),
.C(n_2619),
.Y(n_13227)
);

AND2x4_ASAP7_75t_L g13228 ( 
.A(n_13195),
.B(n_2883),
.Y(n_13228)
);

AOI22xp5_ASAP7_75t_L g13229 ( 
.A1(n_13210),
.A2(n_2622),
.B1(n_2620),
.B2(n_2621),
.Y(n_13229)
);

XOR2xp5_ASAP7_75t_L g13230 ( 
.A(n_13201),
.B(n_2622),
.Y(n_13230)
);

OR3x2_ASAP7_75t_L g13231 ( 
.A(n_13219),
.B(n_13201),
.C(n_13207),
.Y(n_13231)
);

XNOR2xp5_ASAP7_75t_L g13232 ( 
.A(n_13226),
.B(n_13200),
.Y(n_13232)
);

OAI222xp33_ASAP7_75t_L g13233 ( 
.A1(n_13230),
.A2(n_13206),
.B1(n_13205),
.B2(n_2648),
.C1(n_2631),
.C2(n_2656),
.Y(n_13233)
);

XNOR2xp5_ASAP7_75t_L g13234 ( 
.A(n_13220),
.B(n_13205),
.Y(n_13234)
);

NOR2xp33_ASAP7_75t_L g13235 ( 
.A(n_13218),
.B(n_2898),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_13228),
.Y(n_13236)
);

OAI22xp5_ASAP7_75t_L g13237 ( 
.A1(n_13224),
.A2(n_2625),
.B1(n_2626),
.B2(n_2624),
.Y(n_13237)
);

OAI221xp5_ASAP7_75t_L g13238 ( 
.A1(n_13227),
.A2(n_13229),
.B1(n_13225),
.B2(n_13215),
.C(n_13217),
.Y(n_13238)
);

XNOR2xp5_ASAP7_75t_L g13239 ( 
.A(n_13228),
.B(n_2623),
.Y(n_13239)
);

INVx2_ASAP7_75t_L g13240 ( 
.A(n_13221),
.Y(n_13240)
);

AND3x4_ASAP7_75t_L g13241 ( 
.A(n_13223),
.B(n_2627),
.C(n_2628),
.Y(n_13241)
);

INVx2_ASAP7_75t_L g13242 ( 
.A(n_13216),
.Y(n_13242)
);

OR2x2_ASAP7_75t_L g13243 ( 
.A(n_13222),
.B(n_2627),
.Y(n_13243)
);

INVx2_ASAP7_75t_L g13244 ( 
.A(n_13220),
.Y(n_13244)
);

INVxp67_ASAP7_75t_L g13245 ( 
.A(n_13234),
.Y(n_13245)
);

OAI22xp5_ASAP7_75t_L g13246 ( 
.A1(n_13241),
.A2(n_2630),
.B1(n_2628),
.B2(n_2629),
.Y(n_13246)
);

INVx2_ASAP7_75t_L g13247 ( 
.A(n_13239),
.Y(n_13247)
);

OAI22xp5_ASAP7_75t_L g13248 ( 
.A1(n_13231),
.A2(n_2634),
.B1(n_2631),
.B2(n_2633),
.Y(n_13248)
);

BUFx2_ASAP7_75t_L g13249 ( 
.A(n_13243),
.Y(n_13249)
);

O2A1O1Ixp33_ASAP7_75t_L g13250 ( 
.A1(n_13236),
.A2(n_2636),
.B(n_2633),
.C(n_2635),
.Y(n_13250)
);

AOI22x1_ASAP7_75t_L g13251 ( 
.A1(n_13242),
.A2(n_2638),
.B1(n_2639),
.B2(n_2637),
.Y(n_13251)
);

AOI22xp5_ASAP7_75t_L g13252 ( 
.A1(n_13237),
.A2(n_2638),
.B1(n_2635),
.B2(n_2637),
.Y(n_13252)
);

AOI22xp5_ASAP7_75t_L g13253 ( 
.A1(n_13244),
.A2(n_2642),
.B1(n_2640),
.B2(n_2641),
.Y(n_13253)
);

AOI22x1_ASAP7_75t_L g13254 ( 
.A1(n_13240),
.A2(n_2642),
.B1(n_2643),
.B2(n_2641),
.Y(n_13254)
);

INVx1_ASAP7_75t_L g13255 ( 
.A(n_13246),
.Y(n_13255)
);

INVx1_ASAP7_75t_L g13256 ( 
.A(n_13245),
.Y(n_13256)
);

AOI21xp5_ASAP7_75t_L g13257 ( 
.A1(n_13247),
.A2(n_13238),
.B(n_13232),
.Y(n_13257)
);

INVx1_ASAP7_75t_L g13258 ( 
.A(n_13249),
.Y(n_13258)
);

OAI221xp5_ASAP7_75t_L g13259 ( 
.A1(n_13252),
.A2(n_13235),
.B1(n_13233),
.B2(n_2644),
.C(n_2640),
.Y(n_13259)
);

INVx1_ASAP7_75t_SL g13260 ( 
.A(n_13248),
.Y(n_13260)
);

OAI22xp5_ASAP7_75t_L g13261 ( 
.A1(n_13250),
.A2(n_2646),
.B1(n_2643),
.B2(n_2645),
.Y(n_13261)
);

INVx2_ASAP7_75t_L g13262 ( 
.A(n_13251),
.Y(n_13262)
);

OAI322xp33_ASAP7_75t_L g13263 ( 
.A1(n_13256),
.A2(n_13254),
.A3(n_13253),
.B1(n_2652),
.B2(n_2649),
.C1(n_2651),
.C2(n_2645),
.Y(n_13263)
);

XOR2xp5_ASAP7_75t_L g13264 ( 
.A(n_13257),
.B(n_2647),
.Y(n_13264)
);

OAI322xp33_ASAP7_75t_L g13265 ( 
.A1(n_13258),
.A2(n_2655),
.A3(n_2654),
.B1(n_2651),
.B2(n_2647),
.C1(n_2650),
.C2(n_2653),
.Y(n_13265)
);

HB1xp67_ASAP7_75t_L g13266 ( 
.A(n_13259),
.Y(n_13266)
);

INVx1_ASAP7_75t_L g13267 ( 
.A(n_13264),
.Y(n_13267)
);

AO221x2_ASAP7_75t_L g13268 ( 
.A1(n_13266),
.A2(n_13255),
.B1(n_13262),
.B2(n_13261),
.C(n_13260),
.Y(n_13268)
);

OAI331xp33_ASAP7_75t_L g13269 ( 
.A1(n_13267),
.A2(n_13263),
.A3(n_13265),
.B1(n_2659),
.B2(n_2656),
.B3(n_2658),
.C1(n_2654),
.Y(n_13269)
);

AOI22xp5_ASAP7_75t_L g13270 ( 
.A1(n_13269),
.A2(n_13268),
.B1(n_2659),
.B2(n_2655),
.Y(n_13270)
);

NAND3xp33_ASAP7_75t_L g13271 ( 
.A(n_13269),
.B(n_2657),
.C(n_2660),
.Y(n_13271)
);

OR2x6_ASAP7_75t_L g13272 ( 
.A(n_13271),
.B(n_13270),
.Y(n_13272)
);

AOI221xp5_ASAP7_75t_L g13273 ( 
.A1(n_13272),
.A2(n_2662),
.B1(n_2660),
.B2(n_2661),
.C(n_2663),
.Y(n_13273)
);

AOI22xp5_ASAP7_75t_L g13274 ( 
.A1(n_13273),
.A2(n_2665),
.B1(n_2661),
.B2(n_2664),
.Y(n_13274)
);

AOI211xp5_ASAP7_75t_L g13275 ( 
.A1(n_13274),
.A2(n_2667),
.B(n_2664),
.C(n_2666),
.Y(n_13275)
);


endmodule