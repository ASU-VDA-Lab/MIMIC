module real_jpeg_248_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_4),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_69),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_69),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_127),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_6),
.A2(n_54),
.B1(n_56),
.B2(n_127),
.Y(n_249)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_10),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_20),
.B(n_344),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_11),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_12),
.B(n_65),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_12),
.B(n_168),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_12),
.A2(n_13),
.B(n_32),
.C(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_12),
.B(n_37),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_51),
.C(n_54),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_218),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_95),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_12),
.B(n_84),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_32),
.B(n_36),
.C(n_37),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_13),
.B(n_32),
.Y(n_36)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_14),
.A2(n_54),
.B1(n_56),
.B2(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_14),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_15),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_105),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_105),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_15),
.A2(n_54),
.B1(n_56),
.B2(n_105),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_16),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_167),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_16),
.A2(n_54),
.B1(n_56),
.B2(n_167),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_17),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_17),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_17),
.A2(n_43),
.B1(n_54),
.B2(n_56),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_339),
.B(n_342),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_331),
.B(n_335),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_318),
.B(n_330),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_143),
.B(n_315),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_130),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_106),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_26),
.B(n_106),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_87),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_61),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_28),
.A2(n_29),
.B(n_47),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_28),
.B(n_61),
.C(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_30),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_30),
.A2(n_42),
.B1(n_44),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_30),
.A2(n_44),
.B1(n_81),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_30),
.A2(n_184),
.B(n_186),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_30),
.A2(n_186),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_31),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_31),
.A2(n_37),
.B1(n_185),
.B2(n_202),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_31),
.A2(n_37),
.B(n_322),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_32),
.A2(n_33),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g188 ( 
.A1(n_32),
.A2(n_66),
.A3(n_73),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_33),
.B(n_75),
.Y(n_190)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_37),
.B(n_164),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_38),
.A2(n_41),
.B(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_39),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_44),
.A2(n_123),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_44),
.A2(n_163),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_59),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_48),
.A2(n_53),
.B1(n_211),
.B2(n_245),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_48),
.A2(n_213),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_84),
.B1(n_100),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_49),
.A2(n_84),
.B1(n_121),
.B2(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_49),
.A2(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_49),
.B(n_214),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_53),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_53),
.A2(n_234),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_54),
.B(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_78),
.B2(n_86),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_62),
.A2(n_63),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_63),
.B(n_79),
.C(n_83),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_63),
.B(n_134),
.C(n_141),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_72),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_66),
.B1(n_73),
.B2(n_75),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_66),
.A2(n_70),
.B(n_218),
.C(n_227),
.Y(n_226)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_125),
.B(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_72),
.B1(n_77),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_71),
.A2(n_126),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_71),
.A2(n_168),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_71),
.A2(n_168),
.B1(n_325),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_71),
.A2(n_168),
.B(n_333),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_102),
.B(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_82),
.A2(n_83),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_83),
.B(n_135),
.C(n_139),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_84),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_89),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_91),
.B1(n_101),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_96),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_92),
.A2(n_95),
.B1(n_118),
.B2(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_92),
.A2(n_218),
.B(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_93),
.A2(n_94),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_93),
.A2(n_94),
.B1(n_193),
.B2(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_93),
.B(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_93),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_93),
.A2(n_94),
.B1(n_249),
.B2(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_94),
.A2(n_208),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_94),
.B(n_222),
.Y(n_251)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_95),
.A2(n_221),
.B(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_98),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_113),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.C(n_124),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_115),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_124),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_129),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_130),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_142),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_131),
.B(n_142),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_136),
.Y(n_324)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_140),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_169),
.B(n_314),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_145),
.B(n_148),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.C(n_165),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_156),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_157),
.B(n_159),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_195),
.B(n_313),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_171),
.B(n_173),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_180),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_174),
.B(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_180),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_187),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_181),
.B(n_183),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_187),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI31xp33_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_295),
.A3(n_305),
.B(n_310),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_239),
.B(n_294),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_223),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_198),
.B(n_223),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.C(n_215),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_199),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_215),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_219),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_224),
.B(n_236),
.C(n_238),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_225),
.B(n_230),
.C(n_231),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_289),
.B(n_293),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_258),
.B(n_288),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_248),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_270),
.B(n_287),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_281),
.B(n_286),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_276),
.B(n_280),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_279),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_329),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_326),
.C(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_340),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_334),
.Y(n_338)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_341),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule