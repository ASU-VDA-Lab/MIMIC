module real_aes_17915_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_103;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_0), .Y(n_230) );
AND2x4_ASAP7_75t_L g106 ( .A(n_1), .B(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g161 ( .A(n_2), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_3), .Y(n_864) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_5), .B(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g113 ( .A(n_6), .B(n_21), .Y(n_113) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_7), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_8), .A2(n_52), .B1(n_128), .B2(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_8), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_9), .B(n_150), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_10), .B(n_150), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_11), .B(n_198), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_12), .A2(n_81), .B1(n_150), .B2(n_152), .Y(n_249) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_13), .A2(n_36), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_14), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_15), .B(n_188), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_16), .Y(n_611) );
AO32x2_ASAP7_75t_L g246 ( .A1(n_17), .A2(n_141), .A3(n_142), .B1(n_247), .B2(n_250), .Y(n_246) );
AO32x1_ASAP7_75t_L g268 ( .A1(n_17), .A2(n_141), .A3(n_142), .B1(n_247), .B2(n_250), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_18), .B(n_574), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_19), .B(n_141), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_20), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_22), .B(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_23), .A2(n_42), .B1(n_157), .B2(n_188), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_24), .A2(n_90), .B1(n_152), .B2(n_158), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_25), .B(n_172), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_26), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_27), .B(n_205), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_28), .A2(n_61), .B1(n_887), .B2(n_888), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_28), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_29), .A2(n_63), .B1(n_158), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_30), .B(n_150), .Y(n_563) );
INVx2_ASAP7_75t_L g118 ( .A(n_31), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_32), .B(n_154), .Y(n_584) );
BUFx3_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g870 ( .A(n_33), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_34), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_35), .B(n_541), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_37), .B(n_541), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_38), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_39), .B(n_204), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_40), .B(n_574), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_41), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_43), .B(n_553), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_44), .A2(n_76), .B1(n_204), .B2(n_205), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_45), .B(n_239), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_46), .A2(n_189), .B(n_228), .C(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_47), .A2(n_78), .B1(n_150), .B2(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g144 ( .A(n_48), .Y(n_144) );
AND2x4_ASAP7_75t_L g146 ( .A(n_49), .B(n_147), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_50), .A2(n_51), .B1(n_157), .B2(n_158), .Y(n_576) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_52), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_53), .B(n_141), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_54), .B(n_541), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_55), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_56), .B(n_158), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_57), .B(n_152), .Y(n_168) );
INVx1_ASAP7_75t_L g147 ( .A(n_58), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_59), .B(n_141), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_60), .A2(n_228), .B(n_229), .C(n_231), .Y(n_227) );
INVx1_ASAP7_75t_SL g887 ( .A(n_61), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g176 ( .A(n_62), .B(n_152), .C(n_174), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_64), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_65), .B(n_141), .Y(n_567) );
AND2x2_ASAP7_75t_L g233 ( .A(n_66), .B(n_234), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_67), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_68), .B(n_522), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_69), .B(n_154), .C(n_188), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_70), .A2(n_93), .B1(n_150), .B2(n_204), .Y(n_208) );
INVx2_ASAP7_75t_L g155 ( .A(n_71), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_72), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_73), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_74), .B(n_207), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_75), .B(n_150), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_77), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_79), .B(n_192), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_80), .A2(n_88), .B1(n_573), .B2(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_82), .B(n_150), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_83), .B(n_174), .Y(n_173) );
NAND2xp33_ASAP7_75t_SL g539 ( .A(n_84), .B(n_170), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_85), .B(n_186), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_86), .A2(n_100), .B1(n_157), .B2(n_158), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_87), .B(n_205), .Y(n_256) );
INVx1_ASAP7_75t_L g891 ( .A(n_89), .Y(n_891) );
INVx1_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_91), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_92), .B(n_198), .Y(n_262) );
NAND2xp33_ASAP7_75t_L g523 ( .A(n_94), .B(n_170), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_95), .B(n_541), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_96), .B(n_170), .C(n_207), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_97), .B(n_522), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_98), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_99), .B(n_574), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_114), .B(n_890), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
BUFx8_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g892 ( .A(n_105), .Y(n_892) );
AND2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_L g877 ( .A(n_108), .Y(n_877) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
BUFx8_ASAP7_75t_SL g507 ( .A(n_109), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_109), .Y(n_860) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g120 ( .A(n_112), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_113), .Y(n_121) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_122), .B(n_861), .Y(n_114) );
BUFx12f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_SL g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_118), .B(n_877), .Y(n_876) );
INVx3_ASAP7_75t_L g882 ( .A(n_118), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x6_ASAP7_75t_SL g867 ( .A(n_121), .B(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_505), .B1(n_508), .B2(n_859), .Y(n_130) );
XOR2xp5_ASAP7_75t_L g885 ( .A(n_131), .B(n_886), .Y(n_885) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_406), .Y(n_131) );
AND4x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_328), .C(n_361), .D(n_392), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_295), .Y(n_133) );
OAI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_214), .B1(n_263), .B2(n_273), .C(n_282), .Y(n_134) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_135), .A2(n_385), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_178), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_162), .Y(n_137) );
INVx2_ASAP7_75t_L g281 ( .A(n_138), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_138), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g327 ( .A(n_138), .B(n_200), .Y(n_327) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g316 ( .A(n_139), .Y(n_316) );
AOI31xp67_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .A3(n_148), .B(n_159), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_142), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
BUFx3_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_142), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_SL g253 ( .A(n_142), .Y(n_253) );
AND2x4_ASAP7_75t_SL g528 ( .A(n_142), .B(n_145), .Y(n_528) );
INVx1_ASAP7_75t_SL g532 ( .A(n_142), .Y(n_532) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_145), .A2(n_167), .B(n_171), .Y(n_166) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_183), .B(n_190), .Y(n_182) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_534), .B(n_537), .Y(n_533) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_145), .A2(n_547), .B(n_550), .Y(n_546) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_145), .A2(n_561), .B(n_564), .Y(n_560) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_145), .A2(n_583), .B(n_586), .Y(n_582) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_145), .A2(n_640), .B(n_643), .Y(n_639) );
BUFx10_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
INVx1_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_146), .A2(n_201), .A3(n_237), .B(n_242), .Y(n_236) );
BUFx10_ASAP7_75t_L g578 ( .A(n_146), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B1(n_154), .B2(n_156), .Y(n_148) );
INVx3_ASAP7_75t_L g261 ( .A(n_150), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_150), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g589 ( .A(n_150), .Y(n_589) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_151), .Y(n_152) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx1_ASAP7_75t_L g204 ( .A(n_151), .Y(n_204) );
INVx1_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
INVx3_ASAP7_75t_L g522 ( .A(n_151), .Y(n_522) );
INVx1_ASAP7_75t_L g575 ( .A(n_151), .Y(n_575) );
INVx2_ASAP7_75t_SL g205 ( .A(n_152), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_152), .B(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_153), .A2(n_203), .B1(n_206), .B2(n_208), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_153), .A2(n_238), .B1(n_240), .B2(n_241), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_153), .A2(n_259), .B(n_260), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_153), .A2(n_572), .B1(n_576), .B2(n_577), .Y(n_571) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_154), .A2(n_168), .B(n_169), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_154), .A2(n_189), .B1(n_248), .B2(n_249), .Y(n_247) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_185), .B(n_548), .C(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_154), .A2(n_565), .B(n_566), .Y(n_564) );
BUFx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
INVx1_ASAP7_75t_L g207 ( .A(n_155), .Y(n_207) );
INVx1_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_157), .A2(n_188), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g172 ( .A(n_158), .Y(n_172) );
INVx2_ASAP7_75t_L g573 ( .A(n_158), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_158), .A2(n_584), .B(n_585), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_158), .A2(n_522), .B1(n_614), .B2(n_615), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g302 ( .A(n_162), .B(n_292), .Y(n_302) );
OR2x2_ASAP7_75t_L g411 ( .A(n_162), .B(n_180), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_177), .Y(n_162) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_163), .A2(n_166), .B(n_177), .Y(n_280) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_163), .A2(n_546), .B(n_554), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_163), .A2(n_546), .B(n_554), .Y(n_627) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_163), .A2(n_639), .B(n_646), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g664 ( .A1(n_163), .A2(n_639), .B(n_646), .Y(n_664) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g541 ( .A(n_164), .Y(n_541) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx2_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
INVx2_ASAP7_75t_L g553 ( .A(n_170), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_176), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_178), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_200), .Y(n_179) );
INVx1_ASAP7_75t_L g276 ( .A(n_180), .Y(n_276) );
INVx2_ASAP7_75t_SL g353 ( .A(n_180), .Y(n_353) );
BUFx2_ASAP7_75t_L g383 ( .A(n_180), .Y(n_383) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_197), .Y(n_180) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_181), .A2(n_182), .B(n_197), .Y(n_292) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_181), .A2(n_560), .B(n_567), .Y(n_559) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_181), .A2(n_582), .B(n_590), .Y(n_581) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_181), .A2(n_560), .B(n_567), .Y(n_597) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_181), .A2(n_582), .B(n_590), .Y(n_626) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_189), .Y(n_183) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_189), .A2(n_521), .B(n_523), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_189), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_189), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_189), .A2(n_641), .B(n_642), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B1(n_195), .B2(n_196), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_192), .A2(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_193), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_524) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx3_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
INVx2_ASAP7_75t_L g220 ( .A(n_198), .Y(n_220) );
NOR2xp67_ASAP7_75t_SL g606 ( .A(n_198), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_199), .A2(n_571), .A3(n_578), .B(n_579), .Y(n_570) );
AND2x2_ASAP7_75t_L g275 ( .A(n_200), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g294 ( .A(n_200), .Y(n_294) );
OR2x2_ASAP7_75t_L g314 ( .A(n_200), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g355 ( .A(n_200), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_200), .Y(n_366) );
AND2x2_ASAP7_75t_L g373 ( .A(n_200), .B(n_315), .Y(n_373) );
AO31x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .A3(n_209), .B(n_211), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_204), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_SL g250 ( .A(n_210), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_213), .B(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_216), .B(n_244), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_235), .Y(n_216) );
INVx1_ASAP7_75t_L g287 ( .A(n_217), .Y(n_287) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
INVx1_ASAP7_75t_L g308 ( .A(n_218), .Y(n_308) );
INVx1_ASAP7_75t_L g347 ( .A(n_218), .Y(n_347) );
AND2x2_ASAP7_75t_L g377 ( .A(n_218), .B(n_236), .Y(n_377) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g271 ( .A(n_219), .Y(n_271) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_233), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_227), .B(n_232), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_226), .Y(n_222) );
AOI21x1_ASAP7_75t_L g586 ( .A1(n_226), .A2(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g526 ( .A(n_228), .Y(n_526) );
INVx2_ASAP7_75t_L g241 ( .A(n_231), .Y(n_241) );
INVx2_ASAP7_75t_L g577 ( .A(n_231), .Y(n_577) );
INVx1_ASAP7_75t_L g283 ( .A(n_235), .Y(n_283) );
AND2x4_ASAP7_75t_L g332 ( .A(n_235), .B(n_246), .Y(n_332) );
AND2x2_ASAP7_75t_L g342 ( .A(n_235), .B(n_271), .Y(n_342) );
INVx1_ASAP7_75t_L g403 ( .A(n_235), .Y(n_403) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g289 ( .A(n_236), .B(n_268), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_236), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g323 ( .A(n_236), .B(n_268), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_236), .B(n_251), .Y(n_432) );
AOI21x1_ASAP7_75t_L g255 ( .A1(n_241), .A2(n_256), .B(n_257), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_241), .A2(n_644), .B(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_244), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
OR2x2_ASAP7_75t_L g449 ( .A(n_245), .B(n_251), .Y(n_449) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g396 ( .A(n_246), .Y(n_396) );
AND2x2_ASAP7_75t_L g421 ( .A(n_246), .B(n_251), .Y(n_421) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_250), .A2(n_255), .B(n_258), .Y(n_254) );
INVx3_ASAP7_75t_L g272 ( .A(n_251), .Y(n_272) );
AND2x2_ASAP7_75t_L g298 ( .A(n_251), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
INVx1_ASAP7_75t_L g334 ( .A(n_251), .Y(n_334) );
INVx1_ASAP7_75t_L g344 ( .A(n_251), .Y(n_344) );
BUFx2_ASAP7_75t_L g439 ( .A(n_251), .Y(n_439) );
OR2x2_ASAP7_75t_L g467 ( .A(n_251), .B(n_271), .Y(n_467) );
INVxp67_ASAP7_75t_L g484 ( .A(n_251), .Y(n_484) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_262), .Y(n_252) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
AND2x4_ASAP7_75t_L g297 ( .A(n_265), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_265), .B(n_377), .Y(n_458) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g285 ( .A(n_267), .B(n_272), .Y(n_285) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_267), .Y(n_309) );
INVx1_ASAP7_75t_L g433 ( .A(n_267), .Y(n_433) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g346 ( .A(n_268), .Y(n_346) );
AND2x2_ASAP7_75t_L g360 ( .A(n_269), .B(n_323), .Y(n_360) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
OR2x2_ASAP7_75t_L g380 ( .A(n_271), .B(n_346), .Y(n_380) );
INVx1_ASAP7_75t_L g443 ( .A(n_271), .Y(n_443) );
AND2x2_ASAP7_75t_L g386 ( .A(n_272), .B(n_332), .Y(n_386) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
AND2x2_ASAP7_75t_L g389 ( .A(n_275), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
AND2x2_ASAP7_75t_L g293 ( .A(n_278), .B(n_294), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_278), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g391 ( .A(n_280), .B(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g354 ( .A(n_281), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g425 ( .A(n_281), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_286), .C(n_290), .Y(n_282) );
INVx1_ASAP7_75t_L g417 ( .A(n_284), .Y(n_417) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g413 ( .A(n_285), .B(n_377), .Y(n_413) );
INVx1_ASAP7_75t_L g504 ( .A(n_285), .Y(n_504) );
INVx1_ASAP7_75t_L g469 ( .A(n_286), .Y(n_469) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g502 ( .A(n_287), .B(n_421), .Y(n_502) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g319 ( .A(n_289), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g474 ( .A(n_289), .B(n_439), .Y(n_474) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVxp67_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_291), .B(n_326), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_291), .B(n_293), .Y(n_456) );
INVx1_ASAP7_75t_L g339 ( .A(n_292), .Y(n_339) );
INVx2_ASAP7_75t_SL g304 ( .A(n_294), .Y(n_304) );
OR2x2_ASAP7_75t_L g333 ( .A(n_294), .B(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B1(n_305), .B2(n_310), .C(n_317), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_297), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g369 ( .A(n_299), .Y(n_369) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g426 ( .A(n_302), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_302), .B(n_304), .Y(n_464) );
OR2x2_ASAP7_75t_L g446 ( .A(n_303), .B(n_436), .Y(n_446) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g415 ( .A(n_304), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g462 ( .A(n_304), .B(n_391), .Y(n_462) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
AND2x2_ASAP7_75t_L g397 ( .A(n_307), .B(n_320), .Y(n_397) );
BUFx2_ASAP7_75t_L g423 ( .A(n_307), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_311), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g326 ( .A(n_312), .Y(n_326) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g399 ( .A(n_314), .Y(n_399) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_324), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_320), .Y(n_379) );
OR2x2_ASAP7_75t_L g489 ( .A(n_320), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g450 ( .A(n_321), .Y(n_450) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
AND2x2_ASAP7_75t_L g485 ( .A(n_323), .B(n_358), .Y(n_485) );
INVx2_ASAP7_75t_SL g490 ( .A(n_323), .Y(n_490) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g372 ( .A(n_326), .Y(n_372) );
AND2x4_ASAP7_75t_L g348 ( .A(n_327), .B(n_337), .Y(n_348) );
INVx2_ASAP7_75t_L g412 ( .A(n_327), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_327), .B(n_353), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_327), .B(n_383), .Y(n_499) );
AOI221x1_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_335), .B1(n_340), .B2(n_348), .C(n_349), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx2_ASAP7_75t_L g468 ( .A(n_331), .Y(n_468) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_331), .A2(n_476), .B(n_478), .Y(n_475) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g388 ( .A(n_332), .Y(n_388) );
AND2x4_ASAP7_75t_L g442 ( .A(n_332), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g402 ( .A(n_334), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI32xp33_ASAP7_75t_L g447 ( .A1(n_336), .A2(n_445), .A3(n_448), .B1(n_450), .B2(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_337), .B(n_354), .Y(n_470) );
AND2x2_ASAP7_75t_L g486 ( .A(n_337), .B(n_366), .Y(n_486) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_341), .B(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_342), .B(n_484), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_343), .A2(n_419), .B(n_422), .C(n_424), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_356), .B(n_359), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_350), .A2(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_353), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_357), .A2(n_430), .B1(n_434), .B2(n_435), .Y(n_429) );
AND2x2_ASAP7_75t_L g496 ( .A(n_357), .B(n_484), .Y(n_496) );
NOR2xp33_ASAP7_75t_SL g361 ( .A(n_362), .B(n_384), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_374), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_363), .A2(n_473), .B(n_474), .Y(n_472) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g455 ( .A(n_369), .B(n_421), .Y(n_455) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AOI31xp33_ASAP7_75t_L g392 ( .A1(n_372), .A2(n_393), .A3(n_398), .B(n_400), .Y(n_392) );
AND2x2_ASAP7_75t_L g492 ( .A(n_372), .B(n_399), .Y(n_492) );
AND2x2_ASAP7_75t_L g381 ( .A(n_373), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_373), .Y(n_445) );
INVx1_ASAP7_75t_L g479 ( .A(n_373), .Y(n_479) );
OAI21xp33_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_378), .B(n_381), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_377), .B(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_378), .A2(n_461), .B(n_463), .Y(n_460) );
NOR2x1p5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_380), .A2(n_395), .B(n_402), .C(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g414 ( .A(n_383), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g434 ( .A(n_383), .B(n_390), .Y(n_434) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx1_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_414), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g473 ( .A(n_397), .Y(n_473) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_459), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_427), .C(n_437), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_414), .B2(n_417), .C(n_418), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_415), .A2(n_482), .B1(n_485), .B2(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OR2x2_ASAP7_75t_L g478 ( .A(n_426), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g477 ( .A(n_432), .Y(n_477) );
INVx2_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_447), .C(n_453), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g448 ( .A(n_443), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g491 ( .A(n_448), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND4xp75_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_480), .D(n_493), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_469), .B2(n_470), .Y(n_463) );
NAND2x1_ASAP7_75t_SL g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_487), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B(n_492), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B1(n_497), .B2(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_791), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_666), .C(n_706), .D(n_755), .Y(n_510) );
NOR2xp67_ASAP7_75t_L g511 ( .A(n_512), .B(n_617), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_542), .B1(n_591), .B2(n_600), .Y(n_512) );
INVx1_ASAP7_75t_L g787 ( .A(n_513), .Y(n_787) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_514), .B(n_636), .Y(n_703) );
AND2x2_ASAP7_75t_L g734 ( .A(n_514), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_529), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_515), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g658 ( .A(n_515), .Y(n_658) );
AND2x2_ASAP7_75t_L g833 ( .A(n_515), .B(n_701), .Y(n_833) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g602 ( .A(n_516), .Y(n_602) );
AND2x2_ASAP7_75t_L g686 ( .A(n_516), .B(n_648), .Y(n_686) );
AND2x2_ASAP7_75t_L g730 ( .A(n_516), .B(n_637), .Y(n_730) );
OR2x2_ASAP7_75t_L g748 ( .A(n_516), .B(n_749), .Y(n_748) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g652 ( .A(n_517), .B(n_637), .Y(n_652) );
BUFx2_ASAP7_75t_L g709 ( .A(n_517), .Y(n_709) );
OR2x2_ASAP7_75t_L g717 ( .A(n_517), .B(n_675), .Y(n_717) );
INVx1_ASAP7_75t_L g772 ( .A(n_517), .Y(n_772) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_524), .B(n_528), .Y(n_519) );
AND2x2_ASAP7_75t_L g603 ( .A(n_529), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g711 ( .A(n_529), .B(n_688), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_529), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g749 ( .A(n_530), .Y(n_749) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_530), .Y(n_754) );
AND2x2_ASAP7_75t_L g771 ( .A(n_530), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g661 ( .A(n_531), .B(n_605), .Y(n_661) );
INVx1_ASAP7_75t_L g675 ( .A(n_531), .Y(n_675) );
OAI21x1_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_540), .Y(n_531) );
NAND2x1_ASAP7_75t_L g542 ( .A(n_543), .B(n_555), .Y(n_542) );
AND2x4_ASAP7_75t_L g836 ( .A(n_543), .B(n_764), .Y(n_836) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_544), .Y(n_599) );
BUFx3_ASAP7_75t_L g632 ( .A(n_544), .Y(n_632) );
INVx1_ASAP7_75t_L g696 ( .A(n_544), .Y(n_696) );
AND2x2_ASAP7_75t_L g699 ( .A(n_544), .B(n_558), .Y(n_699) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_581), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_544), .Y(n_727) );
AND2x2_ASAP7_75t_L g759 ( .A(n_544), .B(n_626), .Y(n_759) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_568), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g668 ( .A(n_557), .B(n_654), .Y(n_668) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g694 ( .A(n_559), .B(n_681), .Y(n_694) );
AND2x2_ASAP7_75t_L g723 ( .A(n_559), .B(n_570), .Y(n_723) );
OR2x2_ASAP7_75t_L g819 ( .A(n_559), .B(n_570), .Y(n_819) );
AND2x2_ASAP7_75t_L g698 ( .A(n_568), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g847 ( .A(n_568), .Y(n_847) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_569), .Y(n_593) );
OR2x2_ASAP7_75t_L g781 ( .A(n_569), .B(n_595), .Y(n_781) );
INVx1_ASAP7_75t_L g803 ( .A(n_569), .Y(n_803) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_581), .Y(n_569) );
AND2x2_ASAP7_75t_L g621 ( .A(n_570), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g654 ( .A(n_570), .B(n_626), .Y(n_654) );
INVx1_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_570), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_570), .B(n_581), .Y(n_768) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_577), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g607 ( .A(n_578), .Y(n_607) );
AND2x2_ASAP7_75t_L g705 ( .A(n_581), .B(n_627), .Y(n_705) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR3x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .C(n_598), .Y(n_592) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_595), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g653 ( .A(n_595), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g704 ( .A(n_595), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g744 ( .A(n_595), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_595), .B(n_767), .Y(n_799) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g740 ( .A(n_596), .B(n_680), .Y(n_740) );
AND2x2_ASAP7_75t_L g764 ( .A(n_596), .B(n_626), .Y(n_764) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g775 ( .A(n_599), .B(n_654), .Y(n_775) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_602), .B(n_661), .Y(n_840) );
AND2x4_ASAP7_75t_L g832 ( .A(n_603), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_603), .B(n_652), .Y(n_846) );
INVx2_ASAP7_75t_L g648 ( .A(n_604), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_604), .Y(n_651) );
INVx2_ASAP7_75t_L g736 ( .A(n_604), .Y(n_736) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g720 ( .A(n_605), .Y(n_720) );
AOI21x1_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_616), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_655), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_633), .B1(n_649), .B2(n_653), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_628), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g683 ( .A(n_621), .B(n_632), .Y(n_683) );
AND2x2_ASAP7_75t_L g843 ( .A(n_621), .B(n_724), .Y(n_843) );
BUFx2_ASAP7_75t_L g714 ( .A(n_622), .Y(n_714) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g713 ( .A(n_625), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g630 ( .A(n_626), .Y(n_630) );
INVx1_ASAP7_75t_L g680 ( .A(n_626), .Y(n_680) );
INVx1_ASAP7_75t_L g805 ( .A(n_627), .Y(n_805) );
AOI31xp33_ASAP7_75t_L g823 ( .A1(n_628), .A2(n_824), .A3(n_825), .B(n_826), .Y(n_823) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_630), .B(n_723), .Y(n_822) );
INVx2_ASAP7_75t_L g850 ( .A(n_630), .Y(n_850) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_631), .Y(n_665) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g678 ( .A(n_632), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_632), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g808 ( .A(n_632), .B(n_768), .Y(n_808) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_647), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g719 ( .A(n_637), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g688 ( .A(n_638), .Y(n_688) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_651), .Y(n_672) );
INVx1_ASAP7_75t_L g712 ( .A(n_651), .Y(n_712) );
INVx1_ASAP7_75t_L g692 ( .A(n_652), .Y(n_692) );
AND2x2_ASAP7_75t_L g753 ( .A(n_652), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g809 ( .A(n_652), .B(n_736), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_653), .A2(n_726), .B(n_728), .Y(n_725) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_665), .Y(n_655) );
NAND3x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .C(n_662), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g827 ( .A(n_658), .B(n_747), .Y(n_827) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_SL g780 ( .A(n_660), .B(n_692), .Y(n_780) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g700 ( .A(n_661), .B(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_662), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_662), .B(n_771), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_662), .B(n_771), .Y(n_844) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g747 ( .A(n_664), .B(n_720), .Y(n_747) );
AND2x2_ASAP7_75t_L g667 ( .A(n_665), .B(n_668), .Y(n_667) );
AOI221x1_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_669), .B1(n_676), .B2(n_685), .C(n_689), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g848 ( .A1(n_668), .A2(n_849), .A3(n_854), .B1(n_855), .B2(n_857), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_673), .B(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g687 ( .A(n_675), .B(n_688), .Y(n_687) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_675), .Y(n_691) );
OR2x2_ASAP7_75t_L g804 ( .A(n_675), .B(n_805), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .C(n_684), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g726 ( .A(n_679), .B(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g743 ( .A(n_679), .B(n_744), .Y(n_743) );
AND2x4_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_682), .A2(n_779), .B1(n_781), .B2(n_782), .Y(n_778) );
INVx3_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g856 ( .A(n_686), .Y(n_856) );
INVx2_ASAP7_75t_L g701 ( .A(n_688), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_697), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g825 ( .A(n_694), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_695), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_702), .B2(n_704), .Y(n_697) );
AND2x4_ASAP7_75t_L g794 ( .A(n_700), .B(n_709), .Y(n_794) );
INVx1_ASAP7_75t_L g853 ( .A(n_701), .Y(n_853) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g732 ( .A(n_705), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_705), .B(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_705), .B(n_733), .Y(n_824) );
AOI211x1_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_713), .B(n_715), .C(n_741), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR3x2_ASAP7_75t_L g816 ( .A(n_709), .B(n_711), .C(n_712), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_710), .A2(n_732), .B1(n_734), .B2(n_737), .Y(n_731) );
NOR2x1p5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_712), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_711), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
INVx2_ASAP7_75t_L g733 ( .A(n_714), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_721), .B(n_725), .C(n_731), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_723), .B(n_727), .Y(n_738) );
INVx1_ASAP7_75t_L g765 ( .A(n_723), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_723), .B(n_830), .Y(n_838) );
OAI32xp33_ASAP7_75t_L g813 ( .A1(n_724), .A2(n_769), .A3(n_814), .B1(n_816), .B2(n_817), .Y(n_813) );
INVx1_ASAP7_75t_L g830 ( .A(n_724), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_724), .B(n_744), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_727), .B(n_761), .Y(n_796) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g774 ( .A(n_733), .B(n_759), .Y(n_774) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g783 ( .A(n_736), .B(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g751 ( .A(n_739), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B1(n_750), .B2(n_752), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g789 ( .A(n_746), .Y(n_789) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g770 ( .A(n_747), .B(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_747), .B(n_754), .Y(n_858) );
INVx1_ASAP7_75t_SL g784 ( .A(n_748), .Y(n_784) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_778), .C(n_785), .Y(n_755) );
OAI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_769), .B(n_773), .Y(n_756) );
NOR2xp33_ASAP7_75t_SL g757 ( .A(n_758), .B(n_762), .Y(n_757) );
INVxp67_ASAP7_75t_L g790 ( .A(n_758), .Y(n_790) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g815 ( .A(n_760), .Y(n_815) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .C(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g777 ( .A(n_771), .Y(n_777) );
OAI21xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g786 ( .A(n_774), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_779), .A2(n_830), .B1(n_831), .B2(n_834), .C(n_835), .Y(n_829) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI32xp33_ASAP7_75t_L g785 ( .A1(n_782), .A2(n_786), .A3(n_787), .B1(n_788), .B2(n_790), .Y(n_785) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_788), .A2(n_798), .B1(n_799), .B2(n_800), .C(n_806), .Y(n_797) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_810), .C(n_828), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B(n_797), .Y(n_792) );
AOI211x1_ASAP7_75t_L g810 ( .A1(n_793), .A2(n_811), .B(n_813), .C(n_820), .Y(n_810) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2x1_ASAP7_75t_SL g801 ( .A(n_802), .B(n_804), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g812 ( .A(n_803), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AO21x1_ASAP7_75t_L g820 ( .A1(n_809), .A2(n_821), .B(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g854 ( .A(n_825), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_841), .Y(n_828) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI21xp33_ASAP7_75t_SL g835 ( .A1(n_836), .A2(n_837), .B(n_839), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_848), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B(n_845), .Y(n_842) );
NOR2xp67_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g851 ( .A(n_850), .Y(n_851) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx12f_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_878), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_871), .Y(n_862) );
INVxp67_ASAP7_75t_L g889 ( .A(n_863), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_865), .B(n_885), .Y(n_884) );
BUFx12f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx4_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx6_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx10_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_883), .Y(n_878) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
CKINVDCx11_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
BUFx6f_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_889), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
endmodule