module fake_netlist_1_12703_n_782 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_782);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_782;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_96), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
BUFx5_ASAP7_75t_L g103 ( .A(n_100), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_59), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_49), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_68), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_64), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
BUFx10_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_4), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_53), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_28), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_56), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_38), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_42), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_93), .Y(n_121) );
INVxp33_ASAP7_75t_L g122 ( .A(n_95), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_70), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_29), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_32), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_76), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_22), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_1), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_25), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_47), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_7), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_52), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_58), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_9), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_43), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_16), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_7), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_37), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_107), .B(n_0), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_122), .B(n_0), .Y(n_145) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_124), .A2(n_50), .B(n_98), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_132), .B(n_1), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_131), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
INVx2_ASAP7_75t_SL g152 ( .A(n_124), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_103), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_126), .A2(n_127), .B(n_112), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_109), .B(n_2), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_102), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_103), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_103), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_122), .B(n_113), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_113), .B(n_2), .Y(n_161) );
OR2x6_ASAP7_75t_L g162 ( .A(n_160), .B(n_135), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_145), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_160), .B(n_114), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_141), .B(n_126), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_161), .B(n_135), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_161), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_141), .B(n_119), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_142), .B(n_139), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_142), .B(n_129), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_143), .B(n_119), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_154), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_143), .B(n_111), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_163), .B(n_149), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_162), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_165), .B(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_189), .B(n_154), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_177), .B(n_155), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_177), .B(n_155), .Y(n_202) );
OR2x6_ASAP7_75t_L g203 ( .A(n_162), .B(n_102), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_179), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_195), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_171), .B(n_162), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_164), .B(n_115), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_168), .B(n_106), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_196), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_169), .B(n_101), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_183), .B(n_104), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_196), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_182), .B(n_117), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_193), .B(n_103), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_169), .B(n_116), .Y(n_216) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_102), .B1(n_136), .B2(n_120), .C(n_121), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_169), .B(n_118), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_194), .B(n_123), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_186), .B(n_133), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_191), .B(n_134), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_185), .B(n_130), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_185), .B(n_125), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_196), .A2(n_146), .B1(n_102), .B2(n_138), .Y(n_225) );
AND2x4_ASAP7_75t_SL g226 ( .A(n_185), .B(n_128), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g228 ( .A(n_166), .B(n_146), .C(n_137), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_192), .B(n_140), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_192), .B(n_127), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_192), .B(n_146), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_170), .A2(n_174), .B1(n_188), .B2(n_172), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_172), .Y(n_235) );
AND2x6_ASAP7_75t_SL g236 ( .A(n_173), .B(n_3), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_173), .B(n_146), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_174), .B(n_146), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_175), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_175), .B(n_157), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_216), .B(n_176), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_197), .B(n_176), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_232), .A2(n_238), .B(n_237), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_209), .B(n_178), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_197), .A2(n_178), .B(n_188), .C(n_180), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_199), .B(n_180), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_200), .A2(n_190), .B(n_184), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_198), .B(n_181), .Y(n_250) );
INVx5_ASAP7_75t_L g251 ( .A(n_203), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_203), .A2(n_184), .B1(n_181), .B2(n_190), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_199), .B(n_157), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_226), .B(n_131), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_228), .A2(n_187), .B(n_151), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_206), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
NOR3xp33_ASAP7_75t_L g259 ( .A(n_211), .B(n_157), .C(n_4), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_201), .B(n_157), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_202), .B(n_3), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_225), .A2(n_187), .B(n_151), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_207), .A2(n_151), .B(n_150), .C(n_147), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_207), .A2(n_224), .B(n_214), .C(n_219), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_151), .B(n_150), .C(n_147), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_205), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_239), .Y(n_269) );
OAI21x1_ASAP7_75t_SL g270 ( .A1(n_212), .A2(n_5), .B(n_6), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_231), .A2(n_5), .B(n_6), .C(n_8), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_225), .A2(n_151), .B(n_150), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_208), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_210), .A2(n_187), .B(n_151), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_241), .B(n_226), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_245), .A2(n_215), .B(n_213), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_275), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_263), .B(n_235), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_256), .A2(n_213), .B(n_210), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_251), .A2(n_234), .B1(n_233), .B2(n_230), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_222), .B(n_229), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_266), .A2(n_227), .B(n_223), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_256), .A2(n_234), .B(n_240), .Y(n_285) );
O2A1O1Ixp5_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_218), .B(n_221), .C(n_217), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_264), .A2(n_220), .B(n_147), .Y(n_287) );
O2A1O1Ixp5_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_236), .B(n_187), .C(n_150), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_242), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_266), .A2(n_147), .B(n_150), .C(n_12), .Y(n_290) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_243), .A2(n_150), .B(n_147), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_272), .A2(n_55), .B(n_97), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_244), .B(n_10), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_251), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_249), .A2(n_248), .B(n_247), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_276), .A2(n_54), .B(n_94), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_249), .A2(n_51), .B(n_92), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_251), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_252), .B(n_13), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_281), .A2(n_276), .B(n_270), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_296), .A2(n_267), .B(n_262), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_292), .B(n_262), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_277), .B(n_257), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_279), .B(n_257), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_279), .B(n_274), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_287), .A2(n_273), .B(n_269), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_290), .A2(n_265), .B(n_271), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_280), .B(n_274), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_260), .B(n_255), .Y(n_311) );
INVx6_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_300), .A2(n_258), .B1(n_259), .B2(n_246), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_268), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_282), .B(n_268), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_289), .B(n_268), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_295), .A2(n_262), .B1(n_271), .B2(n_253), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_290), .A2(n_261), .B(n_250), .Y(n_320) );
BUFx10_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_278), .A2(n_60), .B(n_14), .Y(n_322) );
BUFx2_ASAP7_75t_R g323 ( .A(n_294), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_299), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_307), .A2(n_297), .B(n_298), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_SL g327 ( .A1(n_319), .A2(n_283), .B(n_288), .C(n_291), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_315), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_316), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_304), .B(n_13), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_307), .A2(n_297), .B(n_293), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_321), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_311), .A2(n_293), .B(n_286), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_313), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_310), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
OA21x2_ASAP7_75t_L g347 ( .A1(n_313), .A2(n_15), .B(n_17), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_315), .B(n_18), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_301), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_19), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_312), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_302), .A2(n_20), .B(n_21), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_334), .B(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_334), .B(n_308), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_330), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_357), .B(n_308), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_357), .B(n_318), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_341), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_341), .B(n_318), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_335), .B(n_316), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_342), .B(n_303), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_329), .B(n_317), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_303), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_329), .B(n_321), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_337), .B(n_320), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_325), .B(n_314), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_332), .B(n_320), .C(n_317), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_329), .B(n_317), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_345), .B(n_320), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_325), .B(n_321), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_336), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_346), .B(n_321), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_350), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_348), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_350), .A2(n_320), .B1(n_317), .B2(n_303), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_345), .B(n_317), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_354), .B(n_323), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_354), .B(n_23), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_352), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_355), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_348), .A2(n_24), .B1(n_26), .B2(n_27), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_344), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_338), .B(n_31), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_338), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_338), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_349), .B(n_33), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_349), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_352), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_347), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_99), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_352), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_347), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_364), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_369), .B(n_352), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_363), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_377), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_361), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_398), .B(n_358), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_374), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_379), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_365), .B(n_352), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_365), .B(n_358), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_370), .B(n_408), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_376), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_370), .B(n_359), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_375), .B(n_359), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_359), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_386), .B(n_339), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_367), .B(n_339), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_401), .B(n_333), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_372), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_401), .B(n_333), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_360), .B(n_326), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_360), .B(n_326), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_362), .B(n_347), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_362), .B(n_347), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_395), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_385), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_366), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_368), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_393), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_410), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_411), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_391), .B(n_356), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_381), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_391), .B(n_356), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_375), .B(n_34), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_381), .B(n_36), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_389), .B(n_39), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_409), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_398), .B(n_327), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_390), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_395), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_373), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_375), .B(n_40), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_409), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_387), .B(n_41), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_387), .B(n_44), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_398), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_383), .B(n_45), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_371), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_387), .B(n_46), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_417), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_371), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_371), .B(n_48), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_402), .A2(n_57), .B1(n_61), .B2(n_62), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_418), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_414), .B(n_63), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_399), .B(n_65), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_399), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_378), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_403), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_399), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_379), .A2(n_67), .B1(n_69), .B2(n_71), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_396), .B(n_73), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_400), .B(n_75), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_403), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_419), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_384), .B(n_78), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_416), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_404), .B(n_79), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_412), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_404), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_420), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_433), .B(n_404), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_434), .B(n_404), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_426), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_476), .B(n_407), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_495), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_433), .B(n_407), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_430), .B(n_80), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_429), .B(n_81), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_441), .B(n_82), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_441), .B(n_83), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_473), .B(n_85), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_486), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_444), .B(n_86), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_465), .B(n_87), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_430), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_444), .B(n_88), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_447), .B(n_89), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_490), .B(n_90), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_432), .B(n_91), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_447), .B(n_475), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_432), .B(n_465), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_493), .B(n_474), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_501), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_474), .B(n_431), .Y(n_533) );
AND2x2_ASAP7_75t_SL g534 ( .A(n_492), .B(n_467), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_483), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_442), .B(n_456), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_427), .B(n_483), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_460), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_431), .B(n_453), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_436), .B(n_485), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_490), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_459), .B(n_461), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_501), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_443), .B(n_446), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_454), .B(n_449), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_437), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_485), .B(n_464), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_437), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_436), .B(n_481), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_462), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_462), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_464), .B(n_466), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_466), .B(n_500), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_435), .B(n_448), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_494), .B(n_449), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_463), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_457), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_448), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_445), .B(n_451), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_451), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_445), .B(n_468), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_436), .B(n_481), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_468), .B(n_503), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_435), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_422), .B(n_428), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_438), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_477), .B(n_479), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_438), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_479), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_457), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_421), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_421), .B(n_422), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_487), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_480), .B(n_478), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_423), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_480), .B(n_470), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_423), .B(n_424), .Y(n_578) );
INVx6_ASAP7_75t_L g579 ( .A(n_487), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_424), .B(n_425), .Y(n_580) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_487), .B(n_481), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_458), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_492), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_425), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_428), .B(n_455), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_505), .B(n_455), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_458), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_471), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_496), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_440), .B(n_489), .Y(n_590) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_467), .B(n_484), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_471), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_489), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_450), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_496), .B(n_450), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_472), .B(n_484), .Y(n_596) );
NOR2xp33_ASAP7_75t_SL g597 ( .A(n_467), .B(n_484), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_496), .B(n_452), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_452), .B(n_506), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_502), .B(n_499), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_504), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_530), .B(n_482), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_519), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_530), .B(n_482), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_583), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_507), .A2(n_499), .B1(n_497), .B2(n_502), .C(n_469), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_523), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
AOI221xp5_ASAP7_75t_SL g609 ( .A1(n_596), .A2(n_469), .B1(n_488), .B2(n_498), .C(n_472), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_590), .Y(n_610) );
AOI32xp33_ASAP7_75t_L g611 ( .A1(n_597), .A2(n_491), .A3(n_504), .B1(n_581), .B2(n_527), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_549), .B(n_491), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_574), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_539), .B(n_533), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_560), .B(n_491), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_522), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_504), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_567), .B(n_569), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_542), .B(n_536), .Y(n_620) );
NAND2x1_ASAP7_75t_L g621 ( .A(n_574), .B(n_579), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_588), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_510), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_536), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_588), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_519), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_546), .B(n_548), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_592), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_545), .B(n_538), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_592), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_556), .B(n_554), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_549), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_529), .B(n_547), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
NAND2x1_ASAP7_75t_L g635 ( .A(n_579), .B(n_549), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_560), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_594), .B(n_565), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_540), .B(n_599), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_594), .B(n_552), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_512), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
NOR2x1_ASAP7_75t_R g642 ( .A(n_596), .B(n_579), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_540), .B(n_562), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_550), .B(n_557), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_551), .B(n_559), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_540), .B(n_531), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_555), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_512), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_561), .B(n_572), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_572), .B(n_573), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_566), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_535), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_526), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_508), .B(n_585), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_526), .B(n_532), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_532), .B(n_543), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_578), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_578), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_541), .A2(n_513), .B1(n_537), .B2(n_591), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_595), .B(n_598), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_563), .B(n_509), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_580), .B(n_543), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_576), .B(n_584), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_580), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_558), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_575), .B(n_577), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_558), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_591), .B(n_570), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_571), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_568), .B(n_564), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_563), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_563), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_537), .B(n_589), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_534), .B(n_600), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_571), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_626), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_660), .A2(n_534), .B1(n_517), .B2(n_514), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_649), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_649), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_619), .Y(n_681) );
NAND2xp33_ASAP7_75t_L g682 ( .A(n_611), .B(n_525), .Y(n_682) );
AOI322xp5_ASAP7_75t_L g683 ( .A1(n_669), .A2(n_511), .A3(n_517), .B1(n_516), .B2(n_524), .C1(n_520), .C2(n_528), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_634), .B(n_593), .Y(n_684) );
NAND2xp33_ASAP7_75t_L g685 ( .A(n_614), .B(n_515), .Y(n_685) );
OAI32xp33_ASAP7_75t_L g686 ( .A1(n_607), .A2(n_528), .A3(n_589), .B1(n_521), .B2(n_518), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_606), .A2(n_517), .B1(n_518), .B2(n_601), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_607), .A2(n_582), .B1(n_587), .B2(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_619), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_636), .B(n_582), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_629), .B(n_587), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_653), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_606), .A2(n_609), .B1(n_675), .B2(n_620), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_621), .A2(n_614), .B(n_635), .C(n_609), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_645), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_612), .B(n_674), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_644), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_651), .B(n_655), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_676), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_644), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_608), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_624), .B(n_613), .Y(n_703) );
AOI32xp33_ASAP7_75t_L g704 ( .A1(n_632), .A2(n_673), .A3(n_674), .B1(n_646), .B2(n_671), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_664), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_647), .B(n_627), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_650), .B(n_659), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_664), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_662), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_652), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_603), .A2(n_612), .B(n_676), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_603), .A2(n_602), .B(n_604), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_639), .Y(n_713) );
NOR2xp67_ASAP7_75t_L g714 ( .A(n_672), .B(n_662), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g715 ( .A1(n_632), .A2(n_673), .B(n_627), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_617), .B(n_623), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_643), .B(n_638), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_639), .A2(n_605), .B(n_665), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_658), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_610), .B(n_631), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_637), .B(n_663), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_694), .A2(n_616), .B1(n_667), .B2(n_641), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_714), .A2(n_633), .B1(n_661), .B2(n_615), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_678), .A2(n_642), .B(n_618), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_697), .B(n_654), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_697), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_713), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_695), .B(n_657), .C(n_656), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_698), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_701), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_677), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_705), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_708), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_709), .B(n_648), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_682), .A2(n_656), .B(n_657), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_690), .Y(n_736) );
OAI21xp5_ASAP7_75t_SL g737 ( .A1(n_704), .A2(n_640), .B(n_625), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_699), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_696), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_712), .B(n_622), .Y(n_740) );
NOR4xp25_ASAP7_75t_L g741 ( .A(n_693), .B(n_628), .C(n_630), .D(n_666), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_715), .B(n_668), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_679), .B(n_670), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_707), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_685), .A2(n_711), .B1(n_686), .B2(n_706), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_724), .A2(n_711), .B(n_718), .Y(n_746) );
AOI221x1_ASAP7_75t_L g747 ( .A1(n_728), .A2(n_680), .B1(n_712), .B2(n_702), .C(n_681), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_745), .B(n_687), .C(n_719), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_722), .B(n_689), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_728), .A2(n_703), .B(n_716), .C(n_710), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g751 ( .A1(n_745), .A2(n_683), .B(n_688), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_L g752 ( .A1(n_737), .A2(n_742), .B(n_741), .C(n_726), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_738), .B(n_720), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_723), .A2(n_692), .B(n_684), .Y(n_754) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_726), .B(n_700), .Y(n_755) );
NOR2xp67_ASAP7_75t_L g756 ( .A(n_735), .B(n_721), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_722), .A2(n_691), .B1(n_717), .B2(n_727), .C(n_744), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_725), .A2(n_731), .B1(n_740), .B2(n_730), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_749), .B(n_729), .Y(n_759) );
NOR3x1_ASAP7_75t_L g760 ( .A(n_751), .B(n_732), .C(n_733), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_748), .B(n_736), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_757), .B(n_739), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_754), .B(n_731), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_756), .B(n_743), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_763), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_761), .B(n_752), .Y(n_766) );
NOR3x1_ASAP7_75t_L g767 ( .A(n_764), .B(n_758), .C(n_747), .Y(n_767) );
XNOR2x1_ASAP7_75t_L g768 ( .A(n_759), .B(n_755), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_765), .B(n_746), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_766), .B(n_760), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_768), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_771), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_769), .B(n_762), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_772), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_773), .Y(n_775) );
NOR2x1p5_ASAP7_75t_L g776 ( .A(n_774), .B(n_775), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_776), .B(n_770), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_777), .B(n_770), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_779), .B(n_770), .Y(n_780) );
OAI21x1_ASAP7_75t_L g781 ( .A1(n_780), .A2(n_750), .B(n_753), .Y(n_781) );
AO21x2_ASAP7_75t_L g782 ( .A1(n_781), .A2(n_767), .B(n_734), .Y(n_782) );
endmodule