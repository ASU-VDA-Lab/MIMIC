module fake_ariane_313_n_7206 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_638, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_7206);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_7206;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_6664;
wire n_1018;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_6539;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_863;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5452;
wire n_5391;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_1389;
wire n_3172;
wire n_4033;
wire n_2659;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_974;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_7007;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_6665;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_1568;
wire n_2919;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_6382;
wire n_670;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_6615;
wire n_6192;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_1163;
wire n_4970;
wire n_3054;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_5858;
wire n_5985;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_688;
wire n_7176;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_1104;
wire n_986;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_4856;
wire n_2618;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_6508;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_1044;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_7076;
wire n_6344;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_3715;
wire n_1593;
wire n_2626;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_6706;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_6551;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_6757;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_6905;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_4230;
wire n_3040;
wire n_6899;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_1261;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_3632;
wire n_2522;
wire n_1344;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_840;
wire n_6575;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_3445;
wire n_2105;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_5844;
wire n_6298;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_774;
wire n_5548;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_1581;
wire n_946;
wire n_757;
wire n_5355;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_7160;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_5360;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_6607;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_6552;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_3728;
wire n_2722;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_4593;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_3429;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_3758;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_6947;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_2855;
wire n_794;
wire n_2848;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_5981;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_6623;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_6390;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_5735;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_6865;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_4818;
wire n_7020;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_5832;
wire n_6254;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_6987;
wire n_877;
wire n_3995;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3568;
wire n_3216;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_982;
wire n_915;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_6139;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_2751;
wire n_3113;
wire n_1622;
wire n_4183;
wire n_1968;
wire n_918;
wire n_5645;
wire n_5020;
wire n_673;
wire n_6455;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_692;
wire n_4457;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7188;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_3278;
wire n_2375;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_6493;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_5887;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3775;
wire n_3148;
wire n_5682;
wire n_684;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_6590;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_6885;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_1752;
wire n_2361;
wire n_3030;
wire n_4538;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_5823;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_6299;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1187;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_672;
wire n_4968;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_5290;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_6394;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_6504;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_6868;
wire n_5131;
wire n_6813;
wire n_5546;
wire n_6294;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_6713;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_2220;
wire n_7044;
wire n_6108;
wire n_6100;
wire n_6800;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_7066;
wire n_5496;
wire n_3104;
wire n_7174;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_5132;
wire n_3498;
wire n_1173;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_6432;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_4293;
wire n_2937;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_5681;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_6591;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_3426;
wire n_2660;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_5420;
wire n_6497;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_7073;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_1804;
wire n_6519;
wire n_4671;
wire n_5989;
wire n_5571;
wire n_4766;
wire n_2272;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_6490;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_7019;
wire n_682;
wire n_5315;
wire n_3708;
wire n_2633;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_979;
wire n_3976;
wire n_3381;
wire n_2546;
wire n_2813;
wire n_897;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_3955;
wire n_1659;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_6971;
wire n_3336;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_5912;
wire n_801;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7107;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_2475;
wire n_1185;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_4412;
wire n_2845;
wire n_2036;
wire n_6923;
wire n_843;
wire n_3358;
wire n_6704;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_5005;
wire n_6126;
wire n_1549;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_5474;
wire n_2767;
wire n_7009;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_1767;
wire n_1040;
wire n_4138;
wire n_3131;
wire n_7083;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_2154;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_1772;
wire n_6879;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_7082;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_4406;
wire n_2180;
wire n_4271;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_6955;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_6832;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_3387;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_977;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_6499;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_6982;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_6400;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_7154;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_7068;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_4549;
wire n_1073;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_6675;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_7056;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_6988;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_804;
wire n_6649;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_6431;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_5659;
wire n_6859;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_6410;
wire n_6473;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_836;
wire n_6975;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_4725;
wire n_2757;
wire n_2312;
wire n_7203;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_6772;
wire n_7088;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_6617;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_6742;
wire n_1467;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_3988;
wire n_2599;
wire n_5022;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3996;
wire n_3761;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_777;
wire n_7095;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_6465;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_6940;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_657;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_1466;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_6825;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_876;
wire n_5872;
wire n_6692;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_3543;
wire n_1324;
wire n_2945;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_6322;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_7089;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_5104;
wire n_6961;
wire n_6792;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_907;
wire n_7118;
wire n_6152;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_6282;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_6737;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_7038;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_1093;
wire n_6518;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_4168;
wire n_1369;
wire n_7036;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_7099;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_3772;
wire n_2891;
wire n_7026;
wire n_4335;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_6436;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_3935;
wire n_2654;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_90),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_475),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_577),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_274),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_523),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_607),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_99),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_384),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_611),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_630),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_492),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_521),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_458),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_399),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_644),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_419),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_202),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_22),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_31),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_126),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_552),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_534),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_546),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_609),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_212),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_359),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_362),
.Y(n_678)
);

CKINVDCx14_ASAP7_75t_R g679 ( 
.A(n_460),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_182),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_30),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_81),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_135),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_103),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_65),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_450),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_485),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_557),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_79),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_548),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_62),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_155),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_257),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_542),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_522),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_378),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_166),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_534),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_552),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_472),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_418),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_123),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_108),
.Y(n_703)
);

BUFx5_ASAP7_75t_L g704 ( 
.A(n_33),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_48),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_362),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_409),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_400),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_169),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_372),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_235),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_316),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_173),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_402),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_29),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_636),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_127),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_444),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_1),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_598),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_191),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_137),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_622),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_185),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_117),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_10),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_536),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_293),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_548),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_572),
.Y(n_731)
);

BUFx8_ASAP7_75t_SL g732 ( 
.A(n_220),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_373),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_257),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_20),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_330),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_382),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_210),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_196),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_303),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_648),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_616),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_505),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_463),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_475),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_537),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_122),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_388),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_392),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_351),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_82),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_274),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_604),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_92),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_95),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_616),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_321),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_296),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_525),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_68),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_575),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_219),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_556),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_414),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_609),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_119),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_80),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_161),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_238),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_9),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_209),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_629),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_451),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_420),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_379),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_587),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_554),
.Y(n_777)
);

CKINVDCx14_ASAP7_75t_R g778 ( 
.A(n_588),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_409),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_148),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_607),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_111),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_389),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_364),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_244),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_615),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_351),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_593),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_47),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_642),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_154),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_442),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_641),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_468),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_93),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_157),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_1),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_102),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_536),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_197),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_162),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_383),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_529),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_190),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_87),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_264),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_384),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_126),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_355),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_193),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_297),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_540),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_647),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_8),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_206),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_216),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_329),
.Y(n_817)
);

BUFx5_ASAP7_75t_L g818 ( 
.A(n_322),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_256),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_281),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_647),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_377),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_258),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_405),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_14),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_374),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_237),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_436),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_372),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_509),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_83),
.Y(n_831)
);

CKINVDCx14_ASAP7_75t_R g832 ( 
.A(n_603),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_8),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_171),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_79),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_278),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_342),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_270),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_438),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_157),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_147),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_18),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_149),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_43),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_92),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_99),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_394),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_136),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_199),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_34),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_151),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_195),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_187),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_149),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_318),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_280),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_566),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_397),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_650),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_645),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_556),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_541),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_20),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_321),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_443),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_77),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_192),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_265),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_287),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_578),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_509),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_482),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_453),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_15),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_595),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_27),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_56),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_43),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_417),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_617),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_265),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_253),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_517),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_25),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_11),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_235),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_593),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_108),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_605),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_356),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_102),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_110),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_579),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_452),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_571),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_170),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_129),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_350),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_242),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_599),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_114),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_78),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_357),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_17),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_527),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_315),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_638),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_640),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_495),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_327),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_96),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_538),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_505),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_645),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_454),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_258),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_200),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_560),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_233),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_443),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_459),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_175),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_270),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_511),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_512),
.Y(n_925)
);

CKINVDCx14_ASAP7_75t_R g926 ( 
.A(n_206),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_639),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_617),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_573),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_560),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_476),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_597),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_459),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_22),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_353),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_363),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_42),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_10),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_50),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_12),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_591),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_308),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_280),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_120),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_547),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_59),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_416),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_318),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_371),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_64),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_426),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_577),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_221),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_175),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_634),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_290),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_367),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_266),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_54),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_196),
.Y(n_960)
);

CKINVDCx16_ASAP7_75t_R g961 ( 
.A(n_341),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_324),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_448),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_131),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_325),
.Y(n_965)
);

CKINVDCx16_ASAP7_75t_R g966 ( 
.A(n_342),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_613),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_319),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_111),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_425),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_231),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_164),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_462),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_85),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_650),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_353),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_177),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_24),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_214),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_323),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_394),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_393),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_500),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_421),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_218),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_544),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_589),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_621),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_502),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_340),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_435),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_596),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_636),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_603),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_314),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_267),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_501),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_208),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_426),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_628),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_510),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_578),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_309),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_493),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_181),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_204),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_344),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_392),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_583),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_515),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_201),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_324),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_565),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_153),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_366),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_234),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_345),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_620),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_403),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_629),
.Y(n_1020)
);

BUFx10_ASAP7_75t_L g1021 ( 
.A(n_402),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_335),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_141),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_133),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_508),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_14),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_227),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_24),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_125),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_619),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_141),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_241),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_295),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_65),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_307),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_53),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_88),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_460),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_388),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_562),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_553),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_13),
.Y(n_1042)
);

CKINVDCx16_ASAP7_75t_R g1043 ( 
.A(n_520),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_457),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_364),
.Y(n_1045)
);

CKINVDCx14_ASAP7_75t_R g1046 ( 
.A(n_176),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_513),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_40),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_10),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_375),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_172),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_314),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_424),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_332),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_228),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_160),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_341),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_611),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_602),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_387),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_516),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_557),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_375),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_635),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_430),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_253),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_133),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_494),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_278),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_312),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_349),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_328),
.Y(n_1072)
);

BUFx10_ASAP7_75t_L g1073 ( 
.A(n_207),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_12),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_604),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_125),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_29),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_53),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_397),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_618),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_101),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_169),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_98),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_483),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_5),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_208),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_434),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_531),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_531),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_606),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_491),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_412),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_249),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_199),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_223),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_408),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_581),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_551),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_6),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_22),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_21),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_138),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_643),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_89),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_606),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_205),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_451),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_563),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_73),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_262),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_541),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_576),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_50),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_334),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_519),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_217),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_621),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_38),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_150),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_146),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_523),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_28),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_203),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_286),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_377),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_33),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_246),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_374),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_461),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_302),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_553),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_46),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_0),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_469),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_498),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_332),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_456),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_511),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_27),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_532),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_156),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_571),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_620),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_90),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_210),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_313),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_241),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_453),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_292),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_171),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_244),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_112),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_46),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_640),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_279),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_385),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_352),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_194),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_434),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_575),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_288),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_586),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_608),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_130),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_277),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_14),
.Y(n_1166)
);

CKINVDCx16_ASAP7_75t_R g1167 ( 
.A(n_601),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_649),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_600),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_204),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_201),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_537),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_468),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_573),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_494),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_479),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_211),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_623),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_608),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_508),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_74),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_477),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_348),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_306),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_45),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_527),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_61),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_31),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_41),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_309),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_181),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_681),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_679),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_679),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_681),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_778),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_778),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_832),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_832),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_681),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1085),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1085),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_926),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_926),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1046),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1085),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1189),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1189),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_1189),
.B(n_0),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_706),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_732),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1046),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_732),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_711),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1189),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_704),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1189),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_704),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_704),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1166),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_711),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_654),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_708),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1166),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_708),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_708),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_654),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_776),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1191),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_706),
.B(n_0),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_730),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_677),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_704),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_730),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_776),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_730),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_762),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_781),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_704),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_781),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_909),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_762),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_762),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_786),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_786),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_786),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_796),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_796),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_757),
.B(n_1),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_796),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_909),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_801),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_801),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_961),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_961),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_801),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_892),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_892),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_966),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_739),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_966),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_892),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1037),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_907),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1037),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_907),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1191),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1043),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_907),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_945),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1043),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_670),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1076),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_945),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_945),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_995),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1076),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1095),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_995),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_995),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_704),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1095),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_757),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_670),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1167),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1010),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1010),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_704),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1010),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_1100),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1067),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_838),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1067),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1067),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1098),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_739),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1098),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1167),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1098),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1157),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

BUFx5_ASAP7_75t_L g1302 ( 
.A(n_1157),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_838),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_704),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1179),
.Y(n_1305)
);

CKINVDCx16_ASAP7_75t_R g1306 ( 
.A(n_1179),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_652),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_677),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1100),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_782),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_707),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_656),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_704),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_704),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_657),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_704),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_658),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_659),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_661),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_669),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_669),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_669),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1000),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_662),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_735),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_664),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_818),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_735),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_818),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_735),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_666),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_653),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_782),
.B(n_2),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_653),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_653),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_667),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_668),
.Y(n_1337)
);

INVxp33_ASAP7_75t_SL g1338 ( 
.A(n_1000),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1100),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_671),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_722),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_722),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_722),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_756),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_756),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_756),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_672),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_860),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_674),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_860),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_675),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_860),
.Y(n_1352)
);

CKINVDCx16_ASAP7_75t_R g1353 ( 
.A(n_696),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_818),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1031),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_864),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1031),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_864),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_676),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_680),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_707),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_686),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_818),
.Y(n_1363)
);

BUFx5_ASAP7_75t_L g1364 ( 
.A(n_874),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_682),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_684),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_687),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_688),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_690),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_691),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_692),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_694),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1072),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_818),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_697),
.Y(n_1375)
);

BUFx5_ASAP7_75t_L g1376 ( 
.A(n_874),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_731),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1072),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_702),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_709),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_710),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1133),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_896),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_731),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_942),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_716),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_963),
.B(n_2),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_818),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_963),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_896),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_963),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_717),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_719),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1133),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_967),
.B(n_2),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_721),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_967),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1064),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_724),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_818),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_967),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_994),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_994),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_994),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1006),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_726),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1006),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1006),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_772),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_728),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1036),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_818),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_772),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1036),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1036),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_733),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_734),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1054),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_736),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1054),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1054),
.B(n_3),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1100),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1100),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1100),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1064),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_818),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1100),
.Y(n_1427)
);

BUFx10_ASAP7_75t_L g1428 ( 
.A(n_686),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_737),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_738),
.Y(n_1430)
);

BUFx2_ASAP7_75t_SL g1431 ( 
.A(n_696),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_904),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_715),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_904),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_741),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_815),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_700),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_660),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_696),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_700),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_742),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_815),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_818),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_744),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_746),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_818),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_686),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_700),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_792),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_747),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_686),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_792),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_816),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_750),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_686),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_792),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_753),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_754),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_822),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_759),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_760),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_761),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_822),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_822),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_857),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_686),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_696),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_857),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_857),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_686),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_765),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_766),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_660),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_871),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_871),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_871),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_767),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_873),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_873),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_873),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_768),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1101),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_771),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_893),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_893),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_893),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_720),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_816),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_931),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_821),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_931),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_812),
.B(n_3),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_775),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_779),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_931),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_780),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_946),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_785),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_713),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_946),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_946),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_965),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_821),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_787),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_965),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_965),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_977),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_788),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_977),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_977),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1004),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_713),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_826),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_791),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_812),
.B(n_3),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_793),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_794),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_713),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_795),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1004),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_798),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1004),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_826),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_802),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_932),
.B(n_4),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_663),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1032),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_803),
.Y(n_1528)
);

XOR2xp5_ASAP7_75t_L g1529 ( 
.A(n_1101),
.B(n_4),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_727),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_805),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1032),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_806),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_770),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1032),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_713),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_851),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1051),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1051),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_851),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_808),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_663),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_932),
.B(n_1027),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_865),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_713),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_811),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1051),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_817),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1057),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_820),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1057),
.Y(n_1551)
);

BUFx5_ASAP7_75t_L g1552 ( 
.A(n_665),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_865),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1057),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1079),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1079),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1079),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1088),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_797),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1088),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1088),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_823),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_866),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1132),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_824),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1132),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_827),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_828),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1132),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1168),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_829),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_713),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1168),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_713),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1168),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_830),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1176),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_831),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1176),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1176),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_718),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_834),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_718),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_665),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_718),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_696),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_835),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_837),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_683),
.B(n_4),
.Y(n_1589)
);

INVxp33_ASAP7_75t_L g1590 ( 
.A(n_683),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_839),
.Y(n_1591)
);

NOR2xp67_ASAP7_75t_L g1592 ( 
.A(n_1027),
.B(n_5),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_718),
.Y(n_1593)
);

NOR2xp67_ASAP7_75t_L g1594 ( 
.A(n_1091),
.B(n_5),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_718),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_843),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_689),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_689),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_866),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_845),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_693),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_894),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_847),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_849),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_718),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_693),
.Y(n_1606)
);

CKINVDCx16_ASAP7_75t_R g1607 ( 
.A(n_748),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_695),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_695),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_698),
.Y(n_1610)
);

CKINVDCx14_ASAP7_75t_R g1611 ( 
.A(n_748),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_850),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_698),
.B(n_6),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_699),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_748),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_699),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_894),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_701),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_814),
.Y(n_1619)
);

BUFx2_ASAP7_75t_SL g1620 ( 
.A(n_748),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_852),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_853),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_701),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_703),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_703),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_718),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_705),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_854),
.Y(n_1628)
);

XOR2x2_ASAP7_75t_L g1629 ( 
.A(n_673),
.B(n_6),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_705),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_714),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_902),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_855),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_819),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_856),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_714),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_723),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_723),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_859),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_861),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_725),
.B(n_7),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_862),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_867),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_819),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_819),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_725),
.Y(n_1646)
);

INVxp33_ASAP7_75t_L g1647 ( 
.A(n_729),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_870),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_729),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_825),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_872),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_877),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_740),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_740),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_743),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_743),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_819),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_902),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_879),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1229),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1207),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1208),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1222),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1227),
.Y(n_1664)
);

CKINVDCx16_ASAP7_75t_R g1665 ( 
.A(n_1203),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1213),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1215),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1217),
.Y(n_1668)
);

CKINVDCx16_ASAP7_75t_R g1669 ( 
.A(n_1353),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1611),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1213),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1232),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1193),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1485),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1290),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1308),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1311),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1332),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1193),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1194),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1194),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1334),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1196),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1455),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1335),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1341),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1342),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1196),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1197),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1343),
.Y(n_1690)
);

CKINVDCx20_ASAP7_75t_R g1691 ( 
.A(n_1361),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1455),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1344),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1345),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1214),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1346),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1197),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1198),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1348),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1350),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1198),
.Y(n_1701)
);

CKINVDCx16_ASAP7_75t_R g1702 ( 
.A(n_1439),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1352),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1356),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1214),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1358),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1339),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1199),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1199),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1272),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1204),
.Y(n_1711)
);

CKINVDCx16_ASAP7_75t_R g1712 ( 
.A(n_1586),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1233),
.Y(n_1713)
);

INVxp33_ASAP7_75t_SL g1714 ( 
.A(n_1431),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1221),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1385),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1204),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1466),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1284),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1205),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1377),
.Y(n_1721)
);

BUFx2_ASAP7_75t_SL g1722 ( 
.A(n_1212),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1389),
.Y(n_1723)
);

INVxp67_ASAP7_75t_SL g1724 ( 
.A(n_1233),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1205),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1391),
.Y(n_1726)
);

CKINVDCx16_ASAP7_75t_R g1727 ( 
.A(n_1607),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1397),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1401),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1382),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1329),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1402),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1403),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1404),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1466),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1405),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1644),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1306),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1394),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1407),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1384),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1307),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1436),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1307),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1408),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1221),
.Y(n_1746)
);

INVxp33_ASAP7_75t_L g1747 ( 
.A(n_1433),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1411),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1312),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1431),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1228),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_1442),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1414),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1415),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_1488),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1418),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1420),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1650),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1223),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1650),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1409),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1225),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1226),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1312),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1329),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1315),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1620),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1354),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1315),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1231),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1234),
.Y(n_1771)
);

CKINVDCx16_ASAP7_75t_R g1772 ( 
.A(n_1620),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1490),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1236),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1237),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1242),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1243),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1244),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1245),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1487),
.Y(n_1780)
);

CKINVDCx20_ASAP7_75t_R g1781 ( 
.A(n_1513),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1523),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1317),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1246),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1247),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1248),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1250),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1228),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_1537),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1317),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1252),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1540),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1553),
.Y(n_1793)
);

CKINVDCx16_ASAP7_75t_R g1794 ( 
.A(n_1211),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1253),
.Y(n_1795)
);

CKINVDCx14_ASAP7_75t_R g1796 ( 
.A(n_1235),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1318),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1256),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1235),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1354),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1257),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1258),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1262),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1264),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1318),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1530),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1413),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1266),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1374),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1309),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1599),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1269),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1270),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1319),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1274),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1275),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1276),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1319),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1545),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1374),
.Y(n_1820)
);

CKINVDCx14_ASAP7_75t_R g1821 ( 
.A(n_1238),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1279),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1238),
.Y(n_1823)
);

INVxp67_ASAP7_75t_SL g1824 ( 
.A(n_1400),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1240),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1280),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1324),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1240),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1286),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1287),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1289),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1324),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1602),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1291),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1293),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1545),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1400),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1326),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1572),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1617),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1294),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1295),
.Y(n_1842)
);

CKINVDCx20_ASAP7_75t_R g1843 ( 
.A(n_1632),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1241),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1297),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1658),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1572),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1412),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1299),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1300),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1574),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1301),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1326),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1331),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1331),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1192),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1195),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1201),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1574),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1202),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1206),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1584),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1597),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1598),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1534),
.Y(n_1865)
);

INVxp33_ASAP7_75t_SL g1866 ( 
.A(n_1336),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1453),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1601),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1559),
.Y(n_1869)
);

INVxp33_ASAP7_75t_SL g1870 ( 
.A(n_1336),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1337),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1503),
.Y(n_1872)
);

INVx4_ASAP7_75t_R g1873 ( 
.A(n_1467),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1241),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1606),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1608),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1609),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1251),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1251),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1610),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1614),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1619),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1337),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1616),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1309),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1618),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1340),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1623),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1340),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1624),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1451),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1625),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1544),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1347),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1627),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1630),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1347),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1631),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1309),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1636),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1349),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1349),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1451),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1637),
.Y(n_1904)
);

CKINVDCx20_ASAP7_75t_R g1905 ( 
.A(n_1563),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1482),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1638),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1646),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1351),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1482),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1254),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1649),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1383),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1654),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1390),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1655),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1656),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1432),
.Y(n_1918)
);

INVxp67_ASAP7_75t_SL g1919 ( 
.A(n_1499),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1434),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1351),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1254),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1200),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1200),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1359),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1302),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1255),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1359),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1302),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_1255),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1302),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1302),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1360),
.Y(n_1933)
);

INVxp67_ASAP7_75t_L g1934 ( 
.A(n_1260),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1302),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1302),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1302),
.Y(n_1937)
);

CKINVDCx16_ASAP7_75t_R g1938 ( 
.A(n_1467),
.Y(n_1938)
);

INVxp33_ASAP7_75t_SL g1939 ( 
.A(n_1360),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1302),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1581),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1365),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1259),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1260),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1364),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1581),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1365),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1259),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1296),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1364),
.Y(n_1950)
);

CKINVDCx16_ASAP7_75t_R g1951 ( 
.A(n_1615),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1366),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1261),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_1261),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1263),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1364),
.Y(n_1956)
);

INVxp67_ASAP7_75t_SL g1957 ( 
.A(n_1499),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1364),
.Y(n_1958)
);

INVxp33_ASAP7_75t_L g1959 ( 
.A(n_1303),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1364),
.Y(n_1960)
);

CKINVDCx20_ASAP7_75t_R g1961 ( 
.A(n_1263),
.Y(n_1961)
);

CKINVDCx16_ASAP7_75t_R g1962 ( 
.A(n_1615),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1364),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1364),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1366),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1364),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1583),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1265),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1367),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1265),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1268),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1367),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1376),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1268),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1376),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1368),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1376),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1296),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1271),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1368),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1369),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1271),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1376),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1369),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1229),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1376),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1310),
.Y(n_1987)
);

CKINVDCx16_ASAP7_75t_R g1988 ( 
.A(n_1310),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1376),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1376),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1398),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1376),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1428),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1320),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1321),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1322),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1512),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1398),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1370),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1325),
.Y(n_2000)
);

INVx1_ASAP7_75t_SL g2001 ( 
.A(n_1273),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1583),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1595),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1328),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1330),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1273),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1437),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1440),
.Y(n_2008)
);

CKINVDCx16_ASAP7_75t_R g2009 ( 
.A(n_1425),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1448),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1449),
.Y(n_2011)
);

CKINVDCx16_ASAP7_75t_R g2012 ( 
.A(n_1425),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1370),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1452),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1371),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1456),
.Y(n_2016)
);

INVxp67_ASAP7_75t_SL g2017 ( 
.A(n_1512),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_1277),
.Y(n_2018)
);

CKINVDCx14_ASAP7_75t_R g2019 ( 
.A(n_1277),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1459),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1463),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1464),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1371),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1465),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1468),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1469),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1372),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1474),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1536),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1536),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1475),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1476),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1595),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1372),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1605),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1478),
.Y(n_2036)
);

INVxp33_ASAP7_75t_L g2037 ( 
.A(n_1373),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1479),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1375),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1923),
.B(n_1589),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1675),
.B(n_1552),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1684),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1710),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1924),
.B(n_1589),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1707),
.B(n_1552),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1684),
.Y(n_2046)
);

OAI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1750),
.A2(n_1249),
.B1(n_1338),
.B2(n_1590),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1692),
.Y(n_2048)
);

BUFx8_ASAP7_75t_L g2049 ( 
.A(n_1695),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1731),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1731),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1674),
.B(n_1589),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1692),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1718),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1718),
.Y(n_2055)
);

OA21x2_ASAP7_75t_L g2056 ( 
.A1(n_1945),
.A2(n_1313),
.B(n_1304),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1739),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1767),
.B(n_1230),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1735),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1735),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1768),
.Y(n_2061)
);

OA21x2_ASAP7_75t_L g2062 ( 
.A1(n_1950),
.A2(n_1316),
.B(n_1314),
.Y(n_2062)
);

BUFx8_ASAP7_75t_L g2063 ( 
.A(n_1705),
.Y(n_2063)
);

BUFx8_ASAP7_75t_L g2064 ( 
.A(n_1715),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1819),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1819),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_1768),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1737),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1926),
.A2(n_1218),
.B(n_1216),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1759),
.B(n_1249),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1810),
.B(n_1552),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1836),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1678),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1682),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1685),
.Y(n_2075)
);

AND2x6_ASAP7_75t_L g2076 ( 
.A(n_1929),
.B(n_1333),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1719),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1686),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1687),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1836),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1839),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1714),
.B(n_1375),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1762),
.B(n_1613),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1810),
.B(n_1714),
.Y(n_2084)
);

INVx5_ASAP7_75t_L g2085 ( 
.A(n_1660),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1839),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1690),
.Y(n_2087)
);

OAI22x1_ASAP7_75t_L g2088 ( 
.A1(n_1739),
.A2(n_1529),
.B1(n_1629),
.B2(n_1220),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1763),
.B(n_1613),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1938),
.B(n_1379),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1693),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1794),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1770),
.B(n_1641),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1847),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1847),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1694),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1772),
.A2(n_1338),
.B1(n_1543),
.B2(n_1282),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1851),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1851),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1696),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1660),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1931),
.A2(n_1218),
.B(n_1216),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1859),
.Y(n_2103)
);

INVxp33_ASAP7_75t_SL g2104 ( 
.A(n_1742),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1699),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1765),
.B(n_1552),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1730),
.B(n_1647),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1771),
.B(n_1641),
.Y(n_2108)
);

INVx4_ASAP7_75t_L g2109 ( 
.A(n_1885),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1700),
.Y(n_2110)
);

CKINVDCx6p67_ASAP7_75t_R g2111 ( 
.A(n_1738),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1859),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1660),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1703),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1951),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1941),
.Y(n_2116)
);

OA21x2_ASAP7_75t_L g2117 ( 
.A1(n_1956),
.A2(n_1239),
.B(n_1219),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1670),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1941),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1962),
.A2(n_1282),
.B1(n_1285),
.B2(n_1278),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1660),
.Y(n_2121)
);

INVx5_ASAP7_75t_L g2122 ( 
.A(n_1985),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1946),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1946),
.Y(n_2124)
);

NAND2xp33_ASAP7_75t_L g2125 ( 
.A(n_1932),
.B(n_1552),
.Y(n_2125)
);

BUFx12f_ASAP7_75t_L g2126 ( 
.A(n_1666),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1967),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1985),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_1758),
.B(n_1379),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1670),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1967),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2002),
.Y(n_2132)
);

INVx5_ASAP7_75t_L g2133 ( 
.A(n_1985),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_1985),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1760),
.A2(n_1806),
.B1(n_1865),
.B2(n_1780),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2002),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1869),
.A2(n_1285),
.B1(n_1298),
.B2(n_1278),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_1935),
.A2(n_1239),
.B(n_1219),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_1882),
.B(n_1380),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2003),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2003),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_SL g2142 ( 
.A1(n_1906),
.A2(n_1529),
.B1(n_937),
.B2(n_952),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2033),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1774),
.B(n_1653),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1747),
.B(n_1380),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_2033),
.Y(n_2146)
);

INVxp67_ASAP7_75t_L g2147 ( 
.A(n_1761),
.Y(n_2147)
);

CKINVDCx20_ASAP7_75t_R g2148 ( 
.A(n_1663),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2035),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2035),
.Y(n_2150)
);

OA21x2_ASAP7_75t_L g2151 ( 
.A1(n_1958),
.A2(n_1288),
.B(n_1281),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_1775),
.B(n_1438),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1800),
.B(n_1552),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1862),
.B(n_1473),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1661),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1742),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1936),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_SL g2158 ( 
.A1(n_1988),
.A2(n_937),
.B1(n_952),
.B2(n_906),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1662),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1960),
.Y(n_2160)
);

OA21x2_ASAP7_75t_L g2161 ( 
.A1(n_1963),
.A2(n_1288),
.B(n_1281),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1964),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1937),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1940),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1885),
.Y(n_2165)
);

CKINVDCx11_ASAP7_75t_R g2166 ( 
.A(n_1911),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_1776),
.B(n_1526),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1667),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1866),
.A2(n_1305),
.B1(n_1298),
.B2(n_1381),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1809),
.B(n_1552),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1899),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1777),
.B(n_1542),
.Y(n_2172)
);

CKINVDCx8_ASAP7_75t_R g2173 ( 
.A(n_1722),
.Y(n_2173)
);

INVx6_ASAP7_75t_L g2174 ( 
.A(n_1993),
.Y(n_2174)
);

INVx4_ASAP7_75t_L g2175 ( 
.A(n_1993),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1966),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1668),
.Y(n_2177)
);

CKINVDCx11_ASAP7_75t_R g2178 ( 
.A(n_1911),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1994),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1778),
.B(n_1387),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1744),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1820),
.B(n_1552),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_2009),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1824),
.B(n_1381),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1673),
.B(n_1679),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1973),
.Y(n_2186)
);

OA21x2_ASAP7_75t_L g2187 ( 
.A1(n_1975),
.A2(n_1363),
.B(n_1327),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1977),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1866),
.B(n_1386),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1983),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1986),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_2012),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1989),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_1990),
.A2(n_1363),
.B(n_1327),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1744),
.Y(n_2195)
);

OA21x2_ASAP7_75t_L g2196 ( 
.A1(n_1992),
.A2(n_1426),
.B(n_1388),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2007),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1704),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1807),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1706),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_1779),
.B(n_1395),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1749),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1995),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1837),
.B(n_1386),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1749),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1848),
.B(n_1392),
.Y(n_2206)
);

BUFx6f_ASAP7_75t_L g2207 ( 
.A(n_1996),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_2000),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_1784),
.B(n_1421),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2008),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_2004),
.Y(n_2211)
);

INVx5_ASAP7_75t_L g2212 ( 
.A(n_1665),
.Y(n_2212)
);

CKINVDCx6p67_ASAP7_75t_R g2213 ( 
.A(n_1669),
.Y(n_2213)
);

BUFx8_ASAP7_75t_SL g2214 ( 
.A(n_1663),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1797),
.Y(n_2215)
);

INVx3_ASAP7_75t_L g2216 ( 
.A(n_2005),
.Y(n_2216)
);

NOR2x1_ASAP7_75t_L g2217 ( 
.A(n_1918),
.B(n_1220),
.Y(n_2217)
);

OA21x2_ASAP7_75t_L g2218 ( 
.A1(n_2010),
.A2(n_1426),
.B(n_1388),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1891),
.B(n_1392),
.Y(n_2219)
);

OA21x2_ASAP7_75t_L g2220 ( 
.A1(n_2011),
.A2(n_1446),
.B(n_1443),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2014),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_1785),
.B(n_1786),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_2016),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_2020),
.Y(n_2224)
);

OAI21x1_ASAP7_75t_L g2225 ( 
.A1(n_1856),
.A2(n_1446),
.B(n_1443),
.Y(n_2225)
);

OA21x2_ASAP7_75t_L g2226 ( 
.A1(n_2021),
.A2(n_1423),
.B(n_1422),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_2022),
.Y(n_2227)
);

OA21x2_ASAP7_75t_L g2228 ( 
.A1(n_2024),
.A2(n_1427),
.B(n_1424),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_2025),
.Y(n_2229)
);

INVx2_ASAP7_75t_SL g2230 ( 
.A(n_1873),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2026),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_2028),
.Y(n_2232)
);

NOR2x1_ASAP7_75t_L g2233 ( 
.A(n_1920),
.B(n_1863),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2031),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_1787),
.B(n_1515),
.Y(n_2235)
);

NOR2x1_ASAP7_75t_L g2236 ( 
.A(n_1864),
.B(n_1868),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_1796),
.A2(n_1305),
.B1(n_1210),
.B2(n_1292),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2032),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_2036),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2038),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1857),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_1664),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1858),
.Y(n_2243)
);

OA21x2_ASAP7_75t_L g2244 ( 
.A1(n_1860),
.A2(n_1626),
.B(n_1605),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1716),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1903),
.B(n_1393),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1723),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1861),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_1791),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1795),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1798),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1801),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_1870),
.A2(n_1396),
.B1(n_1399),
.B2(n_1393),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1726),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1875),
.B(n_1224),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1728),
.Y(n_2256)
);

INVx6_ASAP7_75t_L g2257 ( 
.A(n_1702),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1802),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1803),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1804),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1808),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1812),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1813),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1870),
.A2(n_1939),
.B1(n_2039),
.B2(n_1805),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1815),
.Y(n_2265)
);

BUFx8_ASAP7_75t_SL g2266 ( 
.A(n_1664),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1816),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1817),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1919),
.B(n_1396),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1822),
.B(n_1525),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1826),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1829),
.Y(n_2272)
);

AND2x6_ASAP7_75t_L g2273 ( 
.A(n_1830),
.B(n_1492),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1957),
.B(n_1399),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1831),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1834),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1835),
.Y(n_2277)
);

NOR2x1_ASAP7_75t_L g2278 ( 
.A(n_1876),
.B(n_1224),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1841),
.Y(n_2279)
);

BUFx8_ASAP7_75t_L g2280 ( 
.A(n_1788),
.Y(n_2280)
);

BUFx12f_ASAP7_75t_L g2281 ( 
.A(n_1671),
.Y(n_2281)
);

INVx4_ASAP7_75t_L g2282 ( 
.A(n_1877),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_1842),
.B(n_1592),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1845),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1849),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1880),
.B(n_1480),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_1939),
.B(n_1406),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_1934),
.B(n_1406),
.Y(n_2288)
);

BUFx8_ASAP7_75t_L g2289 ( 
.A(n_1799),
.Y(n_2289)
);

NOR2x1_ASAP7_75t_L g2290 ( 
.A(n_1881),
.B(n_1594),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1850),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1997),
.B(n_1410),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1852),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1729),
.Y(n_2294)
);

CKINVDCx8_ASAP7_75t_R g2295 ( 
.A(n_1712),
.Y(n_2295)
);

BUFx2_ASAP7_75t_L g2296 ( 
.A(n_1944),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1732),
.Y(n_2297)
);

BUFx8_ASAP7_75t_L g2298 ( 
.A(n_1825),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_1733),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1734),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_1736),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1740),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1745),
.Y(n_2303)
);

OAI21x1_ASAP7_75t_L g2304 ( 
.A1(n_1884),
.A2(n_1634),
.B(n_1626),
.Y(n_2304)
);

OR2x6_ASAP7_75t_L g2305 ( 
.A(n_1844),
.B(n_1091),
.Y(n_2305)
);

AND2x6_ASAP7_75t_L g2306 ( 
.A(n_1886),
.B(n_749),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_1888),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1748),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1753),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1754),
.Y(n_2310)
);

CKINVDCx16_ASAP7_75t_R g2311 ( 
.A(n_1727),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1756),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1890),
.Y(n_2313)
);

INVx5_ASAP7_75t_L g2314 ( 
.A(n_1713),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1757),
.Y(n_2315)
);

OA21x2_ASAP7_75t_L g2316 ( 
.A1(n_2017),
.A2(n_1645),
.B(n_1634),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2029),
.B(n_1410),
.Y(n_2317)
);

AND2x6_ASAP7_75t_L g2318 ( 
.A(n_1892),
.B(n_749),
.Y(n_2318)
);

BUFx12f_ASAP7_75t_L g2319 ( 
.A(n_1671),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1895),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1896),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1898),
.Y(n_2322)
);

HB1xp67_ASAP7_75t_L g2323 ( 
.A(n_1949),
.Y(n_2323)
);

INVx5_ASAP7_75t_L g2324 ( 
.A(n_1724),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1900),
.Y(n_2325)
);

INVx4_ASAP7_75t_L g2326 ( 
.A(n_1904),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_1978),
.B(n_1416),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1907),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_1908),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1912),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1914),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_1797),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_1916),
.B(n_1484),
.Y(n_2333)
);

AND2x6_ASAP7_75t_L g2334 ( 
.A(n_1917),
.B(n_752),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2030),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1987),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_1991),
.B(n_1209),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_1673),
.Y(n_2338)
);

HB1xp67_ASAP7_75t_L g2339 ( 
.A(n_1998),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1764),
.Y(n_2340)
);

INVx6_ASAP7_75t_L g2341 ( 
.A(n_1821),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_SL g2342 ( 
.A1(n_1906),
.A2(n_953),
.B1(n_975),
.B2(n_906),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_1766),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_1913),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_1769),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_1874),
.B(n_1283),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1783),
.B(n_1416),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1790),
.B(n_1417),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_2015),
.Y(n_2349)
);

BUFx8_ASAP7_75t_L g2350 ( 
.A(n_1879),
.Y(n_2350)
);

AND2x6_ASAP7_75t_L g2351 ( 
.A(n_1968),
.B(n_752),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1746),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2023),
.B(n_1417),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1751),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_1959),
.B(n_2037),
.Y(n_2355)
);

AND2x4_ASAP7_75t_L g2356 ( 
.A(n_1953),
.B(n_1323),
.Y(n_2356)
);

OA21x2_ASAP7_75t_L g2357 ( 
.A1(n_1915),
.A2(n_1657),
.B(n_1645),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_1805),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_L g2359 ( 
.A(n_1679),
.B(n_1680),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2027),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_2034),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1823),
.Y(n_2362)
);

INVx4_ASAP7_75t_L g2363 ( 
.A(n_1680),
.Y(n_2363)
);

BUFx2_ASAP7_75t_L g2364 ( 
.A(n_1922),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_1681),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_1681),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1683),
.Y(n_2367)
);

OA21x2_ASAP7_75t_L g2368 ( 
.A1(n_1683),
.A2(n_1657),
.B(n_1489),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1688),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1828),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1688),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_SL g2372 ( 
.A1(n_1910),
.A2(n_975),
.B1(n_1005),
.B2(n_953),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1878),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_1970),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1943),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1979),
.Y(n_2376)
);

OAI21x1_ASAP7_75t_L g2377 ( 
.A1(n_1982),
.A2(n_1491),
.B(n_1486),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1689),
.Y(n_2378)
);

BUFx8_ASAP7_75t_SL g2379 ( 
.A(n_1672),
.Y(n_2379)
);

AOI22x1_ASAP7_75t_SL g2380 ( 
.A1(n_1672),
.A2(n_1008),
.B1(n_1022),
.B2(n_1005),
.Y(n_2380)
);

AOI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_1814),
.A2(n_1429),
.B1(n_1430),
.B2(n_1419),
.Y(n_2381)
);

OA21x2_ASAP7_75t_L g2382 ( 
.A1(n_1689),
.A2(n_1497),
.B(n_1495),
.Y(n_2382)
);

CKINVDCx20_ASAP7_75t_R g2383 ( 
.A(n_1676),
.Y(n_2383)
);

OAI22xp5_ASAP7_75t_SL g2384 ( 
.A1(n_1910),
.A2(n_1022),
.B1(n_1024),
.B2(n_1008),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_1697),
.Y(n_2385)
);

BUFx8_ASAP7_75t_L g2386 ( 
.A(n_2019),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_1697),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_1814),
.B(n_1419),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_1698),
.A2(n_1357),
.B1(n_1378),
.B2(n_1355),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2001),
.B(n_1500),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1698),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1701),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_1701),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_1708),
.B(n_1501),
.Y(n_2394)
);

BUFx6f_ASAP7_75t_L g2395 ( 
.A(n_1708),
.Y(n_2395)
);

OAI22x1_ASAP7_75t_R g2396 ( 
.A1(n_1927),
.A2(n_1075),
.B1(n_1090),
.B2(n_1024),
.Y(n_2396)
);

OA21x2_ASAP7_75t_L g2397 ( 
.A1(n_1709),
.A2(n_1505),
.B(n_1502),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_1709),
.B(n_1506),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1711),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_1711),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_1818),
.B(n_1429),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1717),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_1717),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_1818),
.A2(n_1435),
.B1(n_1441),
.B2(n_1430),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_1720),
.B(n_1507),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_1720),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_1725),
.B(n_1435),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_1725),
.B(n_1509),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_1827),
.Y(n_2409)
);

OAI21x1_ASAP7_75t_L g2410 ( 
.A1(n_1827),
.A2(n_1511),
.B(n_1510),
.Y(n_2410)
);

AND2x6_ASAP7_75t_L g2411 ( 
.A(n_1832),
.B(n_755),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1832),
.Y(n_2412)
);

BUFx12f_ASAP7_75t_L g2413 ( 
.A(n_1838),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_1838),
.B(n_1520),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_1853),
.A2(n_1527),
.B(n_1522),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_1853),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_1854),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1854),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_1855),
.B(n_1532),
.Y(n_2419)
);

CKINVDCx11_ASAP7_75t_R g2420 ( 
.A(n_1927),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_1855),
.Y(n_2421)
);

OAI21x1_ASAP7_75t_L g2422 ( 
.A1(n_1871),
.A2(n_1538),
.B(n_1535),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_1871),
.B(n_1539),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1883),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1883),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1887),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_1887),
.B(n_1547),
.Y(n_2427)
);

AND2x2_ASAP7_75t_SL g2428 ( 
.A(n_1889),
.B(n_819),
.Y(n_2428)
);

BUFx12f_ASAP7_75t_L g2429 ( 
.A(n_1889),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_1894),
.B(n_1441),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_1894),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_1897),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_L g2433 ( 
.A(n_1930),
.B(n_1549),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_1897),
.Y(n_2434)
);

INVx3_ASAP7_75t_L g2435 ( 
.A(n_1901),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_1901),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1902),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1902),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_1909),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_1909),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1921),
.Y(n_2441)
);

CKINVDCx8_ASAP7_75t_R g2442 ( 
.A(n_1921),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1925),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1925),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_1928),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1928),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1933),
.B(n_1444),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1933),
.B(n_1444),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_1942),
.B(n_1551),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_1942),
.B(n_1554),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_1947),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1947),
.B(n_1445),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_1952),
.B(n_1445),
.Y(n_2453)
);

INVx5_ASAP7_75t_L g2454 ( 
.A(n_1952),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_1965),
.Y(n_2455)
);

INVx6_ASAP7_75t_L g2456 ( 
.A(n_2039),
.Y(n_2456)
);

OA21x2_ASAP7_75t_L g2457 ( 
.A1(n_1965),
.A2(n_1556),
.B(n_1555),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_1969),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_SL g2459 ( 
.A1(n_1676),
.A2(n_1149),
.B1(n_1075),
.B2(n_1104),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1969),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1972),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1972),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_1976),
.B(n_1450),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_1976),
.A2(n_2013),
.B1(n_1981),
.B2(n_1984),
.Y(n_2464)
);

INVx2_ASAP7_75t_SL g2465 ( 
.A(n_1980),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_1980),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_1981),
.A2(n_833),
.B1(n_863),
.B2(n_842),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1984),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1999),
.B(n_1450),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1999),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2218),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2084),
.B(n_2013),
.Y(n_2472)
);

BUFx6f_ASAP7_75t_L g2473 ( 
.A(n_2050),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2042),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2042),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2046),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2046),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2107),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2060),
.Y(n_2479)
);

NAND2x1p5_ASAP7_75t_L g2480 ( 
.A(n_2212),
.B(n_1557),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2107),
.B(n_1460),
.Y(n_2481)
);

NAND2xp33_ASAP7_75t_L g2482 ( 
.A(n_2412),
.B(n_1454),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_2218),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2048),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2218),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2050),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2060),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_2220),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2052),
.B(n_1948),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_2220),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2086),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2086),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2048),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2127),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2053),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2050),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2050),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2127),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2053),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2136),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2136),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2054),
.Y(n_2502)
);

AND2x4_ASAP7_75t_L g2503 ( 
.A(n_2052),
.B(n_1948),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2220),
.Y(n_2504)
);

OR2x6_ASAP7_75t_L g2505 ( 
.A(n_2230),
.B(n_1558),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2355),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2390),
.B(n_1460),
.Y(n_2507)
);

CKINVDCx20_ASAP7_75t_R g2508 ( 
.A(n_2386),
.Y(n_2508)
);

OA21x2_ASAP7_75t_L g2509 ( 
.A1(n_2304),
.A2(n_1561),
.B(n_1560),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2140),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2140),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2390),
.B(n_1461),
.Y(n_2512)
);

AND2x4_ASAP7_75t_L g2513 ( 
.A(n_2052),
.B(n_1971),
.Y(n_2513)
);

AND2x6_ASAP7_75t_L g2514 ( 
.A(n_2040),
.B(n_755),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2150),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2150),
.Y(n_2516)
);

HB1xp67_ASAP7_75t_L g2517 ( 
.A(n_2355),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2054),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2055),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2055),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2059),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2050),
.Y(n_2522)
);

INVxp67_ASAP7_75t_L g2523 ( 
.A(n_2199),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2059),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2065),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2065),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2066),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2066),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2072),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2072),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2080),
.Y(n_2531)
);

AND2x4_ASAP7_75t_L g2532 ( 
.A(n_2040),
.B(n_2044),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2454),
.B(n_1462),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2454),
.B(n_1462),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2080),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2344),
.B(n_1496),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2081),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2187),
.Y(n_2538)
);

BUFx3_ASAP7_75t_L g2539 ( 
.A(n_2341),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2187),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2068),
.B(n_2330),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2081),
.Y(n_2542)
);

BUFx6f_ASAP7_75t_L g2543 ( 
.A(n_2061),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2094),
.Y(n_2544)
);

INVxp67_ASAP7_75t_L g2545 ( 
.A(n_2077),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2094),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2095),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2095),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2098),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2098),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2099),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2040),
.B(n_2006),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2099),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2330),
.B(n_1454),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2103),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_L g2556 ( 
.A(n_2374),
.B(n_1954),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2044),
.B(n_2435),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2183),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2103),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2112),
.Y(n_2560)
);

AND2x4_ASAP7_75t_L g2561 ( 
.A(n_2044),
.B(n_2018),
.Y(n_2561)
);

INVxp67_ASAP7_75t_L g2562 ( 
.A(n_2043),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2112),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2183),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2092),
.Y(n_2565)
);

OA21x2_ASAP7_75t_L g2566 ( 
.A1(n_2304),
.A2(n_1566),
.B(n_1564),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2116),
.Y(n_2567)
);

BUFx8_ASAP7_75t_L g2568 ( 
.A(n_2192),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2187),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2330),
.B(n_1457),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2116),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2119),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2119),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2123),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2196),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2123),
.Y(n_2576)
);

AND2x2_ASAP7_75t_SL g2577 ( 
.A(n_2428),
.B(n_819),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2344),
.B(n_2083),
.Y(n_2578)
);

OA21x2_ASAP7_75t_L g2579 ( 
.A1(n_2225),
.A2(n_1570),
.B(n_1569),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2124),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2124),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2131),
.Y(n_2582)
);

NAND2xp33_ASAP7_75t_L g2583 ( 
.A(n_2412),
.B(n_1457),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2131),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2435),
.B(n_1954),
.Y(n_2585)
);

OA21x2_ASAP7_75t_L g2586 ( 
.A1(n_2225),
.A2(n_1575),
.B(n_1573),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2335),
.B(n_1458),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2132),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2196),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2132),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2141),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2141),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2143),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2143),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2196),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2149),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2149),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2160),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2244),
.Y(n_2599)
);

AOI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2428),
.A2(n_1104),
.B1(n_1106),
.B2(n_1090),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2117),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2244),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2192),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2244),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2194),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2160),
.Y(n_2606)
);

BUFx3_ASAP7_75t_L g2607 ( 
.A(n_2341),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2454),
.B(n_2412),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2162),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2117),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2435),
.B(n_1955),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2194),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2117),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2057),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2162),
.Y(n_2615)
);

OAI22xp5_ASAP7_75t_SL g2616 ( 
.A1(n_2158),
.A2(n_1112),
.B1(n_1149),
.B2(n_1106),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2335),
.B(n_1458),
.Y(n_2617)
);

OAI21x1_ASAP7_75t_L g2618 ( 
.A1(n_2069),
.A2(n_1579),
.B(n_1577),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2186),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2299),
.B(n_1461),
.Y(n_2620)
);

AND2x4_ASAP7_75t_L g2621 ( 
.A(n_2439),
.B(n_2018),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2151),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2151),
.Y(n_2623)
);

INVx1_ASAP7_75t_SL g2624 ( 
.A(n_2057),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2186),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2151),
.Y(n_2626)
);

OAI21x1_ASAP7_75t_L g2627 ( 
.A1(n_2069),
.A2(n_1580),
.B(n_764),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2188),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2296),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2176),
.Y(n_2630)
);

BUFx6f_ASAP7_75t_L g2631 ( 
.A(n_2176),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2296),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2454),
.B(n_1496),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2341),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2454),
.B(n_1498),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2188),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2161),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2191),
.Y(n_2638)
);

INVx3_ASAP7_75t_L g2639 ( 
.A(n_2161),
.Y(n_2639)
);

OA21x2_ASAP7_75t_L g2640 ( 
.A1(n_2102),
.A2(n_764),
.B(n_758),
.Y(n_2640)
);

NAND2xp33_ASAP7_75t_SL g2641 ( 
.A(n_2412),
.B(n_1961),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2191),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2161),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2211),
.Y(n_2644)
);

BUFx2_ASAP7_75t_L g2645 ( 
.A(n_2346),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2341),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2211),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2102),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2083),
.B(n_1471),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2299),
.B(n_2301),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2412),
.B(n_1471),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2138),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2439),
.B(n_1955),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2211),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2216),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2092),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2346),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2216),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2138),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2316),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2316),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2216),
.Y(n_2662)
);

INVx3_ASAP7_75t_L g2663 ( 
.A(n_2157),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2316),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2238),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2083),
.B(n_1472),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2238),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2238),
.Y(n_2668)
);

NAND2x1_ASAP7_75t_L g2669 ( 
.A(n_2174),
.B(n_1229),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2299),
.B(n_2301),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2301),
.B(n_1472),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2226),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_L g2673 ( 
.A1(n_2377),
.A2(n_769),
.B(n_758),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2240),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2411),
.B(n_1477),
.Y(n_2675)
);

OAI21x1_ASAP7_75t_L g2676 ( 
.A1(n_2377),
.A2(n_773),
.B(n_769),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2226),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2226),
.Y(n_2678)
);

BUFx6f_ASAP7_75t_L g2679 ( 
.A(n_2176),
.Y(n_2679)
);

INVx3_ASAP7_75t_L g2680 ( 
.A(n_2157),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2240),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2157),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2240),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2228),
.Y(n_2684)
);

XNOR2xp5_ASAP7_75t_L g2685 ( 
.A(n_2459),
.B(n_1629),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2228),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2228),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2155),
.Y(n_2688)
);

OR2x2_ASAP7_75t_L g2689 ( 
.A(n_2346),
.B(n_1477),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2155),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2411),
.B(n_1481),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2157),
.Y(n_2692)
);

INVx1_ASAP7_75t_SL g2693 ( 
.A(n_2148),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2159),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2159),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2416),
.B(n_1493),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2168),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2168),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2146),
.Y(n_2699)
);

OA21x2_ASAP7_75t_L g2700 ( 
.A1(n_2106),
.A2(n_774),
.B(n_773),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2177),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2146),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2411),
.B(n_1481),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_2257),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2089),
.B(n_1498),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2356),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2146),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2146),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2146),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2177),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2056),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2179),
.Y(n_2712)
);

BUFx2_ASAP7_75t_L g2713 ( 
.A(n_2356),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2439),
.B(n_1971),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2179),
.Y(n_2715)
);

CKINVDCx16_ASAP7_75t_R g2716 ( 
.A(n_2311),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2197),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2176),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2197),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2411),
.B(n_1483),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2056),
.Y(n_2721)
);

INVx3_ASAP7_75t_L g2722 ( 
.A(n_2157),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2056),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2210),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2210),
.Y(n_2725)
);

BUFx8_ASAP7_75t_L g2726 ( 
.A(n_2126),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2163),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2176),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2145),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2163),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2062),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2356),
.Y(n_2732)
);

INVx3_ASAP7_75t_L g2733 ( 
.A(n_2163),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2089),
.B(n_1504),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2221),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2411),
.B(n_1483),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2190),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2062),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2190),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2062),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2190),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2357),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2357),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2221),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2231),
.Y(n_2745)
);

BUFx6f_ASAP7_75t_L g2746 ( 
.A(n_2190),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2231),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2357),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2190),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_2305),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2234),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2193),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2411),
.B(n_2248),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2193),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2234),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2248),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2248),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2265),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2265),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2265),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2163),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2260),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2089),
.B(n_1508),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2147),
.Y(n_2764)
);

INVx1_ASAP7_75t_SL g2765 ( 
.A(n_2148),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2451),
.B(n_2006),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2163),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2203),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2164),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2093),
.B(n_1508),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_L g2771 ( 
.A1(n_2071),
.A2(n_777),
.B(n_774),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2260),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2193),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2261),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2282),
.B(n_1493),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2203),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2203),
.Y(n_2777)
);

CKINVDCx20_ASAP7_75t_R g2778 ( 
.A(n_2386),
.Y(n_2778)
);

NAND2xp33_ASAP7_75t_SL g2779 ( 
.A(n_2416),
.B(n_1961),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2261),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2203),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2268),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2203),
.Y(n_2783)
);

BUFx2_ASAP7_75t_L g2784 ( 
.A(n_2305),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2416),
.B(n_1517),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2207),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2268),
.Y(n_2787)
);

HB1xp67_ASAP7_75t_L g2788 ( 
.A(n_2323),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2271),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2271),
.Y(n_2790)
);

OA21x2_ASAP7_75t_L g2791 ( 
.A1(n_2153),
.A2(n_783),
.B(n_777),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2279),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2279),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2284),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2164),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2284),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2207),
.Y(n_2797)
);

NAND2xp33_ASAP7_75t_L g2798 ( 
.A(n_2416),
.B(n_1494),
.Y(n_2798)
);

HB1xp67_ASAP7_75t_L g2799 ( 
.A(n_2339),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2321),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2193),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2321),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2207),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2207),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2242),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2193),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2207),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2282),
.B(n_1494),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2282),
.B(n_1504),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2325),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2208),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2208),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2325),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2241),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2164),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2241),
.Y(n_2816)
);

BUFx6f_ASAP7_75t_L g2817 ( 
.A(n_2164),
.Y(n_2817)
);

OAI21x1_ASAP7_75t_L g2818 ( 
.A1(n_2170),
.A2(n_784),
.B(n_783),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2164),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2250),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2250),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2251),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2093),
.B(n_2108),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2251),
.Y(n_2824)
);

HB1xp67_ASAP7_75t_L g2825 ( 
.A(n_2242),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2252),
.Y(n_2826)
);

NAND2x1p5_ASAP7_75t_L g2827 ( 
.A(n_2212),
.B(n_784),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2257),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2208),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2208),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2252),
.Y(n_2831)
);

INVx1_ASAP7_75t_SL g2832 ( 
.A(n_2383),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2208),
.Y(n_2833)
);

AOI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2306),
.A2(n_1153),
.B1(n_1177),
.B2(n_1112),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2223),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2223),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2051),
.Y(n_2837)
);

AND2x4_ASAP7_75t_L g2838 ( 
.A(n_2451),
.B(n_2466),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2383),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2267),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2267),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2326),
.B(n_1514),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2223),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2051),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2223),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2093),
.B(n_2108),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2326),
.B(n_1514),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2275),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2275),
.Y(n_2849)
);

OAI21x1_ASAP7_75t_L g2850 ( 
.A1(n_2182),
.A2(n_2415),
.B(n_2410),
.Y(n_2850)
);

HB1xp67_ASAP7_75t_L g2851 ( 
.A(n_2214),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2276),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2410),
.A2(n_799),
.B(n_790),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2223),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2276),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2277),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2224),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2277),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2285),
.Y(n_2859)
);

BUFx2_ASAP7_75t_L g2860 ( 
.A(n_2305),
.Y(n_2860)
);

HB1xp67_ASAP7_75t_L g2861 ( 
.A(n_2214),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2285),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2224),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2291),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2224),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2291),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2451),
.B(n_1974),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2224),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2224),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2466),
.B(n_1974),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2320),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2320),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2322),
.Y(n_2873)
);

OA21x2_ASAP7_75t_L g2874 ( 
.A1(n_2415),
.A2(n_799),
.B(n_790),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2322),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2227),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2305),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2331),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2331),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_2115),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2227),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2051),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2108),
.B(n_1546),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2297),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2297),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2300),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2300),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2115),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2303),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2303),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2309),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2189),
.B(n_1516),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2309),
.Y(n_2893)
);

AND2x6_ASAP7_75t_L g2894 ( 
.A(n_2414),
.B(n_2427),
.Y(n_2894)
);

BUFx3_ASAP7_75t_L g2895 ( 
.A(n_2257),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2287),
.B(n_1516),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2310),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2310),
.Y(n_2898)
);

INVxp67_ASAP7_75t_L g2899 ( 
.A(n_2266),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_2416),
.B(n_2421),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2227),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2227),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2326),
.B(n_1517),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2041),
.Y(n_2904)
);

INVxp67_ASAP7_75t_L g2905 ( 
.A(n_2266),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2227),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2229),
.Y(n_2907)
);

OAI22xp33_ASAP7_75t_R g2908 ( 
.A1(n_2430),
.A2(n_673),
.B1(n_685),
.B2(n_678),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2154),
.B(n_1524),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2229),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2421),
.B(n_1524),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2045),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2154),
.B(n_1528),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2294),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2229),
.Y(n_2915)
);

HB1xp67_ASAP7_75t_L g2916 ( 
.A(n_2379),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2229),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2474),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2892),
.B(n_2466),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2630),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2630),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2484),
.Y(n_2922)
);

OR2x6_ASAP7_75t_L g2923 ( 
.A(n_2532),
.B(n_2230),
.Y(n_2923)
);

INVx3_ASAP7_75t_L g2924 ( 
.A(n_2630),
.Y(n_2924)
);

NAND2xp33_ASAP7_75t_L g2925 ( 
.A(n_2894),
.B(n_2421),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2896),
.B(n_2463),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2645),
.Y(n_2927)
);

AO22x2_ASAP7_75t_L g2928 ( 
.A1(n_2600),
.A2(n_2380),
.B1(n_2396),
.B2(n_2414),
.Y(n_2928)
);

NAND2xp33_ASAP7_75t_L g2929 ( 
.A(n_2894),
.B(n_2421),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2474),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_L g2931 ( 
.A1(n_2600),
.A2(n_2351),
.B1(n_2457),
.B2(n_2397),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2484),
.Y(n_2932)
);

INVx2_ASAP7_75t_SL g2933 ( 
.A(n_2532),
.Y(n_2933)
);

INVx3_ASAP7_75t_L g2934 ( 
.A(n_2630),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2493),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2475),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2493),
.Y(n_2937)
);

INVx4_ASAP7_75t_L g2938 ( 
.A(n_2630),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2729),
.B(n_2419),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2475),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2495),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2495),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2476),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2499),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2499),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2532),
.B(n_2421),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2577),
.A2(n_2306),
.B1(n_2334),
.B2(n_2318),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2502),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2502),
.Y(n_2949)
);

INVx3_ASAP7_75t_L g2950 ( 
.A(n_2630),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2838),
.B(n_2419),
.Y(n_2951)
);

OR2x2_ASAP7_75t_L g2952 ( 
.A(n_2693),
.B(n_2364),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2472),
.B(n_2104),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2476),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2477),
.Y(n_2955)
);

BUFx8_ASAP7_75t_SL g2956 ( 
.A(n_2508),
.Y(n_2956)
);

AND2x6_ASAP7_75t_L g2957 ( 
.A(n_2532),
.B(n_2440),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2477),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2520),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2520),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2521),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2624),
.B(n_2104),
.Y(n_2962)
);

OR2x2_ASAP7_75t_L g2963 ( 
.A(n_2765),
.B(n_2364),
.Y(n_2963)
);

INVx3_ASAP7_75t_L g2964 ( 
.A(n_2631),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2521),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2631),
.Y(n_2966)
);

INVx2_ASAP7_75t_SL g2967 ( 
.A(n_2704),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2479),
.Y(n_2968)
);

INVxp67_ASAP7_75t_SL g2969 ( 
.A(n_2631),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2631),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2631),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2524),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2556),
.B(n_2156),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2524),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2631),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2479),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2557),
.B(n_2440),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2523),
.B(n_2181),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2487),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2487),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2689),
.B(n_2195),
.Y(n_2981)
);

INVx5_ASAP7_75t_L g2982 ( 
.A(n_2679),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2525),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2689),
.B(n_2195),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2491),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2491),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2557),
.B(n_2440),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2492),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2525),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2565),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_2557),
.B(n_2440),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2679),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2531),
.Y(n_2993)
);

INVx3_ASAP7_75t_L g2994 ( 
.A(n_2679),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2531),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2679),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2838),
.B(n_2423),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2577),
.A2(n_2351),
.B1(n_2457),
.B2(n_2397),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2492),
.Y(n_2999)
);

INVx2_ASAP7_75t_SL g3000 ( 
.A(n_2704),
.Y(n_3000)
);

BUFx2_ASAP7_75t_L g3001 ( 
.A(n_2564),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2535),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2535),
.Y(n_3003)
);

OR2x6_ASAP7_75t_L g3004 ( 
.A(n_2505),
.B(n_2257),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2838),
.B(n_2423),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2494),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2494),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2498),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2498),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2577),
.A2(n_2351),
.B1(n_2457),
.B2(n_2397),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2500),
.Y(n_3011)
);

CKINVDCx6p67_ASAP7_75t_R g3012 ( 
.A(n_2716),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2542),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2542),
.Y(n_3014)
);

CKINVDCx20_ASAP7_75t_R g3015 ( 
.A(n_2716),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2500),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2823),
.B(n_2449),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2544),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2562),
.B(n_2202),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_SL g3020 ( 
.A(n_2557),
.B(n_2440),
.Y(n_3020)
);

INVx3_ASAP7_75t_L g3021 ( 
.A(n_2679),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2544),
.Y(n_3022)
);

NOR3xp33_ASAP7_75t_L g3023 ( 
.A(n_2536),
.B(n_2359),
.C(n_2205),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2549),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2501),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2838),
.B(n_2449),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2549),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2679),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2501),
.Y(n_3029)
);

INVx5_ASAP7_75t_L g3030 ( 
.A(n_2718),
.Y(n_3030)
);

INVx3_ASAP7_75t_L g3031 ( 
.A(n_2718),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2507),
.B(n_2455),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2550),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_SL g3034 ( 
.A(n_2507),
.B(n_2455),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2550),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2571),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2510),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2510),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2511),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2571),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2511),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2574),
.Y(n_3042)
);

BUFx2_ASAP7_75t_L g3043 ( 
.A(n_2564),
.Y(n_3043)
);

INVx4_ASAP7_75t_L g3044 ( 
.A(n_2718),
.Y(n_3044)
);

HB1xp67_ASAP7_75t_L g3045 ( 
.A(n_2713),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2908),
.A2(n_2894),
.B1(n_2616),
.B2(n_2834),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2515),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2574),
.Y(n_3048)
);

INVx8_ASAP7_75t_L g3049 ( 
.A(n_2894),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2908),
.A2(n_2351),
.B1(n_2382),
.B2(n_2318),
.Y(n_3050)
);

INVxp67_ASAP7_75t_L g3051 ( 
.A(n_2764),
.Y(n_3051)
);

AO22x2_ASAP7_75t_L g3052 ( 
.A1(n_2834),
.A2(n_2380),
.B1(n_2427),
.B2(n_2414),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2512),
.B(n_2445),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2580),
.Y(n_3054)
);

XNOR2xp5_ASAP7_75t_L g3055 ( 
.A(n_2685),
.B(n_2088),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2823),
.B(n_2450),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2515),
.Y(n_3057)
);

NAND2xp33_ASAP7_75t_L g3058 ( 
.A(n_2894),
.B(n_2445),
.Y(n_3058)
);

BUFx3_ASAP7_75t_L g3059 ( 
.A(n_2828),
.Y(n_3059)
);

BUFx10_ASAP7_75t_L g3060 ( 
.A(n_2585),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2656),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2894),
.B(n_2512),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2894),
.B(n_2450),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2516),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2516),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2718),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2598),
.Y(n_3067)
);

INVx2_ASAP7_75t_SL g3068 ( 
.A(n_2828),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2688),
.B(n_2338),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2775),
.B(n_2445),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2580),
.Y(n_3071)
);

OR2x6_ASAP7_75t_L g3072 ( 
.A(n_2505),
.B(n_2445),
.Y(n_3072)
);

CKINVDCx6p67_ASAP7_75t_R g3073 ( 
.A(n_2778),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2581),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2581),
.Y(n_3075)
);

CKINVDCx20_ASAP7_75t_R g3076 ( 
.A(n_2726),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_SL g3077 ( 
.A(n_2552),
.Y(n_3077)
);

OAI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2657),
.A2(n_2205),
.B1(n_2215),
.B2(n_2202),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2593),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_SL g3080 ( 
.A1(n_2616),
.A2(n_2342),
.B1(n_2384),
.B2(n_2372),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_SL g3081 ( 
.A(n_2808),
.B(n_2445),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2598),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2593),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_SL g3084 ( 
.A1(n_2585),
.A2(n_2142),
.B1(n_2351),
.B2(n_2455),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2688),
.B(n_2338),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2718),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2594),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2594),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2518),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2690),
.B(n_2338),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2518),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2606),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2519),
.Y(n_3093)
);

AND2x2_ASAP7_75t_SL g3094 ( 
.A(n_2753),
.B(n_2382),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2606),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2690),
.B(n_2366),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2519),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2609),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2694),
.B(n_2366),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2609),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2694),
.B(n_2366),
.Y(n_3101)
);

INVx1_ASAP7_75t_SL g3102 ( 
.A(n_2558),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2615),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2526),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2695),
.B(n_2400),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_2809),
.B(n_2455),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2615),
.Y(n_3107)
);

NAND2xp33_ASAP7_75t_R g3108 ( 
.A(n_2585),
.B(n_2215),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_2726),
.Y(n_3109)
);

INVx3_ASAP7_75t_L g3110 ( 
.A(n_2718),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2846),
.B(n_2578),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_2726),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2526),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2603),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2895),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2619),
.Y(n_3116)
);

OAI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2706),
.A2(n_2358),
.B1(n_2434),
.B2(n_2332),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2619),
.Y(n_3118)
);

INVx6_ASAP7_75t_L g3119 ( 
.A(n_2728),
.Y(n_3119)
);

HB1xp67_ASAP7_75t_L g3120 ( 
.A(n_2732),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2527),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2514),
.A2(n_2306),
.B1(n_2334),
.B2(n_2318),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2842),
.B(n_2455),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_2847),
.B(n_2365),
.Y(n_3124)
);

OA22x2_ASAP7_75t_L g3125 ( 
.A1(n_2846),
.A2(n_2685),
.B1(n_2088),
.B2(n_2750),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2545),
.B(n_2332),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2527),
.Y(n_3127)
);

INVx2_ASAP7_75t_SL g3128 ( 
.A(n_2895),
.Y(n_3128)
);

NAND3xp33_ASAP7_75t_L g3129 ( 
.A(n_2482),
.B(n_2407),
.C(n_2460),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2528),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_SL g3131 ( 
.A(n_2552),
.Y(n_3131)
);

NAND3xp33_ASAP7_75t_L g3132 ( 
.A(n_2583),
.B(n_2461),
.C(n_2460),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2728),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_SL g3134 ( 
.A(n_2552),
.Y(n_3134)
);

AOI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_2514),
.A2(n_2306),
.B1(n_2334),
.B2(n_2318),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2903),
.B(n_2365),
.Y(n_3136)
);

INVx3_ASAP7_75t_L g3137 ( 
.A(n_2728),
.Y(n_3137)
);

BUFx10_ASAP7_75t_L g3138 ( 
.A(n_2585),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2528),
.Y(n_3139)
);

BUFx6f_ASAP7_75t_L g3140 ( 
.A(n_2728),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2529),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2695),
.B(n_2400),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2625),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2529),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2530),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2530),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2537),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2537),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2539),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2578),
.B(n_2365),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2625),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2546),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2536),
.B(n_2358),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_2728),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2697),
.B(n_2400),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2546),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2547),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2628),
.Y(n_3158)
);

INVx5_ASAP7_75t_L g3159 ( 
.A(n_2728),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2547),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2628),
.Y(n_3161)
);

OR2x2_ASAP7_75t_L g3162 ( 
.A(n_2832),
.B(n_2434),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2636),
.Y(n_3163)
);

CKINVDCx5p33_ASAP7_75t_R g3164 ( 
.A(n_2726),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2636),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2697),
.B(n_2408),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2638),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2638),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2698),
.B(n_2701),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2909),
.B(n_2070),
.Y(n_3170)
);

OR2x6_ASAP7_75t_L g3171 ( 
.A(n_2505),
.B(n_2365),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2548),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2642),
.Y(n_3173)
);

HB1xp67_ASAP7_75t_L g3174 ( 
.A(n_2629),
.Y(n_3174)
);

NAND2xp33_ASAP7_75t_L g3175 ( 
.A(n_2737),
.B(n_2340),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2642),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_2909),
.B(n_2070),
.Y(n_3177)
);

NOR3xp33_ASAP7_75t_L g3178 ( 
.A(n_2614),
.B(n_2359),
.C(n_2465),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2548),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2551),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_2913),
.A2(n_2351),
.B1(n_2382),
.B2(n_2318),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2551),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2553),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2553),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2555),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_2913),
.A2(n_2318),
.B1(n_2334),
.B2(n_2306),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2555),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2559),
.Y(n_3188)
);

BUFx10_ASAP7_75t_L g3189 ( 
.A(n_2611),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2559),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2632),
.B(n_2465),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2560),
.Y(n_3192)
);

NAND2xp33_ASAP7_75t_L g3193 ( 
.A(n_2737),
.B(n_2340),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2560),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2563),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2563),
.Y(n_3196)
);

INVxp33_ASAP7_75t_L g3197 ( 
.A(n_2805),
.Y(n_3197)
);

BUFx6f_ASAP7_75t_L g3198 ( 
.A(n_2737),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_2737),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2567),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_2554),
.B(n_2365),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2567),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_SL g3203 ( 
.A(n_2827),
.B(n_2413),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2737),
.Y(n_3204)
);

INVx1_ASAP7_75t_SL g3205 ( 
.A(n_2788),
.Y(n_3205)
);

INVx3_ASAP7_75t_L g3206 ( 
.A(n_2737),
.Y(n_3206)
);

BUFx2_ASAP7_75t_L g3207 ( 
.A(n_2568),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2570),
.B(n_2385),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2572),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2572),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2698),
.B(n_2408),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2573),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2573),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2576),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2576),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2582),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2582),
.Y(n_3217)
);

NAND2xp33_ASAP7_75t_L g3218 ( 
.A(n_2739),
.B(n_2340),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_2701),
.B(n_2070),
.Y(n_3219)
);

BUFx3_ASAP7_75t_L g3220 ( 
.A(n_2539),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2584),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2588),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2588),
.Y(n_3223)
);

INVx4_ASAP7_75t_L g3224 ( 
.A(n_2739),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2590),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2590),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2591),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2591),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2592),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2478),
.B(n_2456),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2620),
.B(n_2385),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_2671),
.B(n_2385),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2592),
.Y(n_3233)
);

BUFx6f_ASAP7_75t_L g3234 ( 
.A(n_2739),
.Y(n_3234)
);

INVx5_ASAP7_75t_L g3235 ( 
.A(n_2739),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2596),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_2481),
.B(n_2456),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2596),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2597),
.Y(n_3239)
);

INVx3_ASAP7_75t_L g3240 ( 
.A(n_2739),
.Y(n_3240)
);

BUFx2_ASAP7_75t_L g3241 ( 
.A(n_2568),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2597),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_2618),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2710),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2710),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2712),
.B(n_2409),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2481),
.B(n_2456),
.Y(n_3247)
);

INVx5_ASAP7_75t_L g3248 ( 
.A(n_2739),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_2741),
.Y(n_3249)
);

BUFx10_ASAP7_75t_L g3250 ( 
.A(n_2611),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_2741),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_2799),
.B(n_2456),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2607),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2618),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2712),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2715),
.Y(n_3256)
);

BUFx6f_ASAP7_75t_L g3257 ( 
.A(n_2741),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2715),
.B(n_2409),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2579),
.Y(n_3259)
);

INVx5_ASAP7_75t_L g3260 ( 
.A(n_2741),
.Y(n_3260)
);

NOR2xp33_ASAP7_75t_L g3261 ( 
.A(n_2506),
.B(n_2464),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_2579),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_2514),
.A2(n_2306),
.B1(n_2334),
.B2(n_2273),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2579),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2517),
.B(n_2264),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2579),
.Y(n_3266)
);

INVx4_ASAP7_75t_L g3267 ( 
.A(n_2741),
.Y(n_3267)
);

INVx5_ASAP7_75t_L g3268 ( 
.A(n_2741),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_2607),
.B(n_2212),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2762),
.Y(n_3270)
);

BUFx6f_ASAP7_75t_L g3271 ( 
.A(n_2746),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2586),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2586),
.Y(n_3273)
);

INVx1_ASAP7_75t_SL g3274 ( 
.A(n_2825),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2762),
.B(n_2772),
.Y(n_3275)
);

BUFx6f_ASAP7_75t_L g3276 ( 
.A(n_2746),
.Y(n_3276)
);

BUFx3_ASAP7_75t_L g3277 ( 
.A(n_2634),
.Y(n_3277)
);

AOI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_2514),
.A2(n_2334),
.B1(n_2273),
.B2(n_2076),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_2586),
.Y(n_3279)
);

CKINVDCx5p33_ASAP7_75t_R g3280 ( 
.A(n_2568),
.Y(n_3280)
);

INVx3_ASAP7_75t_L g3281 ( 
.A(n_2746),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2772),
.Y(n_3282)
);

HB1xp67_ASAP7_75t_L g3283 ( 
.A(n_2839),
.Y(n_3283)
);

NAND2xp33_ASAP7_75t_SL g3284 ( 
.A(n_2587),
.B(n_2340),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2774),
.B(n_2431),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_2634),
.B(n_2385),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_2646),
.B(n_2212),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2774),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2586),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2613),
.Y(n_3290)
);

OAI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_2617),
.A2(n_2442),
.B1(n_2385),
.B2(n_2402),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2613),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2780),
.B(n_2431),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2780),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2782),
.Y(n_3295)
);

BUFx6f_ASAP7_75t_L g3296 ( 
.A(n_2746),
.Y(n_3296)
);

BUFx6f_ASAP7_75t_L g3297 ( 
.A(n_2746),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2782),
.Y(n_3298)
);

INVx2_ASAP7_75t_SL g3299 ( 
.A(n_2646),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2787),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2787),
.B(n_2432),
.Y(n_3301)
);

INVx4_ASAP7_75t_SL g3302 ( 
.A(n_2514),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_2649),
.B(n_2442),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_2746),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_2789),
.B(n_2255),
.Y(n_3305)
);

INVx3_ASAP7_75t_L g3306 ( 
.A(n_2749),
.Y(n_3306)
);

BUFx6f_ASAP7_75t_L g3307 ( 
.A(n_2749),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2622),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2789),
.B(n_2255),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2649),
.B(n_2461),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_2552),
.B(n_2395),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_2561),
.B(n_2395),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_2622),
.Y(n_3313)
);

BUFx6f_ASAP7_75t_L g3314 ( 
.A(n_2749),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2790),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2623),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2790),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2792),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_2792),
.B(n_2427),
.Y(n_3319)
);

BUFx6f_ASAP7_75t_L g3320 ( 
.A(n_2749),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2793),
.Y(n_3321)
);

INVxp33_ASAP7_75t_L g3322 ( 
.A(n_2666),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_2623),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_2626),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2794),
.Y(n_3325)
);

OR2x6_ASAP7_75t_L g3326 ( 
.A(n_2505),
.B(n_2395),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_2794),
.B(n_2432),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2796),
.B(n_2436),
.Y(n_3328)
);

INVx2_ASAP7_75t_SL g3329 ( 
.A(n_2505),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2561),
.B(n_2395),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2626),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_2637),
.Y(n_3332)
);

NAND2xp33_ASAP7_75t_L g3333 ( 
.A(n_2749),
.B(n_2340),
.Y(n_3333)
);

INVx5_ASAP7_75t_L g3334 ( 
.A(n_2749),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_2637),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_2643),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_2643),
.Y(n_3337)
);

XOR2xp5_ASAP7_75t_L g3338 ( 
.A(n_2561),
.B(n_1677),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_2752),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2796),
.Y(n_3340)
);

AND2x6_ASAP7_75t_L g3341 ( 
.A(n_2752),
.B(n_2395),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2871),
.Y(n_3342)
);

INVx5_ASAP7_75t_L g3343 ( 
.A(n_2752),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_2827),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2871),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_2752),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_2509),
.Y(n_3347)
);

BUFx6f_ASAP7_75t_L g3348 ( 
.A(n_2752),
.Y(n_3348)
);

CKINVDCx5p33_ASAP7_75t_R g3349 ( 
.A(n_2568),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2509),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2509),
.Y(n_3351)
);

BUFx6f_ASAP7_75t_L g3352 ( 
.A(n_2754),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_2509),
.Y(n_3353)
);

BUFx2_ASAP7_75t_L g3354 ( 
.A(n_2489),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_2666),
.B(n_2462),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2872),
.B(n_2873),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_2566),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_2872),
.B(n_2144),
.Y(n_3358)
);

CKINVDCx5p33_ASAP7_75t_R g3359 ( 
.A(n_2851),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_2754),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2873),
.B(n_2436),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_2561),
.B(n_2402),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2566),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2875),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_2566),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_2875),
.Y(n_3366)
);

OAI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_2750),
.A2(n_2402),
.B1(n_2363),
.B2(n_2343),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_2754),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_2566),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_2861),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2705),
.B(n_2462),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_2878),
.B(n_2144),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2538),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2878),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2879),
.B(n_2441),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_2538),
.Y(n_3376)
);

BUFx3_ASAP7_75t_L g3377 ( 
.A(n_2754),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2879),
.B(n_2144),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2538),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2705),
.B(n_2402),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2884),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2884),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2885),
.B(n_2441),
.Y(n_3383)
);

INVx3_ASAP7_75t_L g3384 ( 
.A(n_2754),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2885),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2538),
.Y(n_3386)
);

INVx4_ASAP7_75t_SL g3387 ( 
.A(n_2514),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2540),
.Y(n_3388)
);

INVx4_ASAP7_75t_SL g3389 ( 
.A(n_2957),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3244),
.B(n_2886),
.Y(n_3390)
);

INVx2_ASAP7_75t_SL g3391 ( 
.A(n_3012),
.Y(n_3391)
);

INVx2_ASAP7_75t_SL g3392 ( 
.A(n_3012),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3089),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3305),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3305),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_2952),
.B(n_2336),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_3001),
.Y(n_3397)
);

XOR2xp5_ASAP7_75t_L g3398 ( 
.A(n_3076),
.B(n_1677),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3170),
.B(n_2734),
.Y(n_3399)
);

AND2x6_ASAP7_75t_L g3400 ( 
.A(n_3278),
.B(n_2721),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3309),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3358),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3372),
.Y(n_3403)
);

INVxp33_ASAP7_75t_L g3404 ( 
.A(n_3338),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3372),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_R g3406 ( 
.A(n_3280),
.B(n_2118),
.Y(n_3406)
);

NOR2xp67_ASAP7_75t_L g3407 ( 
.A(n_2990),
.B(n_2212),
.Y(n_3407)
);

NOR2xp67_ASAP7_75t_L g3408 ( 
.A(n_2990),
.B(n_2363),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3378),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3378),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3244),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3245),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3245),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3255),
.Y(n_3414)
);

INVxp33_ASAP7_75t_L g3415 ( 
.A(n_3338),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3255),
.Y(n_3416)
);

BUFx6f_ASAP7_75t_L g3417 ( 
.A(n_3059),
.Y(n_3417)
);

CKINVDCx20_ASAP7_75t_R g3418 ( 
.A(n_2956),
.Y(n_3418)
);

INVx2_ASAP7_75t_SL g3419 ( 
.A(n_3001),
.Y(n_3419)
);

AND2x6_ASAP7_75t_L g3420 ( 
.A(n_3278),
.B(n_3263),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3170),
.B(n_2734),
.Y(n_3421)
);

INVx2_ASAP7_75t_SL g3422 ( 
.A(n_3043),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3256),
.Y(n_3423)
);

INVx2_ASAP7_75t_SL g3424 ( 
.A(n_3043),
.Y(n_3424)
);

XOR2xp5_ASAP7_75t_L g3425 ( 
.A(n_3015),
.B(n_1691),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3256),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3270),
.Y(n_3427)
);

XOR2xp5_ASAP7_75t_L g3428 ( 
.A(n_3061),
.B(n_1721),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3291),
.B(n_2754),
.Y(n_3429)
);

XOR2xp5_ASAP7_75t_L g3430 ( 
.A(n_3109),
.B(n_1721),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3270),
.Y(n_3431)
);

INVxp33_ASAP7_75t_L g3432 ( 
.A(n_2978),
.Y(n_3432)
);

INVx4_ASAP7_75t_SL g3433 ( 
.A(n_2957),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_2926),
.B(n_2470),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3282),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3177),
.B(n_2763),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3282),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_3263),
.B(n_2773),
.Y(n_3438)
);

OAI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3169),
.A2(n_2627),
.B(n_2850),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3288),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3177),
.B(n_2763),
.Y(n_3441)
);

CKINVDCx16_ASAP7_75t_R g3442 ( 
.A(n_3108),
.Y(n_3442)
);

OAI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3275),
.A2(n_2627),
.B(n_2850),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3111),
.B(n_2770),
.Y(n_3444)
);

BUFx6f_ASAP7_75t_L g3445 ( 
.A(n_3059),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3288),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3089),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3322),
.B(n_2470),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3294),
.Y(n_3449)
);

INVx4_ASAP7_75t_SL g3450 ( 
.A(n_2957),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3295),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3295),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3111),
.B(n_2770),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_2982),
.B(n_3030),
.Y(n_3454)
);

XOR2xp5_ASAP7_75t_L g3455 ( 
.A(n_3109),
.B(n_1741),
.Y(n_3455)
);

INVxp67_ASAP7_75t_SL g3456 ( 
.A(n_2920),
.Y(n_3456)
);

INVx2_ASAP7_75t_SL g3457 ( 
.A(n_3280),
.Y(n_3457)
);

NAND2xp33_ASAP7_75t_R g3458 ( 
.A(n_3349),
.B(n_2118),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3298),
.Y(n_3459)
);

CKINVDCx20_ASAP7_75t_R g3460 ( 
.A(n_3073),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3265),
.B(n_2047),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3300),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3300),
.Y(n_3463)
);

INVxp33_ASAP7_75t_L g3464 ( 
.A(n_3126),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3315),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3315),
.Y(n_3466)
);

OR2x2_ASAP7_75t_SL g3467 ( 
.A(n_3162),
.B(n_2916),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3317),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3153),
.B(n_2883),
.Y(n_3469)
);

OR2x2_ASAP7_75t_L g3470 ( 
.A(n_2952),
.B(n_2963),
.Y(n_3470)
);

XOR2xp5_ASAP7_75t_L g3471 ( 
.A(n_3112),
.B(n_1741),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3317),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3318),
.B(n_2886),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3318),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3321),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3321),
.Y(n_3476)
);

AND2x4_ASAP7_75t_L g3477 ( 
.A(n_2933),
.B(n_2784),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_3261),
.B(n_2458),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3325),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3325),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3340),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3340),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3342),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3091),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3342),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3345),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3345),
.Y(n_3487)
);

CKINVDCx20_ASAP7_75t_R g3488 ( 
.A(n_3073),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3364),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3017),
.B(n_2883),
.Y(n_3490)
);

NOR2xp33_ASAP7_75t_L g3491 ( 
.A(n_2953),
.B(n_2458),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3364),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3366),
.Y(n_3493)
);

XOR2x2_ASAP7_75t_L g3494 ( 
.A(n_3055),
.B(n_2135),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3366),
.Y(n_3495)
);

XOR2x2_ASAP7_75t_L g3496 ( 
.A(n_3055),
.B(n_2097),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3374),
.Y(n_3497)
);

BUFx12f_ASAP7_75t_L g3498 ( 
.A(n_3112),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3374),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3017),
.B(n_2489),
.Y(n_3500)
);

CKINVDCx20_ASAP7_75t_R g3501 ( 
.A(n_3164),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3381),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_2973),
.B(n_2468),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3381),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3091),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3382),
.Y(n_3506)
);

CKINVDCx20_ASAP7_75t_R g3507 ( 
.A(n_3164),
.Y(n_3507)
);

NOR2xp33_ASAP7_75t_L g3508 ( 
.A(n_2939),
.B(n_2468),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3093),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3385),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3056),
.B(n_2489),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3385),
.Y(n_3512)
);

CKINVDCx20_ASAP7_75t_R g3513 ( 
.A(n_3349),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3067),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3067),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3082),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3097),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3097),
.Y(n_3518)
);

CKINVDCx20_ASAP7_75t_R g3519 ( 
.A(n_3359),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3082),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3104),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_3359),
.Y(n_3522)
);

INVxp67_ASAP7_75t_L g3523 ( 
.A(n_3174),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3092),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3104),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3113),
.Y(n_3526)
);

INVx1_ASAP7_75t_SL g3527 ( 
.A(n_3102),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3092),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_2919),
.A2(n_2670),
.B(n_2650),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3056),
.B(n_2981),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3095),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3095),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_SL g3533 ( 
.A(n_3049),
.B(n_2363),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3098),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3098),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3100),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3100),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_2918),
.B(n_2887),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_L g3539 ( 
.A(n_3310),
.B(n_2402),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3103),
.Y(n_3540)
);

OAI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3356),
.A2(n_2676),
.B(n_2673),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3103),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3107),
.Y(n_3543)
);

OAI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3166),
.A2(n_2676),
.B(n_2673),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3113),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3107),
.Y(n_3546)
);

AND2x2_ASAP7_75t_SL g3547 ( 
.A(n_3046),
.B(n_2798),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_SL g3548 ( 
.A(n_2982),
.B(n_2773),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3116),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3116),
.Y(n_3550)
);

NOR2xp67_ASAP7_75t_L g3551 ( 
.A(n_3129),
.B(n_2413),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3118),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3118),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3143),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3143),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_3370),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3151),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3151),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_2933),
.B(n_2784),
.Y(n_3559)
);

OAI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3211),
.A2(n_2912),
.B(n_2904),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3158),
.Y(n_3561)
);

INVxp67_ASAP7_75t_SL g3562 ( 
.A(n_2920),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3158),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3161),
.Y(n_3564)
);

CKINVDCx5p33_ASAP7_75t_R g3565 ( 
.A(n_3370),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_L g3566 ( 
.A(n_3355),
.B(n_2611),
.Y(n_3566)
);

NAND2x1p5_ASAP7_75t_L g3567 ( 
.A(n_3269),
.B(n_2773),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3161),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3163),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3163),
.Y(n_3570)
);

XOR2xp5_ASAP7_75t_L g3571 ( 
.A(n_2928),
.B(n_1743),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3165),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3165),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3167),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3371),
.B(n_2611),
.Y(n_3575)
);

BUFx6f_ASAP7_75t_L g3576 ( 
.A(n_3059),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3167),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3168),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3168),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3269),
.B(n_2860),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_2962),
.Y(n_3581)
);

INVxp67_ASAP7_75t_SL g3582 ( 
.A(n_2920),
.Y(n_3582)
);

BUFx6f_ASAP7_75t_L g3583 ( 
.A(n_3115),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3173),
.Y(n_3584)
);

INVx2_ASAP7_75t_SL g3585 ( 
.A(n_3114),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_2984),
.B(n_2489),
.Y(n_3586)
);

XOR2x2_ASAP7_75t_L g3587 ( 
.A(n_3125),
.B(n_2253),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3173),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3176),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3176),
.Y(n_3590)
);

BUFx2_ASAP7_75t_L g3591 ( 
.A(n_2963),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2918),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3019),
.B(n_2503),
.Y(n_3593)
);

XOR2xp5_ASAP7_75t_L g3594 ( 
.A(n_2928),
.B(n_1743),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_2930),
.Y(n_3595)
);

XNOR2xp5_ASAP7_75t_L g3596 ( 
.A(n_2928),
.B(n_1752),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_2936),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2936),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3121),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2940),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2940),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2943),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_2943),
.B(n_2954),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_2954),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_2955),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_2955),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_2958),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_2958),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_2968),
.B(n_2887),
.Y(n_3609)
);

BUFx8_ASAP7_75t_L g3610 ( 
.A(n_3077),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2968),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_2928),
.B(n_2503),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_2976),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2976),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_2979),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_2979),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_2980),
.Y(n_3617)
);

INVxp33_ASAP7_75t_L g3618 ( 
.A(n_3162),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2980),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3121),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3354),
.B(n_2503),
.Y(n_3621)
);

AND2x6_ASAP7_75t_L g3622 ( 
.A(n_3122),
.B(n_2731),
.Y(n_3622)
);

XOR2xp5_ASAP7_75t_L g3623 ( 
.A(n_3207),
.B(n_1752),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3354),
.B(n_2503),
.Y(n_3624)
);

AND2x6_ASAP7_75t_L g3625 ( 
.A(n_3122),
.B(n_2711),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_2985),
.Y(n_3626)
);

AOI21x1_ASAP7_75t_L g3627 ( 
.A1(n_3243),
.A2(n_2853),
.B(n_2900),
.Y(n_3627)
);

INVx1_ASAP7_75t_SL g3628 ( 
.A(n_3205),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_2986),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_2986),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2988),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3303),
.B(n_2513),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_2988),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_2927),
.B(n_2513),
.Y(n_3634)
);

XOR2x2_ASAP7_75t_SL g3635 ( 
.A(n_3080),
.B(n_2389),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3127),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_2999),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_3274),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_2999),
.Y(n_3639)
);

XOR2xp5_ASAP7_75t_L g3640 ( 
.A(n_3207),
.B(n_1755),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3006),
.Y(n_3641)
);

AND2x2_ASAP7_75t_SL g3642 ( 
.A(n_3050),
.B(n_2860),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_3115),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3007),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3007),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3008),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3008),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3127),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3009),
.Y(n_3649)
);

XOR2xp5_ASAP7_75t_L g3650 ( 
.A(n_3241),
.B(n_1755),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3009),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3062),
.B(n_2621),
.Y(n_3652)
);

INVx2_ASAP7_75t_SL g3653 ( 
.A(n_3241),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3011),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3011),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3016),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3016),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3025),
.Y(n_3658)
);

CKINVDCx20_ASAP7_75t_R g3659 ( 
.A(n_3283),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3025),
.B(n_2889),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3029),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3029),
.Y(n_3662)
);

CKINVDCx5p33_ASAP7_75t_R g3663 ( 
.A(n_3077),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3037),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3037),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3038),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3130),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3063),
.B(n_2621),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3038),
.B(n_2889),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3039),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3039),
.Y(n_3671)
);

CKINVDCx20_ASAP7_75t_R g3672 ( 
.A(n_3051),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_2951),
.B(n_2997),
.Y(n_3673)
);

XOR2xp5_ASAP7_75t_L g3674 ( 
.A(n_3052),
.B(n_1773),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3041),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3041),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3045),
.B(n_2513),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3047),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3047),
.Y(n_3679)
);

CKINVDCx20_ASAP7_75t_R g3680 ( 
.A(n_3120),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3057),
.Y(n_3681)
);

OR2x2_ASAP7_75t_L g3682 ( 
.A(n_3078),
.B(n_2336),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3057),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_3077),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3064),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3064),
.Y(n_3686)
);

OAI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_3069),
.A2(n_2912),
.B(n_2904),
.Y(n_3687)
);

INVx1_ASAP7_75t_SL g3688 ( 
.A(n_3005),
.Y(n_3688)
);

XNOR2xp5_ASAP7_75t_L g3689 ( 
.A(n_3052),
.B(n_1773),
.Y(n_3689)
);

INVxp33_ASAP7_75t_SL g3690 ( 
.A(n_3237),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_L g3691 ( 
.A(n_3026),
.B(n_2621),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3065),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3065),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_3247),
.B(n_2621),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3183),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3183),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3184),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3117),
.B(n_2653),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3052),
.B(n_2513),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3052),
.B(n_2653),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3219),
.B(n_3319),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3184),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3187),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3130),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3187),
.Y(n_3705)
);

XOR2x2_ASAP7_75t_L g3706 ( 
.A(n_3125),
.B(n_2381),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3191),
.B(n_2653),
.Y(n_3707)
);

NAND2x1p5_ASAP7_75t_L g3708 ( 
.A(n_3269),
.B(n_2773),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3188),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3188),
.Y(n_3710)
);

XOR2xp5_ASAP7_75t_L g3711 ( 
.A(n_3084),
.B(n_1781),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3219),
.B(n_2653),
.Y(n_3712)
);

CKINVDCx20_ASAP7_75t_R g3713 ( 
.A(n_3252),
.Y(n_3713)
);

OR2x2_ASAP7_75t_L g3714 ( 
.A(n_3197),
.B(n_2111),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3192),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3192),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3319),
.B(n_2870),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3139),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3200),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3060),
.B(n_2870),
.Y(n_3720)
);

NOR2xp67_ASAP7_75t_L g3721 ( 
.A(n_3129),
.B(n_2429),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3200),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3212),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3212),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3213),
.Y(n_3725)
);

CKINVDCx20_ASAP7_75t_R g3726 ( 
.A(n_3115),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_3175),
.A2(n_2125),
.B(n_2605),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_3230),
.B(n_2714),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3213),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_L g3730 ( 
.A(n_3032),
.B(n_2714),
.Y(n_3730)
);

BUFx6f_ASAP7_75t_L g3731 ( 
.A(n_3149),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3214),
.Y(n_3732)
);

BUFx8_ASAP7_75t_L g3733 ( 
.A(n_3131),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3214),
.B(n_2890),
.Y(n_3734)
);

INVxp33_ASAP7_75t_L g3735 ( 
.A(n_3023),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3215),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3060),
.B(n_2870),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3215),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3217),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3217),
.Y(n_3740)
);

NOR2xp33_ASAP7_75t_L g3741 ( 
.A(n_3034),
.B(n_2714),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3222),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3222),
.Y(n_3743)
);

XOR2xp5_ASAP7_75t_L g3744 ( 
.A(n_3125),
.B(n_1781),
.Y(n_3744)
);

BUFx2_ASAP7_75t_L g3745 ( 
.A(n_3004),
.Y(n_3745)
);

XOR2xp5_ASAP7_75t_L g3746 ( 
.A(n_3269),
.B(n_1782),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3223),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3223),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3225),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3225),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3227),
.Y(n_3751)
);

NAND2xp33_ASAP7_75t_R g3752 ( 
.A(n_3004),
.B(n_2130),
.Y(n_3752)
);

INVxp67_ASAP7_75t_SL g3753 ( 
.A(n_2920),
.Y(n_3753)
);

XNOR2x2_ASAP7_75t_L g3754 ( 
.A(n_3311),
.B(n_2467),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3227),
.B(n_2890),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3053),
.B(n_2714),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3228),
.Y(n_3757)
);

XOR2xp5_ASAP7_75t_L g3758 ( 
.A(n_3287),
.B(n_1782),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3228),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3060),
.B(n_2766),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3229),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3229),
.Y(n_3762)
);

INVx4_ASAP7_75t_SL g3763 ( 
.A(n_2957),
.Y(n_3763)
);

INVxp33_ASAP7_75t_L g3764 ( 
.A(n_3178),
.Y(n_3764)
);

INVx1_ASAP7_75t_SL g3765 ( 
.A(n_3287),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3139),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3233),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3233),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3246),
.B(n_2766),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3238),
.Y(n_3770)
);

XOR2xp5_ASAP7_75t_L g3771 ( 
.A(n_3287),
.B(n_1789),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3238),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_3258),
.B(n_2766),
.Y(n_3773)
);

NOR2xp67_ASAP7_75t_L g3774 ( 
.A(n_3132),
.B(n_2429),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3239),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3239),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3587),
.A2(n_2931),
.B1(n_3134),
.B2(n_3131),
.Y(n_3777)
);

AND2x4_ASAP7_75t_L g3778 ( 
.A(n_3580),
.B(n_3287),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3478),
.B(n_2139),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3478),
.B(n_2129),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3393),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3727),
.A2(n_2929),
.B(n_2925),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3461),
.B(n_2766),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3447),
.Y(n_3784)
);

AOI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3706),
.A2(n_3134),
.B1(n_3131),
.B2(n_3181),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3434),
.B(n_2417),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3484),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3394),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3434),
.B(n_2343),
.Y(n_3789)
);

AOI22xp33_ASAP7_75t_L g3790 ( 
.A1(n_3461),
.A2(n_3134),
.B1(n_2779),
.B2(n_2641),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3727),
.A2(n_3058),
.B(n_3193),
.Y(n_3791)
);

INVx5_ASAP7_75t_L g3792 ( 
.A(n_3622),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3503),
.B(n_2343),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3503),
.B(n_3491),
.Y(n_3794)
);

OAI21xp33_ASAP7_75t_L g3795 ( 
.A1(n_3539),
.A2(n_2327),
.B(n_2288),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3539),
.B(n_2343),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3674),
.A2(n_1177),
.B1(n_1180),
.B2(n_1153),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3505),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3509),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3395),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3690),
.B(n_2343),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3530),
.B(n_2867),
.Y(n_3802)
);

NOR3xp33_ASAP7_75t_L g3803 ( 
.A(n_3491),
.B(n_3132),
.C(n_2387),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3399),
.B(n_2867),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_SL g3805 ( 
.A(n_3566),
.B(n_2345),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_R g3806 ( 
.A(n_3406),
.B(n_2295),
.Y(n_3806)
);

BUFx6f_ASAP7_75t_L g3807 ( 
.A(n_3417),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_L g3808 ( 
.A(n_3566),
.B(n_2378),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3575),
.B(n_2345),
.Y(n_3809)
);

BUFx8_ASAP7_75t_L g3810 ( 
.A(n_3498),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3575),
.B(n_2345),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3508),
.B(n_2345),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3581),
.B(n_2345),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3728),
.B(n_2349),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_SL g3815 ( 
.A(n_3728),
.B(n_2349),
.Y(n_3815)
);

INVx2_ASAP7_75t_SL g3816 ( 
.A(n_3610),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_L g3817 ( 
.A1(n_3496),
.A2(n_1186),
.B1(n_1180),
.B2(n_2867),
.Y(n_3817)
);

AOI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3694),
.A2(n_2870),
.B1(n_2867),
.B2(n_2399),
.Y(n_3818)
);

NOR3xp33_ASAP7_75t_L g3819 ( 
.A(n_3698),
.B(n_2399),
.C(n_2387),
.Y(n_3819)
);

OAI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3752),
.A2(n_3698),
.B1(n_2947),
.B2(n_3701),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3401),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3508),
.B(n_2349),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3469),
.B(n_2349),
.Y(n_3823)
);

OAI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3752),
.A2(n_2947),
.B1(n_3171),
.B2(n_3072),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3411),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3444),
.B(n_2349),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3412),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3432),
.B(n_2367),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_3432),
.B(n_2361),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_3726),
.Y(n_3830)
);

INVx2_ASAP7_75t_SL g3831 ( 
.A(n_3610),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3517),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3413),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3464),
.B(n_2361),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_SL g3835 ( 
.A(n_3638),
.B(n_2295),
.Y(n_3835)
);

CKINVDCx5p33_ASAP7_75t_R g3836 ( 
.A(n_3418),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3453),
.B(n_2361),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3490),
.B(n_2361),
.Y(n_3838)
);

OAI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3701),
.A2(n_3171),
.B1(n_3326),
.B2(n_3072),
.Y(n_3839)
);

NOR2xp67_ASAP7_75t_L g3840 ( 
.A(n_3585),
.B(n_2126),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_3687),
.A2(n_3333),
.B(n_3218),
.Y(n_3841)
);

NAND3xp33_ASAP7_75t_L g3842 ( 
.A(n_3694),
.B(n_2361),
.C(n_2404),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_3464),
.B(n_2367),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3396),
.B(n_2360),
.Y(n_3844)
);

O2A1O1Ixp33_ASAP7_75t_L g3845 ( 
.A1(n_3682),
.A2(n_2401),
.B(n_2447),
.C(n_2388),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3414),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3416),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3421),
.B(n_2360),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3423),
.Y(n_3849)
);

OAI221xp5_ASAP7_75t_L g3850 ( 
.A1(n_3448),
.A2(n_2169),
.B1(n_2424),
.B2(n_2425),
.C(n_2418),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3426),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3436),
.B(n_2369),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3441),
.B(n_2369),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3547),
.B(n_3203),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_3691),
.B(n_2371),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3427),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3470),
.B(n_2371),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3431),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3769),
.B(n_2391),
.Y(n_3859)
);

OR2x2_ASAP7_75t_L g3860 ( 
.A(n_3591),
.B(n_2877),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3586),
.B(n_2877),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_3691),
.B(n_2391),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3435),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3769),
.B(n_2392),
.Y(n_3864)
);

O2A1O1Ixp5_ASAP7_75t_L g3865 ( 
.A1(n_3735),
.A2(n_3284),
.B(n_3070),
.C(n_3106),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3518),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3547),
.B(n_3203),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_3688),
.B(n_3367),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3688),
.B(n_3713),
.Y(n_3869)
);

BUFx6f_ASAP7_75t_L g3870 ( 
.A(n_3417),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3521),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3773),
.B(n_2392),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3773),
.B(n_2393),
.Y(n_3873)
);

OAI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3673),
.A2(n_2403),
.B1(n_2406),
.B2(n_2393),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3628),
.B(n_2403),
.Y(n_3875)
);

OR2x6_ASAP7_75t_L g3876 ( 
.A(n_3580),
.B(n_3049),
.Y(n_3876)
);

OR2x6_ASAP7_75t_L g3877 ( 
.A(n_3745),
.B(n_3049),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3618),
.B(n_2406),
.Y(n_3878)
);

NOR2x1p5_ASAP7_75t_L g3879 ( 
.A(n_3556),
.B(n_2111),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3593),
.A2(n_2437),
.B1(n_2438),
.B2(n_2426),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3628),
.B(n_2394),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3527),
.B(n_2443),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3527),
.B(n_2444),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3525),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_SL g3885 ( 
.A(n_3442),
.B(n_2379),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3437),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3440),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3446),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3707),
.B(n_2446),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3449),
.Y(n_3890)
);

NOR2xp33_ASAP7_75t_L g3891 ( 
.A(n_3618),
.B(n_2448),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3673),
.B(n_3329),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3526),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_L g3894 ( 
.A(n_3668),
.B(n_2452),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3687),
.A2(n_3171),
.B(n_3072),
.Y(n_3895)
);

BUFx6f_ASAP7_75t_SL g3896 ( 
.A(n_3391),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3448),
.B(n_2469),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3397),
.B(n_2347),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3451),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3635),
.B(n_3329),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3419),
.B(n_2348),
.Y(n_3901)
);

AOI221xp5_ASAP7_75t_L g3902 ( 
.A1(n_3428),
.A2(n_2237),
.B1(n_2337),
.B2(n_1521),
.C(n_1531),
.Y(n_3902)
);

OAI221xp5_ASAP7_75t_L g3903 ( 
.A1(n_3551),
.A2(n_2120),
.B1(n_2137),
.B2(n_2353),
.C(n_2185),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3422),
.B(n_2370),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3545),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_3632),
.B(n_2982),
.Y(n_3906)
);

NOR2x1p5_ASAP7_75t_L g3907 ( 
.A(n_3565),
.B(n_2213),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3452),
.Y(n_3908)
);

NOR2xp33_ASAP7_75t_SL g3909 ( 
.A(n_3519),
.B(n_2281),
.Y(n_3909)
);

NAND3xp33_ASAP7_75t_L g3910 ( 
.A(n_3406),
.B(n_2063),
.C(n_2049),
.Y(n_3910)
);

INVxp67_ASAP7_75t_SL g3911 ( 
.A(n_3603),
.Y(n_3911)
);

INVx4_ASAP7_75t_L g3912 ( 
.A(n_3389),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3459),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3689),
.A2(n_1186),
.B1(n_2719),
.B2(n_2717),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_SL g3915 ( 
.A(n_3774),
.B(n_2982),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3599),
.Y(n_3916)
);

NOR3xp33_ASAP7_75t_L g3917 ( 
.A(n_3730),
.B(n_3330),
.C(n_3312),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3424),
.B(n_2370),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3668),
.B(n_2082),
.Y(n_3919)
);

NOR3xp33_ASAP7_75t_L g3920 ( 
.A(n_3730),
.B(n_3362),
.C(n_2453),
.Y(n_3920)
);

NOR3xp33_ASAP7_75t_L g3921 ( 
.A(n_3741),
.B(n_3380),
.C(n_2696),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_3652),
.B(n_2090),
.Y(n_3922)
);

AOI22xp33_ASAP7_75t_L g3923 ( 
.A1(n_3744),
.A2(n_2717),
.B1(n_2724),
.B2(n_2719),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3620),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3636),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3402),
.B(n_2373),
.Y(n_3926)
);

NOR2xp33_ASAP7_75t_L g3927 ( 
.A(n_3652),
.B(n_2281),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3648),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3462),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3403),
.B(n_2375),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3667),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3704),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3405),
.B(n_2375),
.Y(n_3933)
);

INVx3_ASAP7_75t_L g3934 ( 
.A(n_3567),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3463),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3672),
.B(n_1789),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3712),
.B(n_3717),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3389),
.B(n_2982),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3389),
.B(n_2982),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3409),
.B(n_2376),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3410),
.B(n_2376),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3718),
.Y(n_3942)
);

AOI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_3494),
.A2(n_2319),
.B1(n_1793),
.B2(n_1811),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3523),
.B(n_3285),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_L g3945 ( 
.A(n_3417),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_SL g3946 ( 
.A(n_3433),
.B(n_3450),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3766),
.Y(n_3947)
);

AOI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3458),
.A2(n_2319),
.B1(n_1793),
.B2(n_1811),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3523),
.B(n_3293),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3500),
.B(n_3511),
.Y(n_3950)
);

AOI22xp5_ASAP7_75t_L g3951 ( 
.A1(n_3458),
.A2(n_1833),
.B1(n_1840),
.B2(n_1792),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3514),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3465),
.Y(n_3953)
);

NAND3xp33_ASAP7_75t_L g3954 ( 
.A(n_3741),
.B(n_2063),
.C(n_2049),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_SL g3955 ( 
.A(n_3433),
.B(n_3030),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3634),
.B(n_3301),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3466),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_L g3958 ( 
.A(n_3621),
.B(n_2880),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3677),
.B(n_3327),
.Y(n_3959)
);

OR2x6_ASAP7_75t_L g3960 ( 
.A(n_3477),
.B(n_3049),
.Y(n_3960)
);

BUFx6f_ASAP7_75t_SL g3961 ( 
.A(n_3392),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3515),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3624),
.B(n_3328),
.Y(n_3963)
);

BUFx6f_ASAP7_75t_SL g3964 ( 
.A(n_3457),
.Y(n_3964)
);

INVx3_ASAP7_75t_L g3965 ( 
.A(n_3567),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3516),
.Y(n_3966)
);

INVx3_ASAP7_75t_L g3967 ( 
.A(n_3708),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3520),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3433),
.B(n_3030),
.Y(n_3969)
);

OAI221xp5_ASAP7_75t_L g3970 ( 
.A1(n_3721),
.A2(n_2433),
.B1(n_2352),
.B2(n_2362),
.C(n_2354),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3450),
.B(n_3030),
.Y(n_3971)
);

NAND2x1_ASAP7_75t_L g3972 ( 
.A(n_3445),
.B(n_3341),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_3735),
.B(n_2888),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3612),
.B(n_2394),
.Y(n_3974)
);

BUFx3_ASAP7_75t_L g3975 ( 
.A(n_3460),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3571),
.A2(n_2725),
.B1(n_2735),
.B2(n_2724),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3700),
.B(n_2394),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3468),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3603),
.B(n_3361),
.Y(n_3979)
);

CKINVDCx5p33_ASAP7_75t_R g3980 ( 
.A(n_3522),
.Y(n_3980)
);

NOR2xp33_ASAP7_75t_L g3981 ( 
.A(n_3764),
.B(n_3004),
.Y(n_3981)
);

BUFx6f_ASAP7_75t_L g3982 ( 
.A(n_3445),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3472),
.B(n_3375),
.Y(n_3983)
);

BUFx6f_ASAP7_75t_SL g3984 ( 
.A(n_3653),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3594),
.A2(n_2735),
.B1(n_2744),
.B2(n_2725),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3404),
.B(n_2398),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3450),
.B(n_3763),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3474),
.B(n_3383),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3404),
.B(n_2398),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3746),
.B(n_2398),
.Y(n_3990)
);

O2A1O1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3756),
.A2(n_2785),
.B(n_2911),
.C(n_2651),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3475),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3415),
.B(n_2405),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3415),
.B(n_2405),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3476),
.Y(n_3995)
);

AOI22xp5_ASAP7_75t_L g3996 ( 
.A1(n_3680),
.A2(n_1833),
.B1(n_1840),
.B2(n_1792),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_L g3997 ( 
.A(n_3765),
.B(n_3004),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3479),
.Y(n_3998)
);

HB1xp67_ASAP7_75t_SL g3999 ( 
.A(n_3733),
.Y(n_3999)
);

INVx5_ASAP7_75t_L g4000 ( 
.A(n_3622),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3480),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3524),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3481),
.B(n_2337),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_3763),
.B(n_3030),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3482),
.B(n_2337),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3528),
.Y(n_4006)
);

OAI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_3390),
.A2(n_3072),
.B1(n_3326),
.B2(n_3171),
.Y(n_4007)
);

HB1xp67_ASAP7_75t_L g4008 ( 
.A(n_3456),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3483),
.B(n_2167),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3765),
.B(n_3004),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3485),
.B(n_2167),
.Y(n_4011)
);

NOR2xp33_ASAP7_75t_L g4012 ( 
.A(n_3659),
.B(n_2130),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3486),
.Y(n_4013)
);

OR2x6_ASAP7_75t_L g4014 ( 
.A(n_3477),
.B(n_3049),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3763),
.B(n_3030),
.Y(n_4015)
);

INVx2_ASAP7_75t_SL g4016 ( 
.A(n_3733),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3531),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3487),
.B(n_2152),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_SL g4019 ( 
.A(n_3445),
.B(n_3159),
.Y(n_4019)
);

OR2x2_ASAP7_75t_L g4020 ( 
.A(n_3758),
.B(n_2213),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3489),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3576),
.B(n_3583),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3532),
.Y(n_4023)
);

NOR3xp33_ASAP7_75t_L g4024 ( 
.A(n_3756),
.B(n_3150),
.C(n_2946),
.Y(n_4024)
);

AOI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3425),
.A2(n_1846),
.B1(n_1843),
.B2(n_2166),
.Y(n_4025)
);

A2O1A1Ixp33_ASAP7_75t_L g4026 ( 
.A1(n_3560),
.A2(n_3135),
.B(n_3186),
.C(n_3090),
.Y(n_4026)
);

NOR2xp33_ASAP7_75t_L g4027 ( 
.A(n_3771),
.B(n_3060),
.Y(n_4027)
);

NOR2xp67_ASAP7_75t_L g4028 ( 
.A(n_3408),
.B(n_2899),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3534),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3492),
.B(n_2152),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3493),
.B(n_2152),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_R g4032 ( 
.A(n_3501),
.B(n_2173),
.Y(n_4032)
);

BUFx6f_ASAP7_75t_L g4033 ( 
.A(n_3576),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_SL g4034 ( 
.A(n_3576),
.B(n_3159),
.Y(n_4034)
);

NOR3xp33_ASAP7_75t_L g4035 ( 
.A(n_3560),
.B(n_2987),
.C(n_2977),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3720),
.B(n_3138),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_L g4037 ( 
.A(n_3737),
.B(n_3138),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3495),
.Y(n_4038)
);

AOI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3430),
.A2(n_1846),
.B1(n_1843),
.B2(n_2166),
.Y(n_4039)
);

BUFx6f_ASAP7_75t_L g4040 ( 
.A(n_3583),
.Y(n_4040)
);

AOI22xp33_ASAP7_75t_L g4041 ( 
.A1(n_3711),
.A2(n_2745),
.B1(n_2747),
.B2(n_2744),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3535),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3497),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3583),
.B(n_3159),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3536),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3499),
.Y(n_4046)
);

OAI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3390),
.A2(n_3171),
.B1(n_3326),
.B2(n_3072),
.Y(n_4047)
);

BUFx6f_ASAP7_75t_L g4048 ( 
.A(n_3643),
.Y(n_4048)
);

INVx3_ASAP7_75t_L g4049 ( 
.A(n_3708),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3760),
.B(n_3455),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3502),
.B(n_2167),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3537),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3504),
.B(n_3506),
.Y(n_4053)
);

OAI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3529),
.A2(n_2691),
.B(n_2675),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3510),
.B(n_2172),
.Y(n_4055)
);

NOR3x1_ASAP7_75t_L g4056 ( 
.A(n_3714),
.B(n_2420),
.C(n_2178),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3512),
.B(n_2172),
.Y(n_4057)
);

AO221x1_ASAP7_75t_L g4058 ( 
.A1(n_3731),
.A2(n_3368),
.B1(n_3066),
.B2(n_3140),
.C(n_2975),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3731),
.B(n_3159),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_3731),
.B(n_3235),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_SL g4061 ( 
.A(n_3533),
.B(n_3235),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3592),
.B(n_3595),
.Y(n_4062)
);

A2O1A1Ixp33_ASAP7_75t_L g4063 ( 
.A1(n_3473),
.A2(n_3135),
.B(n_3096),
.C(n_3099),
.Y(n_4063)
);

INVxp67_ASAP7_75t_L g4064 ( 
.A(n_3559),
.Y(n_4064)
);

NOR2xp67_ASAP7_75t_L g4065 ( 
.A(n_3407),
.B(n_2905),
.Y(n_4065)
);

INVxp67_ASAP7_75t_L g4066 ( 
.A(n_3559),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_SL g4067 ( 
.A(n_3533),
.B(n_3235),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3473),
.B(n_3235),
.Y(n_4068)
);

INVx3_ASAP7_75t_L g4069 ( 
.A(n_3622),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3540),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3542),
.Y(n_4071)
);

NOR2xp33_ASAP7_75t_L g4072 ( 
.A(n_3471),
.B(n_3138),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3699),
.B(n_2217),
.Y(n_4073)
);

NOR2xp67_ASAP7_75t_L g4074 ( 
.A(n_3663),
.B(n_3299),
.Y(n_4074)
);

INVxp67_ASAP7_75t_L g4075 ( 
.A(n_3754),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3543),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3597),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3538),
.B(n_3235),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3546),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3549),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3550),
.Y(n_4081)
);

NOR2xp67_ASAP7_75t_L g4082 ( 
.A(n_3684),
.B(n_3299),
.Y(n_4082)
);

INVx2_ASAP7_75t_SL g4083 ( 
.A(n_3507),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3598),
.B(n_2049),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_SL g4085 ( 
.A(n_3538),
.B(n_3235),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3623),
.B(n_2278),
.Y(n_4086)
);

O2A1O1Ixp5_ASAP7_75t_L g4087 ( 
.A1(n_3429),
.A2(n_3081),
.B(n_3124),
.C(n_3123),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3552),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_3596),
.A2(n_2747),
.B1(n_2751),
.B2(n_2745),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3600),
.B(n_2063),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3601),
.B(n_2064),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3640),
.B(n_2058),
.Y(n_4092)
);

NOR2xp33_ASAP7_75t_L g4093 ( 
.A(n_3650),
.B(n_3138),
.Y(n_4093)
);

AOI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3513),
.A2(n_2178),
.B1(n_2420),
.B2(n_2280),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_3642),
.B(n_3189),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3553),
.Y(n_4096)
);

AOI22xp5_ASAP7_75t_L g4097 ( 
.A1(n_3398),
.A2(n_2280),
.B1(n_2289),
.B2(n_2064),
.Y(n_4097)
);

INVx2_ASAP7_75t_SL g4098 ( 
.A(n_3488),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3602),
.B(n_2064),
.Y(n_4099)
);

AND2x4_ASAP7_75t_L g4100 ( 
.A(n_3604),
.B(n_3149),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3605),
.B(n_2280),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3554),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3606),
.B(n_2289),
.Y(n_4103)
);

NAND3xp33_ASAP7_75t_L g4104 ( 
.A(n_3609),
.B(n_2298),
.C(n_2289),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_3642),
.B(n_3189),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_3420),
.A2(n_2755),
.B1(n_2800),
.B2(n_2751),
.Y(n_4106)
);

INVx2_ASAP7_75t_SL g4107 ( 
.A(n_3607),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3608),
.Y(n_4108)
);

O2A1O1Ixp5_ASAP7_75t_L g4109 ( 
.A1(n_3429),
.A2(n_3136),
.B(n_3208),
.C(n_3201),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_3555),
.Y(n_4110)
);

INVx2_ASAP7_75t_SL g4111 ( 
.A(n_3611),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3557),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3613),
.B(n_2298),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3614),
.B(n_3615),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_SL g4115 ( 
.A(n_3609),
.B(n_3248),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_L g4116 ( 
.A(n_3660),
.B(n_3189),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3622),
.Y(n_4117)
);

INVxp67_ASAP7_75t_L g4118 ( 
.A(n_3616),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3617),
.B(n_2298),
.Y(n_4119)
);

OAI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_3529),
.A2(n_2720),
.B(n_2703),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3619),
.B(n_2350),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_SL g4122 ( 
.A(n_3660),
.B(n_3248),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3626),
.Y(n_4123)
);

NOR2xp33_ASAP7_75t_L g4124 ( 
.A(n_3669),
.B(n_3189),
.Y(n_4124)
);

AOI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3420),
.A2(n_2800),
.B1(n_2802),
.B2(n_2755),
.Y(n_4125)
);

A2O1A1Ixp33_ASAP7_75t_L g4126 ( 
.A1(n_3669),
.A2(n_3101),
.B(n_3105),
.C(n_3085),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_3467),
.B(n_3250),
.Y(n_4127)
);

AND2x4_ASAP7_75t_SL g4128 ( 
.A(n_3629),
.B(n_2923),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_3630),
.B(n_2350),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3631),
.B(n_2891),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3633),
.B(n_3637),
.Y(n_4131)
);

NAND2x1_ASAP7_75t_L g4132 ( 
.A(n_3558),
.B(n_3341),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3639),
.B(n_2891),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3641),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3644),
.B(n_2893),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3645),
.B(n_2897),
.Y(n_4136)
);

OAI22xp5_ASAP7_75t_SL g4137 ( 
.A1(n_3646),
.A2(n_2173),
.B1(n_1872),
.B2(n_1893),
.Y(n_4137)
);

INVx6_ASAP7_75t_L g4138 ( 
.A(n_3778),
.Y(n_4138)
);

AOI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_3808),
.A2(n_3326),
.B1(n_2957),
.B2(n_3420),
.Y(n_4139)
);

INVx1_ASAP7_75t_SL g4140 ( 
.A(n_4032),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_SL g4141 ( 
.A1(n_3808),
.A2(n_1872),
.B1(n_1893),
.B2(n_1867),
.Y(n_4141)
);

AND2x4_ASAP7_75t_L g4142 ( 
.A(n_3778),
.B(n_3960),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3781),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_3797),
.A2(n_1905),
.B1(n_1867),
.B2(n_2180),
.Y(n_4144)
);

NOR3xp33_ASAP7_75t_L g4145 ( 
.A(n_3795),
.B(n_2534),
.C(n_2533),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3911),
.B(n_3647),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3952),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3962),
.Y(n_4148)
);

BUFx3_ASAP7_75t_L g4149 ( 
.A(n_3830),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_3807),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3911),
.B(n_3649),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_3784),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3794),
.B(n_3651),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3979),
.B(n_3654),
.Y(n_4154)
);

HB1xp67_ASAP7_75t_L g4155 ( 
.A(n_4107),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3966),
.Y(n_4156)
);

INVx2_ASAP7_75t_SL g4157 ( 
.A(n_3879),
.Y(n_4157)
);

INVx2_ASAP7_75t_SL g4158 ( 
.A(n_3907),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3968),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4002),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4006),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_SL g4162 ( 
.A(n_3855),
.B(n_3250),
.Y(n_4162)
);

HB1xp67_ASAP7_75t_L g4163 ( 
.A(n_4111),
.Y(n_4163)
);

BUFx12f_ASAP7_75t_L g4164 ( 
.A(n_3836),
.Y(n_4164)
);

NAND2x1p5_ASAP7_75t_L g4165 ( 
.A(n_3912),
.B(n_3248),
.Y(n_4165)
);

INVx2_ASAP7_75t_SL g4166 ( 
.A(n_3975),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4017),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4023),
.Y(n_4168)
);

INVx1_ASAP7_75t_SL g4169 ( 
.A(n_3806),
.Y(n_4169)
);

AND2x4_ASAP7_75t_L g4170 ( 
.A(n_3960),
.B(n_3655),
.Y(n_4170)
);

INVx1_ASAP7_75t_SL g4171 ( 
.A(n_3835),
.Y(n_4171)
);

NOR3xp33_ASAP7_75t_SL g4172 ( 
.A(n_3980),
.B(n_1521),
.C(n_1519),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4029),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4042),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4045),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4052),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3787),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4070),
.Y(n_4178)
);

INVxp67_ASAP7_75t_L g4179 ( 
.A(n_3936),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4075),
.B(n_3656),
.Y(n_4180)
);

INVx2_ASAP7_75t_SL g4181 ( 
.A(n_3816),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_SL g4182 ( 
.A(n_3862),
.B(n_3142),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_3797),
.A2(n_1905),
.B1(n_2201),
.B2(n_2180),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3798),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4071),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_R g4186 ( 
.A(n_3999),
.B(n_2386),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_3799),
.Y(n_4187)
);

BUFx2_ASAP7_75t_L g4188 ( 
.A(n_3807),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4076),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4075),
.B(n_3657),
.Y(n_4190)
);

BUFx6f_ASAP7_75t_L g4191 ( 
.A(n_3807),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_3869),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3819),
.B(n_3894),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_3809),
.B(n_3155),
.Y(n_4194)
);

HB1xp67_ASAP7_75t_L g4195 ( 
.A(n_4008),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_3960),
.B(n_3658),
.Y(n_4196)
);

BUFx3_ASAP7_75t_L g4197 ( 
.A(n_3810),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_3789),
.B(n_2920),
.Y(n_4198)
);

O2A1O1Ixp33_ASAP7_75t_L g4199 ( 
.A1(n_3779),
.A2(n_3020),
.B(n_2991),
.C(n_678),
.Y(n_4199)
);

INVx3_ASAP7_75t_L g4200 ( 
.A(n_3912),
.Y(n_4200)
);

NOR3xp33_ASAP7_75t_SL g4201 ( 
.A(n_3850),
.B(n_1531),
.C(n_1528),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3894),
.B(n_3661),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_SL g4203 ( 
.A(n_3927),
.B(n_3786),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4079),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4116),
.B(n_4124),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4080),
.Y(n_4206)
);

OR2x6_ASAP7_75t_L g4207 ( 
.A(n_4014),
.B(n_3438),
.Y(n_4207)
);

BUFx12f_ASAP7_75t_L g4208 ( 
.A(n_3810),
.Y(n_4208)
);

NAND3xp33_ASAP7_75t_SL g4209 ( 
.A(n_3780),
.B(n_712),
.C(n_685),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4116),
.B(n_3662),
.Y(n_4210)
);

CKINVDCx5p33_ASAP7_75t_R g4211 ( 
.A(n_3999),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_3914),
.A2(n_2180),
.B1(n_2209),
.B2(n_2201),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4124),
.B(n_3664),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4081),
.Y(n_4214)
);

AOI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_3914),
.A2(n_2201),
.B1(n_2209),
.B2(n_2998),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4088),
.Y(n_4216)
);

AND2x6_ASAP7_75t_L g4217 ( 
.A(n_4069),
.B(n_3665),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_3832),
.Y(n_4218)
);

OR2x6_ASAP7_75t_L g4219 ( 
.A(n_4014),
.B(n_3438),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4096),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_4118),
.B(n_3666),
.Y(n_4221)
);

INVx3_ASAP7_75t_L g4222 ( 
.A(n_3807),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4118),
.B(n_3670),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_3802),
.B(n_712),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3866),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_3793),
.B(n_2975),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_4014),
.B(n_3671),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_3871),
.Y(n_4228)
);

BUFx2_ASAP7_75t_L g4229 ( 
.A(n_3870),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4102),
.Y(n_4230)
);

BUFx3_ASAP7_75t_L g4231 ( 
.A(n_3831),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4110),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_3963),
.B(n_3675),
.Y(n_4233)
);

AND2x4_ASAP7_75t_L g4234 ( 
.A(n_3876),
.B(n_3676),
.Y(n_4234)
);

AOI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3900),
.A2(n_3922),
.B1(n_3919),
.B2(n_3783),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3859),
.B(n_3678),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3864),
.B(n_3679),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_3804),
.B(n_745),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3872),
.B(n_3681),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_3870),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3884),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4112),
.Y(n_4242)
);

AOI211xp5_ASAP7_75t_L g4243 ( 
.A1(n_3903),
.A2(n_3902),
.B(n_3922),
.C(n_3842),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_3825),
.Y(n_4244)
);

AOI22xp33_ASAP7_75t_L g4245 ( 
.A1(n_3817),
.A2(n_2209),
.B1(n_3010),
.B2(n_2810),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_3873),
.B(n_3683),
.Y(n_4246)
);

AOI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_3919),
.A2(n_2058),
.B1(n_1541),
.B2(n_1546),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_3812),
.B(n_2975),
.Y(n_4248)
);

AO21x1_ASAP7_75t_L g4249 ( 
.A1(n_3820),
.A2(n_3232),
.B(n_3231),
.Y(n_4249)
);

INVx2_ASAP7_75t_SL g4250 ( 
.A(n_4016),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3893),
.Y(n_4251)
);

AND2x2_ASAP7_75t_L g4252 ( 
.A(n_3861),
.B(n_745),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3827),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3822),
.B(n_3685),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3833),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_3905),
.Y(n_4256)
);

OR2x4_ASAP7_75t_L g4257 ( 
.A(n_3828),
.B(n_3561),
.Y(n_4257)
);

HB1xp67_ASAP7_75t_L g4258 ( 
.A(n_3860),
.Y(n_4258)
);

NOR2xp33_ASAP7_75t_L g4259 ( 
.A(n_4012),
.B(n_1533),
.Y(n_4259)
);

BUFx12f_ASAP7_75t_L g4260 ( 
.A(n_4083),
.Y(n_4260)
);

AO22x1_ASAP7_75t_L g4261 ( 
.A1(n_4056),
.A2(n_3341),
.B1(n_916),
.B2(n_954),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3846),
.B(n_3686),
.Y(n_4262)
);

NAND2x1p5_ASAP7_75t_L g4263 ( 
.A(n_3946),
.B(n_3248),
.Y(n_4263)
);

INVx8_ASAP7_75t_L g4264 ( 
.A(n_3876),
.Y(n_4264)
);

NAND2x1p5_ASAP7_75t_L g4265 ( 
.A(n_3987),
.B(n_3248),
.Y(n_4265)
);

NOR2xp33_ASAP7_75t_L g4266 ( 
.A(n_4012),
.B(n_1533),
.Y(n_4266)
);

INVx5_ASAP7_75t_L g4267 ( 
.A(n_3876),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3847),
.B(n_3692),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3849),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_3916),
.Y(n_4270)
);

INVx3_ASAP7_75t_L g4271 ( 
.A(n_3870),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3851),
.B(n_3693),
.Y(n_4272)
);

CKINVDCx5p33_ASAP7_75t_R g4273 ( 
.A(n_3964),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3856),
.Y(n_4274)
);

AO22x1_ASAP7_75t_L g4275 ( 
.A1(n_4093),
.A2(n_3341),
.B1(n_916),
.B2(n_954),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_3858),
.B(n_3863),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3886),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3887),
.Y(n_4278)
);

AOI21xp5_ASAP7_75t_L g4279 ( 
.A1(n_3841),
.A2(n_3541),
.B(n_3544),
.Y(n_4279)
);

HB1xp67_ASAP7_75t_L g4280 ( 
.A(n_4100),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_SL g4281 ( 
.A(n_3790),
.B(n_2975),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3888),
.Y(n_4282)
);

AOI22xp33_ASAP7_75t_L g4283 ( 
.A1(n_3817),
.A2(n_2810),
.B1(n_2813),
.B2(n_2802),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_3924),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3890),
.B(n_3772),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3899),
.Y(n_4286)
);

OAI22xp5_ASAP7_75t_SL g4287 ( 
.A1(n_4039),
.A2(n_751),
.B1(n_804),
.B2(n_763),
.Y(n_4287)
);

NOR2x2_ASAP7_75t_L g4288 ( 
.A(n_3885),
.B(n_2923),
.Y(n_4288)
);

OAI22xp33_ASAP7_75t_L g4289 ( 
.A1(n_3818),
.A2(n_2923),
.B1(n_2736),
.B2(n_2827),
.Y(n_4289)
);

AOI22xp33_ASAP7_75t_L g4290 ( 
.A1(n_3777),
.A2(n_2814),
.B1(n_2816),
.B2(n_2813),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_3986),
.B(n_751),
.Y(n_4291)
);

OR2x6_ASAP7_75t_L g4292 ( 
.A(n_3877),
.B(n_2923),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3908),
.Y(n_4293)
);

A2O1A1Ixp33_ASAP7_75t_L g4294 ( 
.A1(n_3845),
.A2(n_2898),
.B(n_2897),
.C(n_3734),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_3925),
.Y(n_4295)
);

INVx4_ASAP7_75t_L g4296 ( 
.A(n_3964),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3913),
.Y(n_4297)
);

A2O1A1Ixp33_ASAP7_75t_L g4298 ( 
.A1(n_3803),
.A2(n_2898),
.B(n_3734),
.C(n_3755),
.Y(n_4298)
);

INVx4_ASAP7_75t_L g4299 ( 
.A(n_3896),
.Y(n_4299)
);

NAND2x1p5_ASAP7_75t_L g4300 ( 
.A(n_3792),
.B(n_3248),
.Y(n_4300)
);

NOR2xp67_ASAP7_75t_L g4301 ( 
.A(n_3910),
.B(n_3260),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_3989),
.B(n_3993),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3929),
.B(n_3757),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3935),
.Y(n_4304)
);

AND2x4_ASAP7_75t_L g4305 ( 
.A(n_4064),
.B(n_3563),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_3953),
.B(n_3759),
.Y(n_4306)
);

BUFx6f_ASAP7_75t_L g4307 ( 
.A(n_3870),
.Y(n_4307)
);

CKINVDCx20_ASAP7_75t_R g4308 ( 
.A(n_3996),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3957),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_3978),
.B(n_3761),
.Y(n_4310)
);

INVx1_ASAP7_75t_SL g4311 ( 
.A(n_4098),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_3928),
.Y(n_4312)
);

INVxp67_ASAP7_75t_L g4313 ( 
.A(n_3828),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3992),
.B(n_3995),
.Y(n_4314)
);

AOI22xp33_ASAP7_75t_L g4315 ( 
.A1(n_3777),
.A2(n_2816),
.B1(n_2820),
.B2(n_2814),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_3788),
.Y(n_4316)
);

CKINVDCx5p33_ASAP7_75t_R g4317 ( 
.A(n_3896),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_SL g4318 ( 
.A(n_3790),
.B(n_2975),
.Y(n_4318)
);

OR2x6_ASAP7_75t_L g4319 ( 
.A(n_3877),
.B(n_2923),
.Y(n_4319)
);

AND2x4_ASAP7_75t_L g4320 ( 
.A(n_4064),
.B(n_3564),
.Y(n_4320)
);

NOR2x2_ASAP7_75t_L g4321 ( 
.A(n_3909),
.B(n_2294),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_3800),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_3931),
.Y(n_4323)
);

INVx5_ASAP7_75t_L g4324 ( 
.A(n_3877),
.Y(n_4324)
);

OR2x6_ASAP7_75t_L g4325 ( 
.A(n_3895),
.B(n_3755),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_3998),
.B(n_3740),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_3932),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_3857),
.B(n_3568),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4001),
.B(n_3743),
.Y(n_4329)
);

AOI22xp5_ASAP7_75t_L g4330 ( 
.A1(n_3973),
.A2(n_1548),
.B1(n_1550),
.B2(n_1541),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4013),
.B(n_3748),
.Y(n_4331)
);

INVx1_ASAP7_75t_SL g4332 ( 
.A(n_3882),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4021),
.B(n_3749),
.Y(n_4333)
);

OAI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_3990),
.A2(n_763),
.B1(n_836),
.B2(n_804),
.Y(n_4334)
);

INVx3_ASAP7_75t_L g4335 ( 
.A(n_3945),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_SL g4336 ( 
.A(n_3803),
.B(n_3066),
.Y(n_4336)
);

NOR2x1_ASAP7_75t_L g4337 ( 
.A(n_3813),
.B(n_3286),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4038),
.B(n_3762),
.Y(n_4338)
);

AOI22xp33_ASAP7_75t_L g4339 ( 
.A1(n_3923),
.A2(n_2821),
.B1(n_2822),
.B2(n_2820),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_3942),
.Y(n_4340)
);

BUFx6f_ASAP7_75t_L g4341 ( 
.A(n_3945),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_SL g4342 ( 
.A(n_3823),
.B(n_3066),
.Y(n_4342)
);

NOR2xp33_ASAP7_75t_L g4343 ( 
.A(n_4025),
.B(n_1548),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4043),
.Y(n_4344)
);

BUFx3_ASAP7_75t_L g4345 ( 
.A(n_3945),
.Y(n_4345)
);

INVx4_ASAP7_75t_L g4346 ( 
.A(n_3961),
.Y(n_4346)
);

OAI22xp5_ASAP7_75t_SL g4347 ( 
.A1(n_4094),
.A2(n_836),
.B1(n_858),
.B2(n_846),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_SL g4348 ( 
.A(n_3854),
.B(n_3066),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_3947),
.Y(n_4349)
);

NOR2x1p5_ASAP7_75t_L g4350 ( 
.A(n_4104),
.B(n_3149),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4046),
.Y(n_4351)
);

BUFx12f_ASAP7_75t_L g4352 ( 
.A(n_4020),
.Y(n_4352)
);

BUFx2_ASAP7_75t_L g4353 ( 
.A(n_3982),
.Y(n_4353)
);

BUFx6f_ASAP7_75t_L g4354 ( 
.A(n_3982),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_3867),
.B(n_3066),
.Y(n_4355)
);

BUFx6f_ASAP7_75t_SL g4356 ( 
.A(n_3982),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4077),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_3951),
.B(n_1550),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4108),
.B(n_3729),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4123),
.Y(n_4360)
);

INVx3_ASAP7_75t_SL g4361 ( 
.A(n_3881),
.Y(n_4361)
);

CKINVDCx8_ASAP7_75t_R g4362 ( 
.A(n_3982),
.Y(n_4362)
);

OAI22xp33_ASAP7_75t_L g4363 ( 
.A1(n_3880),
.A2(n_846),
.B1(n_1053),
.B2(n_858),
.Y(n_4363)
);

OAI21xp33_ASAP7_75t_SL g4364 ( 
.A1(n_4058),
.A2(n_3811),
.B(n_3805),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_3961),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_3948),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4134),
.B(n_3738),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_L g4368 ( 
.A(n_3943),
.B(n_3973),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_4066),
.B(n_3569),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3821),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_3981),
.A2(n_1565),
.B1(n_1567),
.B2(n_1562),
.Y(n_4371)
);

OAI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4106),
.A2(n_3747),
.B1(n_3750),
.B2(n_3742),
.Y(n_4372)
);

BUFx6f_ASAP7_75t_L g4373 ( 
.A(n_4033),
.Y(n_4373)
);

INVx3_ASAP7_75t_L g4374 ( 
.A(n_4033),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_3983),
.B(n_3751),
.Y(n_4375)
);

INVx6_ASAP7_75t_L g4376 ( 
.A(n_4033),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3988),
.B(n_3767),
.Y(n_4377)
);

NOR2xp33_ASAP7_75t_L g4378 ( 
.A(n_3891),
.B(n_1562),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4053),
.B(n_3768),
.Y(n_4379)
);

HB1xp67_ASAP7_75t_L g4380 ( 
.A(n_4033),
.Y(n_4380)
);

INVx3_ASAP7_75t_L g4381 ( 
.A(n_4040),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_3984),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4062),
.Y(n_4383)
);

INVx4_ASAP7_75t_L g4384 ( 
.A(n_3984),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4114),
.Y(n_4385)
);

CKINVDCx5p33_ASAP7_75t_R g4386 ( 
.A(n_4137),
.Y(n_4386)
);

AO22x1_ASAP7_75t_L g4387 ( 
.A1(n_4093),
.A2(n_1105),
.B1(n_1160),
.B2(n_1053),
.Y(n_4387)
);

NOR2xp33_ASAP7_75t_L g4388 ( 
.A(n_3891),
.B(n_1565),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_4040),
.Y(n_4389)
);

INVx3_ASAP7_75t_L g4390 ( 
.A(n_4040),
.Y(n_4390)
);

NOR2xp33_ASAP7_75t_L g4391 ( 
.A(n_3843),
.B(n_1567),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4131),
.B(n_3570),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4130),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_3956),
.B(n_3710),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_3994),
.B(n_1105),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_3791),
.A2(n_3541),
.B(n_3544),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_SL g4397 ( 
.A1(n_3792),
.A2(n_3622),
.B1(n_3625),
.B2(n_3400),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4133),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4135),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4136),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_SL g4401 ( 
.A(n_3897),
.B(n_3140),
.Y(n_4401)
);

CKINVDCx14_ASAP7_75t_R g4402 ( 
.A(n_4097),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3944),
.Y(n_4403)
);

NOR2xp33_ASAP7_75t_L g4404 ( 
.A(n_3843),
.B(n_1568),
.Y(n_4404)
);

BUFx3_ASAP7_75t_L g4405 ( 
.A(n_4048),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_SL g4406 ( 
.A(n_3820),
.B(n_3140),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_3814),
.B(n_3140),
.Y(n_4407)
);

OAI221xp5_ASAP7_75t_L g4408 ( 
.A1(n_3874),
.A2(n_1160),
.B1(n_807),
.B2(n_810),
.C(n_809),
.Y(n_4408)
);

INVx2_ASAP7_75t_SL g4409 ( 
.A(n_4048),
.Y(n_4409)
);

NAND2x2_ASAP7_75t_L g4410 ( 
.A(n_3838),
.B(n_3220),
.Y(n_4410)
);

INVx5_ASAP7_75t_L g4411 ( 
.A(n_3792),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_3958),
.B(n_748),
.Y(n_4412)
);

INVxp67_ASAP7_75t_SL g4413 ( 
.A(n_3997),
.Y(n_4413)
);

HB1xp67_ASAP7_75t_L g4414 ( 
.A(n_4048),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4106),
.A2(n_3732),
.B1(n_3736),
.B2(n_3725),
.Y(n_4415)
);

BUFx6f_ASAP7_75t_L g4416 ( 
.A(n_4048),
.Y(n_4416)
);

INVx5_ASAP7_75t_L g4417 ( 
.A(n_3792),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_3959),
.B(n_4125),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3949),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_3923),
.A2(n_2822),
.B1(n_2824),
.B2(n_2821),
.Y(n_4420)
);

CKINVDCx20_ASAP7_75t_R g4421 ( 
.A(n_4050),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_SL g4422 ( 
.A(n_3815),
.B(n_3878),
.Y(n_4422)
);

AOI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_3782),
.A2(n_3443),
.B(n_3439),
.Y(n_4423)
);

NOR3xp33_ASAP7_75t_SL g4424 ( 
.A(n_3801),
.B(n_1571),
.C(n_1568),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3926),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4063),
.A2(n_3443),
.B(n_3439),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3930),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_4125),
.B(n_3572),
.Y(n_4428)
);

AOI22xp33_ASAP7_75t_L g4429 ( 
.A1(n_4089),
.A2(n_2826),
.B1(n_2831),
.B2(n_2824),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_3958),
.B(n_789),
.Y(n_4430)
);

AOI22xp5_ASAP7_75t_L g4431 ( 
.A1(n_3981),
.A2(n_1576),
.B1(n_1578),
.B2(n_1571),
.Y(n_4431)
);

CKINVDCx5p33_ASAP7_75t_R g4432 ( 
.A(n_4086),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3933),
.Y(n_4433)
);

BUFx3_ASAP7_75t_L g4434 ( 
.A(n_3883),
.Y(n_4434)
);

NAND2xp33_ASAP7_75t_SL g4435 ( 
.A(n_3826),
.B(n_3140),
.Y(n_4435)
);

NAND2xp33_ASAP7_75t_SL g4436 ( 
.A(n_3837),
.B(n_3198),
.Y(n_4436)
);

BUFx4f_ASAP7_75t_L g4437 ( 
.A(n_3934),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_SL g4438 ( 
.A(n_3878),
.B(n_3198),
.Y(n_4438)
);

OAI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_4000),
.A2(n_3715),
.B1(n_3716),
.B2(n_3709),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_3940),
.Y(n_4440)
);

INVx3_ASAP7_75t_L g4441 ( 
.A(n_3972),
.Y(n_4441)
);

NOR2xp33_ASAP7_75t_L g4442 ( 
.A(n_4084),
.B(n_1576),
.Y(n_4442)
);

BUFx4f_ASAP7_75t_L g4443 ( 
.A(n_3934),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3941),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4092),
.B(n_3974),
.Y(n_4445)
);

CKINVDCx5p33_ASAP7_75t_R g4446 ( 
.A(n_4050),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_SL g4447 ( 
.A(n_4000),
.B(n_3198),
.Y(n_4447)
);

INVx4_ASAP7_75t_L g4448 ( 
.A(n_3965),
.Y(n_4448)
);

BUFx3_ASAP7_75t_L g4449 ( 
.A(n_3875),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_3997),
.B(n_3722),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4010),
.B(n_3723),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4000),
.A2(n_3739),
.B1(n_3770),
.B2(n_3724),
.Y(n_4452)
);

AND2x4_ASAP7_75t_L g4453 ( 
.A(n_4128),
.B(n_3573),
.Y(n_4453)
);

OAI21xp33_ASAP7_75t_SL g4454 ( 
.A1(n_3796),
.A2(n_3548),
.B(n_2608),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_3852),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_4000),
.B(n_3198),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4010),
.B(n_3776),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_3977),
.B(n_3937),
.Y(n_4458)
);

INVxp67_ASAP7_75t_L g4459 ( 
.A(n_3904),
.Y(n_4459)
);

BUFx4f_ASAP7_75t_L g4460 ( 
.A(n_3965),
.Y(n_4460)
);

OR2x2_ASAP7_75t_L g4461 ( 
.A(n_4073),
.B(n_3574),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_3892),
.B(n_3584),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_3853),
.Y(n_4463)
);

INVx3_ASAP7_75t_L g4464 ( 
.A(n_4069),
.Y(n_4464)
);

NAND2xp33_ASAP7_75t_L g4465 ( 
.A(n_3898),
.B(n_3198),
.Y(n_4465)
);

INVx2_ASAP7_75t_SL g4466 ( 
.A(n_4022),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4047),
.B(n_3589),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4047),
.B(n_3590),
.Y(n_4468)
);

BUFx6f_ASAP7_75t_L g4469 ( 
.A(n_3967),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4003),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4117),
.B(n_3695),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4117),
.B(n_3696),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4095),
.B(n_3697),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4005),
.Y(n_4474)
);

NOR2xp33_ASAP7_75t_L g4475 ( 
.A(n_4090),
.B(n_1578),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_3848),
.Y(n_4476)
);

NAND2xp33_ASAP7_75t_L g4477 ( 
.A(n_3901),
.B(n_3204),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4009),
.Y(n_4478)
);

O2A1O1Ixp5_ASAP7_75t_L g4479 ( 
.A1(n_3829),
.A2(n_3548),
.B(n_3454),
.C(n_3456),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4095),
.B(n_3703),
.Y(n_4480)
);

AND2x4_ASAP7_75t_L g4481 ( 
.A(n_3967),
.B(n_3577),
.Y(n_4481)
);

AO22x1_ASAP7_75t_L g4482 ( 
.A1(n_4027),
.A2(n_884),
.B1(n_885),
.B2(n_876),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4105),
.B(n_3578),
.Y(n_4483)
);

OAI22xp5_ASAP7_75t_SL g4484 ( 
.A1(n_4072),
.A2(n_891),
.B1(n_895),
.B2(n_655),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4011),
.Y(n_4485)
);

BUFx3_ASAP7_75t_L g4486 ( 
.A(n_4049),
.Y(n_4486)
);

OAI21x1_ASAP7_75t_L g4487 ( 
.A1(n_4054),
.A2(n_3627),
.B(n_3254),
.Y(n_4487)
);

AND3x1_ASAP7_75t_L g4488 ( 
.A(n_4072),
.B(n_807),
.C(n_800),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_3844),
.Y(n_4489)
);

HB1xp67_ASAP7_75t_L g4490 ( 
.A(n_3918),
.Y(n_4490)
);

INVx2_ASAP7_75t_SL g4491 ( 
.A(n_4091),
.Y(n_4491)
);

INVxp67_ASAP7_75t_SL g4492 ( 
.A(n_3824),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_3950),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_3920),
.B(n_3204),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4018),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_3920),
.B(n_3204),
.Y(n_4496)
);

BUFx6f_ASAP7_75t_L g4497 ( 
.A(n_4049),
.Y(n_4497)
);

AOI22xp5_ASAP7_75t_L g4498 ( 
.A1(n_3937),
.A2(n_1587),
.B1(n_1588),
.B2(n_1582),
.Y(n_4498)
);

AOI22xp5_ASAP7_75t_L g4499 ( 
.A1(n_4027),
.A2(n_4127),
.B1(n_4007),
.B2(n_3954),
.Y(n_4499)
);

NOR2xp33_ASAP7_75t_L g4500 ( 
.A(n_4099),
.B(n_1582),
.Y(n_4500)
);

INVx3_ASAP7_75t_L g4501 ( 
.A(n_4132),
.Y(n_4501)
);

NOR2xp67_ASAP7_75t_L g4502 ( 
.A(n_3970),
.B(n_3260),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_3889),
.B(n_789),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4030),
.Y(n_4504)
);

AND2x2_ASAP7_75t_SL g4505 ( 
.A(n_3785),
.B(n_3094),
.Y(n_4505)
);

AOI22xp5_ASAP7_75t_L g4506 ( 
.A1(n_4041),
.A2(n_1588),
.B1(n_1591),
.B2(n_1587),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_4101),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_SL g4508 ( 
.A(n_3917),
.B(n_3234),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4031),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4105),
.B(n_3579),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_3839),
.B(n_3588),
.Y(n_4511)
);

INVx5_ASAP7_75t_L g4512 ( 
.A(n_3839),
.Y(n_4512)
);

CKINVDCx6p67_ASAP7_75t_R g4513 ( 
.A(n_4103),
.Y(n_4513)
);

AND2x4_ASAP7_75t_L g4514 ( 
.A(n_4074),
.B(n_3702),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_SL g4515 ( 
.A(n_3917),
.B(n_3921),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4403),
.B(n_3705),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_4362),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_4193),
.A2(n_4067),
.B(n_4061),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4419),
.B(n_3719),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4316),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4351),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4193),
.A2(n_3582),
.B(n_3562),
.Y(n_4522)
);

INVx11_ASAP7_75t_L g4523 ( 
.A(n_4164),
.Y(n_4523)
);

CKINVDCx20_ASAP7_75t_R g4524 ( 
.A(n_4186),
.Y(n_4524)
);

OAI21xp5_ASAP7_75t_L g4525 ( 
.A1(n_4243),
.A2(n_4026),
.B(n_3865),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4302),
.B(n_4089),
.Y(n_4526)
);

AOI22xp5_ASAP7_75t_L g4527 ( 
.A1(n_4368),
.A2(n_4041),
.B1(n_3785),
.B2(n_3921),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4490),
.B(n_4258),
.Y(n_4528)
);

NOR2x1_ASAP7_75t_L g4529 ( 
.A(n_4384),
.B(n_4299),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4383),
.B(n_3775),
.Y(n_4530)
);

AOI22xp33_ASAP7_75t_L g4531 ( 
.A1(n_4141),
.A2(n_3976),
.B1(n_3985),
.B2(n_3868),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4458),
.B(n_3976),
.Y(n_4532)
);

OAI321xp33_ASAP7_75t_L g4533 ( 
.A1(n_4408),
.A2(n_3985),
.A3(n_810),
.B1(n_800),
.B2(n_840),
.C(n_813),
.Y(n_4533)
);

INVxp67_ASAP7_75t_L g4534 ( 
.A(n_4434),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_4298),
.A2(n_3582),
.B(n_3562),
.Y(n_4535)
);

AOI22xp5_ASAP7_75t_L g4536 ( 
.A1(n_4347),
.A2(n_4036),
.B1(n_4037),
.B2(n_3840),
.Y(n_4536)
);

NOR2xp33_ASAP7_75t_L g4537 ( 
.A(n_4259),
.B(n_4266),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4322),
.Y(n_4538)
);

OAI22xp5_ASAP7_75t_L g4539 ( 
.A1(n_4235),
.A2(n_4051),
.B1(n_4057),
.B2(n_4055),
.Y(n_4539)
);

AOI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_4488),
.A2(n_4287),
.B1(n_4358),
.B2(n_4343),
.Y(n_4540)
);

BUFx6f_ASAP7_75t_L g4541 ( 
.A(n_4437),
.Y(n_4541)
);

INVx3_ASAP7_75t_L g4542 ( 
.A(n_4170),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4385),
.B(n_4113),
.Y(n_4543)
);

NAND2x1p5_ASAP7_75t_L g4544 ( 
.A(n_4411),
.B(n_3915),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4313),
.B(n_4119),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4202),
.B(n_4121),
.Y(n_4546)
);

AOI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4439),
.A2(n_3753),
.B(n_4068),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4276),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4202),
.B(n_4129),
.Y(n_4549)
);

BUFx8_ASAP7_75t_L g4550 ( 
.A(n_4208),
.Y(n_4550)
);

O2A1O1Ixp5_ASAP7_75t_L g4551 ( 
.A1(n_4515),
.A2(n_3834),
.B(n_3865),
.C(n_4087),
.Y(n_4551)
);

AOI21xp5_ASAP7_75t_L g4552 ( 
.A1(n_4452),
.A2(n_4085),
.B(n_4078),
.Y(n_4552)
);

NOR3xp33_ASAP7_75t_L g4553 ( 
.A(n_4482),
.B(n_3991),
.C(n_813),
.Y(n_4553)
);

A2O1A1Ixp33_ASAP7_75t_L g4554 ( 
.A1(n_4201),
.A2(n_4037),
.B(n_4036),
.C(n_4087),
.Y(n_4554)
);

INVx3_ASAP7_75t_SL g4555 ( 
.A(n_4211),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_SL g4556 ( 
.A(n_4203),
.B(n_4082),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_SL g4557 ( 
.A(n_4205),
.B(n_4024),
.Y(n_4557)
);

O2A1O1Ixp33_ASAP7_75t_SL g4558 ( 
.A1(n_4205),
.A2(n_2635),
.B(n_2633),
.C(n_841),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4440),
.B(n_4035),
.Y(n_4559)
);

AOI21xp5_ASAP7_75t_L g4560 ( 
.A1(n_4452),
.A2(n_4122),
.B(n_4115),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4445),
.B(n_3906),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_4197),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_SL g4563 ( 
.A(n_4502),
.B(n_4301),
.Y(n_4563)
);

OA21x2_ASAP7_75t_L g4564 ( 
.A1(n_4279),
.A2(n_4109),
.B(n_4120),
.Y(n_4564)
);

AOI21xp33_ASAP7_75t_L g4565 ( 
.A1(n_4408),
.A2(n_4109),
.B(n_2422),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4276),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_SL g4567 ( 
.A(n_4499),
.B(n_4024),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4398),
.B(n_4035),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4378),
.B(n_1591),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_4399),
.B(n_3400),
.Y(n_4570)
);

OAI21xp5_ASAP7_75t_L g4571 ( 
.A1(n_4388),
.A2(n_4126),
.B(n_2422),
.Y(n_4571)
);

AND2x4_ASAP7_75t_L g4572 ( 
.A(n_4324),
.B(n_4267),
.Y(n_4572)
);

OAI22xp5_ASAP7_75t_L g4573 ( 
.A1(n_4139),
.A2(n_891),
.B1(n_895),
.B2(n_655),
.Y(n_4573)
);

AOI21x1_ASAP7_75t_L g4574 ( 
.A1(n_4275),
.A2(n_4034),
.B(n_4019),
.Y(n_4574)
);

OAI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_4391),
.A2(n_4404),
.B(n_4294),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_4465),
.A2(n_3939),
.B(n_3938),
.Y(n_4576)
);

AOI21xp5_ASAP7_75t_L g4577 ( 
.A1(n_4477),
.A2(n_3969),
.B(n_3955),
.Y(n_4577)
);

AOI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4182),
.A2(n_4396),
.B(n_4426),
.Y(n_4578)
);

HB1xp67_ASAP7_75t_L g4579 ( 
.A(n_4195),
.Y(n_4579)
);

AOI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4396),
.A2(n_4004),
.B(n_3971),
.Y(n_4580)
);

A2O1A1Ixp33_ASAP7_75t_L g4581 ( 
.A1(n_4442),
.A2(n_4500),
.B(n_4475),
.C(n_4247),
.Y(n_4581)
);

OAI21x1_ASAP7_75t_L g4582 ( 
.A1(n_4487),
.A2(n_3254),
.B(n_3243),
.Y(n_4582)
);

CKINVDCx10_ASAP7_75t_R g4583 ( 
.A(n_4356),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_SL g4584 ( 
.A(n_4437),
.B(n_4065),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4400),
.B(n_3400),
.Y(n_4585)
);

INVx5_ASAP7_75t_L g4586 ( 
.A(n_4411),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4493),
.B(n_3400),
.Y(n_4587)
);

OR2x6_ASAP7_75t_SL g4588 ( 
.A(n_4273),
.B(n_897),
.Y(n_4588)
);

AOI22x1_ASAP7_75t_L g4589 ( 
.A1(n_4296),
.A2(n_898),
.B1(n_899),
.B2(n_897),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4459),
.B(n_3400),
.Y(n_4590)
);

AOI21xp5_ASAP7_75t_L g4591 ( 
.A1(n_4426),
.A2(n_4325),
.B(n_4435),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4314),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_L g4593 ( 
.A1(n_4141),
.A2(n_2826),
.B1(n_2840),
.B2(n_2831),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4425),
.B(n_3625),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4143),
.Y(n_4595)
);

AOI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4325),
.A2(n_4015),
.B(n_4044),
.Y(n_4596)
);

BUFx6f_ASAP7_75t_L g4597 ( 
.A(n_4443),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4314),
.Y(n_4598)
);

OAI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4506),
.A2(n_4371),
.B1(n_4431),
.B2(n_4330),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_SL g4600 ( 
.A(n_4443),
.B(n_4460),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_SL g4601 ( 
.A(n_4460),
.B(n_4028),
.Y(n_4601)
);

AOI21xp33_ASAP7_75t_L g4602 ( 
.A1(n_4199),
.A2(n_2791),
.B(n_2700),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4427),
.B(n_3625),
.Y(n_4603)
);

BUFx6f_ASAP7_75t_L g4604 ( 
.A(n_4150),
.Y(n_4604)
);

AOI22xp5_ASAP7_75t_L g4605 ( 
.A1(n_4363),
.A2(n_3625),
.B1(n_3387),
.B2(n_3302),
.Y(n_4605)
);

AOI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_4436),
.A2(n_4060),
.B(n_4059),
.Y(n_4606)
);

INVx3_ASAP7_75t_SL g4607 ( 
.A(n_4317),
.Y(n_4607)
);

O2A1O1Ixp33_ASAP7_75t_L g4608 ( 
.A1(n_4209),
.A2(n_809),
.B(n_844),
.C(n_840),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4433),
.B(n_3625),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4444),
.B(n_4153),
.Y(n_4610)
);

AOI22x1_ASAP7_75t_L g4611 ( 
.A1(n_4296),
.A2(n_4382),
.B1(n_4365),
.B2(n_4384),
.Y(n_4611)
);

NAND3xp33_ASAP7_75t_L g4612 ( 
.A(n_4498),
.B(n_912),
.C(n_848),
.Y(n_4612)
);

AOI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_4406),
.A2(n_3268),
.B(n_3260),
.Y(n_4613)
);

AND2x4_ASAP7_75t_SL g4614 ( 
.A(n_4142),
.B(n_3234),
.Y(n_4614)
);

INVx3_ASAP7_75t_L g4615 ( 
.A(n_4170),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4152),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4280),
.B(n_841),
.Y(n_4617)
);

INVxp67_ASAP7_75t_L g4618 ( 
.A(n_4155),
.Y(n_4618)
);

AOI21xp5_ASAP7_75t_L g4619 ( 
.A1(n_4423),
.A2(n_3268),
.B(n_3260),
.Y(n_4619)
);

O2A1O1Ixp5_ASAP7_75t_L g4620 ( 
.A1(n_4249),
.A2(n_2840),
.B(n_2848),
.C(n_2841),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4177),
.Y(n_4621)
);

NOR2xp33_ASAP7_75t_L g4622 ( 
.A(n_4179),
.B(n_1596),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4153),
.B(n_3242),
.Y(n_4623)
);

AOI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4397),
.A2(n_3268),
.B(n_3260),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4184),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4180),
.B(n_3242),
.Y(n_4626)
);

AOI21xp33_ASAP7_75t_L g4627 ( 
.A1(n_4180),
.A2(n_4190),
.B(n_4470),
.Y(n_4627)
);

AO21x1_ASAP7_75t_L g4628 ( 
.A1(n_4190),
.A2(n_848),
.B(n_844),
.Y(n_4628)
);

INVxp67_ASAP7_75t_L g4629 ( 
.A(n_4163),
.Y(n_4629)
);

OAI22xp5_ASAP7_75t_L g4630 ( 
.A1(n_4397),
.A2(n_899),
.B1(n_900),
.B2(n_898),
.Y(n_4630)
);

AOI22xp5_ASAP7_75t_L g4631 ( 
.A1(n_4209),
.A2(n_3302),
.B1(n_3387),
.B2(n_938),
.Y(n_4631)
);

OR2x2_ASAP7_75t_L g4632 ( 
.A(n_4461),
.B(n_2700),
.Y(n_4632)
);

INVx3_ASAP7_75t_L g4633 ( 
.A(n_4196),
.Y(n_4633)
);

AOI21x1_ASAP7_75t_L g4634 ( 
.A1(n_4401),
.A2(n_2874),
.B(n_2818),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4393),
.B(n_3141),
.Y(n_4635)
);

NOR2xp67_ASAP7_75t_L g4636 ( 
.A(n_4299),
.B(n_3268),
.Y(n_4636)
);

OAI21xp5_ASAP7_75t_L g4637 ( 
.A1(n_4454),
.A2(n_2853),
.B(n_2818),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_4149),
.B(n_1596),
.Y(n_4638)
);

BUFx8_ASAP7_75t_L g4639 ( 
.A(n_4260),
.Y(n_4639)
);

AOI22xp33_ASAP7_75t_L g4640 ( 
.A1(n_4505),
.A2(n_2841),
.B1(n_2849),
.B2(n_2848),
.Y(n_4640)
);

OAI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_4215),
.A2(n_901),
.B1(n_903),
.B2(n_900),
.Y(n_4641)
);

BUFx6f_ASAP7_75t_L g4642 ( 
.A(n_4150),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_4146),
.A2(n_3343),
.B(n_3334),
.Y(n_4643)
);

AOI22x1_ASAP7_75t_L g4644 ( 
.A1(n_4346),
.A2(n_903),
.B1(n_905),
.B2(n_901),
.Y(n_4644)
);

AND2x4_ASAP7_75t_L g4645 ( 
.A(n_4324),
.B(n_3377),
.Y(n_4645)
);

BUFx2_ASAP7_75t_L g4646 ( 
.A(n_4257),
.Y(n_4646)
);

BUFx6f_ASAP7_75t_L g4647 ( 
.A(n_4150),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4151),
.A2(n_4456),
.B(n_4447),
.Y(n_4648)
);

AOI22xp5_ASAP7_75t_L g4649 ( 
.A1(n_4366),
.A2(n_3302),
.B1(n_3387),
.B2(n_940),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_SL g4650 ( 
.A(n_4364),
.B(n_3234),
.Y(n_4650)
);

AOI22xp5_ASAP7_75t_L g4651 ( 
.A1(n_4308),
.A2(n_3302),
.B1(n_3387),
.B2(n_978),
.Y(n_4651)
);

AOI22x1_ASAP7_75t_L g4652 ( 
.A1(n_4346),
.A2(n_908),
.B1(n_910),
.B2(n_905),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4151),
.A2(n_3343),
.B(n_3334),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4244),
.Y(n_4654)
);

AOI22xp5_ASAP7_75t_L g4655 ( 
.A1(n_4421),
.A2(n_1026),
.B1(n_1028),
.B2(n_934),
.Y(n_4655)
);

AOI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4336),
.A2(n_3343),
.B(n_3334),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4455),
.B(n_3144),
.Y(n_4657)
);

AOI21xp5_ASAP7_75t_L g4658 ( 
.A1(n_4154),
.A2(n_3343),
.B(n_3334),
.Y(n_4658)
);

AOI21xp5_ASAP7_75t_L g4659 ( 
.A1(n_4154),
.A2(n_3343),
.B(n_3334),
.Y(n_4659)
);

O2A1O1Ixp5_ASAP7_75t_L g4660 ( 
.A1(n_4494),
.A2(n_4496),
.B(n_4508),
.C(n_4355),
.Y(n_4660)
);

OAI21xp5_ASAP7_75t_L g4661 ( 
.A1(n_4479),
.A2(n_2771),
.B(n_3344),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4187),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4463),
.B(n_4233),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4253),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4233),
.B(n_4476),
.Y(n_4665)
);

AOI21x1_ASAP7_75t_L g4666 ( 
.A1(n_4248),
.A2(n_2874),
.B(n_2771),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4328),
.B(n_3144),
.Y(n_4667)
);

AOI21xp5_ASAP7_75t_L g4668 ( 
.A1(n_4194),
.A2(n_2969),
.B(n_3234),
.Y(n_4668)
);

AO21x1_ASAP7_75t_L g4669 ( 
.A1(n_4422),
.A2(n_869),
.B(n_868),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4255),
.Y(n_4670)
);

AOI21xp5_ASAP7_75t_L g4671 ( 
.A1(n_4372),
.A2(n_3257),
.B(n_3251),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4372),
.A2(n_3257),
.B(n_3251),
.Y(n_4672)
);

OAI22xp5_ASAP7_75t_L g4673 ( 
.A1(n_4245),
.A2(n_4213),
.B1(n_4210),
.B2(n_4212),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4305),
.B(n_868),
.Y(n_4674)
);

INVx2_ASAP7_75t_L g4675 ( 
.A(n_4218),
.Y(n_4675)
);

NAND3xp33_ASAP7_75t_L g4676 ( 
.A(n_4387),
.B(n_889),
.C(n_878),
.Y(n_4676)
);

AOI21xp5_ASAP7_75t_L g4677 ( 
.A1(n_4415),
.A2(n_3257),
.B(n_3251),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4394),
.B(n_3145),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4305),
.B(n_869),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4394),
.B(n_3145),
.Y(n_4680)
);

OAI22xp5_ASAP7_75t_L g4681 ( 
.A1(n_4210),
.A2(n_910),
.B1(n_924),
.B2(n_908),
.Y(n_4681)
);

INVx4_ASAP7_75t_L g4682 ( 
.A(n_4191),
.Y(n_4682)
);

AOI21xp5_ASAP7_75t_L g4683 ( 
.A1(n_4415),
.A2(n_3257),
.B(n_3251),
.Y(n_4683)
);

OAI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4479),
.A2(n_4145),
.B(n_4412),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4257),
.Y(n_4685)
);

INVxp67_ASAP7_75t_L g4686 ( 
.A(n_4252),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4320),
.B(n_875),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_SL g4688 ( 
.A(n_4213),
.B(n_3271),
.Y(n_4688)
);

OAI22x1_ASAP7_75t_L g4689 ( 
.A1(n_4361),
.A2(n_1049),
.B1(n_1074),
.B2(n_1042),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4320),
.B(n_875),
.Y(n_4690)
);

AOI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4417),
.A2(n_3276),
.B(n_3271),
.Y(n_4691)
);

NAND2x1p5_ASAP7_75t_L g4692 ( 
.A(n_4417),
.B(n_3377),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4417),
.A2(n_3276),
.B(n_3271),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4269),
.Y(n_4694)
);

AOI21xp33_ASAP7_75t_L g4695 ( 
.A1(n_4474),
.A2(n_2791),
.B(n_2700),
.Y(n_4695)
);

BUFx3_ASAP7_75t_L g4696 ( 
.A(n_4231),
.Y(n_4696)
);

AOI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4198),
.A2(n_3296),
.B(n_3276),
.Y(n_4697)
);

NAND3xp33_ASAP7_75t_L g4698 ( 
.A(n_4424),
.B(n_920),
.C(n_881),
.Y(n_4698)
);

INVx2_ASAP7_75t_L g4699 ( 
.A(n_4225),
.Y(n_4699)
);

O2A1O1Ixp33_ASAP7_75t_L g4700 ( 
.A1(n_4334),
.A2(n_878),
.B(n_887),
.C(n_886),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4478),
.B(n_3146),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4485),
.B(n_3146),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4504),
.B(n_3147),
.Y(n_4703)
);

CKINVDCx20_ASAP7_75t_R g4704 ( 
.A(n_4446),
.Y(n_4704)
);

AOI22xp5_ASAP7_75t_L g4705 ( 
.A1(n_4386),
.A2(n_1099),
.B1(n_1122),
.B2(n_1077),
.Y(n_4705)
);

NAND2x1p5_ASAP7_75t_L g4706 ( 
.A(n_4267),
.B(n_3377),
.Y(n_4706)
);

O2A1O1Ixp33_ASAP7_75t_L g4707 ( 
.A1(n_4430),
.A2(n_881),
.B(n_887),
.C(n_886),
.Y(n_4707)
);

NOR2xp33_ASAP7_75t_L g4708 ( 
.A(n_4166),
.B(n_4311),
.Y(n_4708)
);

INVx1_ASAP7_75t_SL g4709 ( 
.A(n_4188),
.Y(n_4709)
);

AOI21xp5_ASAP7_75t_L g4710 ( 
.A1(n_4226),
.A2(n_3297),
.B(n_3296),
.Y(n_4710)
);

OAI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4503),
.A2(n_4289),
.B(n_4428),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4509),
.B(n_4489),
.Y(n_4712)
);

AOI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4254),
.A2(n_3297),
.B(n_3296),
.Y(n_4713)
);

NAND2xp5_ASAP7_75t_SL g4714 ( 
.A(n_4514),
.B(n_3297),
.Y(n_4714)
);

NOR2xp33_ASAP7_75t_L g4715 ( 
.A(n_4181),
.B(n_1600),
.Y(n_4715)
);

INVx5_ASAP7_75t_L g4716 ( 
.A(n_4217),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_4514),
.B(n_3307),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4332),
.B(n_3147),
.Y(n_4718)
);

AO21x1_ASAP7_75t_L g4719 ( 
.A1(n_4221),
.A2(n_912),
.B(n_889),
.Y(n_4719)
);

O2A1O1Ixp33_ASAP7_75t_SL g4720 ( 
.A1(n_4157),
.A2(n_919),
.B(n_920),
.C(n_914),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4369),
.B(n_914),
.Y(n_4721)
);

AOI22x1_ASAP7_75t_L g4722 ( 
.A1(n_4350),
.A2(n_1190),
.B1(n_924),
.B2(n_1600),
.Y(n_4722)
);

NOR2xp33_ASAP7_75t_L g4723 ( 
.A(n_4250),
.B(n_1603),
.Y(n_4723)
);

INVx11_ASAP7_75t_L g4724 ( 
.A(n_4352),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_SL g4725 ( 
.A(n_4418),
.B(n_4507),
.Y(n_4725)
);

BUFx6f_ASAP7_75t_L g4726 ( 
.A(n_4191),
.Y(n_4726)
);

AOI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_4254),
.A2(n_3314),
.B(n_3307),
.Y(n_4727)
);

AND2x6_ASAP7_75t_L g4728 ( 
.A(n_4464),
.B(n_2921),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4450),
.B(n_3148),
.Y(n_4729)
);

AO22x1_ASAP7_75t_L g4730 ( 
.A1(n_4217),
.A2(n_919),
.B1(n_936),
.B2(n_918),
.Y(n_4730)
);

AOI21x1_ASAP7_75t_L g4731 ( 
.A1(n_4261),
.A2(n_2874),
.B(n_2791),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_4513),
.B(n_1603),
.Y(n_4732)
);

NOR2xp33_ASAP7_75t_L g4733 ( 
.A(n_4140),
.B(n_1604),
.Y(n_4733)
);

A2O1A1Ixp33_ASAP7_75t_L g4734 ( 
.A1(n_4418),
.A2(n_1139),
.B(n_1188),
.C(n_1126),
.Y(n_4734)
);

NOR2xp67_ASAP7_75t_L g4735 ( 
.A(n_4158),
.B(n_2938),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4228),
.Y(n_4736)
);

NAND2x1_ASAP7_75t_L g4737 ( 
.A(n_4217),
.B(n_3119),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4450),
.B(n_3148),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4451),
.B(n_4457),
.Y(n_4739)
);

NOR2xp33_ASAP7_75t_R g4740 ( 
.A(n_4432),
.B(n_3220),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_L g4741 ( 
.A1(n_4512),
.A2(n_2849),
.B1(n_2855),
.B2(n_2852),
.Y(n_4741)
);

AOI22xp5_ASAP7_75t_L g4742 ( 
.A1(n_4484),
.A2(n_1612),
.B1(n_1621),
.B2(n_1604),
.Y(n_4742)
);

INVx4_ASAP7_75t_L g4743 ( 
.A(n_4191),
.Y(n_4743)
);

AOI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_4375),
.A2(n_4377),
.B(n_4379),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4241),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4274),
.Y(n_4746)
);

NOR2xp33_ASAP7_75t_L g4747 ( 
.A(n_4192),
.B(n_1612),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4457),
.B(n_3152),
.Y(n_4748)
);

AOI21xp5_ASAP7_75t_L g4749 ( 
.A1(n_4377),
.A2(n_3314),
.B(n_3307),
.Y(n_4749)
);

OAI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_4512),
.A2(n_1190),
.B1(n_936),
.B2(n_939),
.Y(n_4750)
);

INVx3_ASAP7_75t_L g4751 ( 
.A(n_4196),
.Y(n_4751)
);

OAI22xp5_ASAP7_75t_L g4752 ( 
.A1(n_4512),
.A2(n_939),
.B1(n_941),
.B2(n_918),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4277),
.Y(n_4753)
);

AOI21xp5_ASAP7_75t_L g4754 ( 
.A1(n_4379),
.A2(n_3314),
.B(n_3307),
.Y(n_4754)
);

AOI21x1_ASAP7_75t_L g4755 ( 
.A1(n_4438),
.A2(n_4407),
.B(n_4342),
.Y(n_4755)
);

OAI21xp5_ASAP7_75t_L g4756 ( 
.A1(n_4428),
.A2(n_3344),
.B(n_2855),
.Y(n_4756)
);

AOI22xp5_ASAP7_75t_L g4757 ( 
.A1(n_4402),
.A2(n_1622),
.B1(n_1628),
.B2(n_1621),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4495),
.B(n_3156),
.Y(n_4758)
);

BUFx2_ASAP7_75t_L g4759 ( 
.A(n_4229),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4392),
.B(n_3156),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4251),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_SL g4762 ( 
.A(n_4491),
.B(n_3314),
.Y(n_4762)
);

OAI22xp5_ASAP7_75t_L g4763 ( 
.A1(n_4512),
.A2(n_4283),
.B1(n_4221),
.B2(n_4223),
.Y(n_4763)
);

AOI21xp5_ASAP7_75t_L g4764 ( 
.A1(n_4392),
.A2(n_3339),
.B(n_3320),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4449),
.B(n_3157),
.Y(n_4765)
);

A2O1A1Ixp33_ASAP7_75t_L g4766 ( 
.A1(n_4492),
.A2(n_948),
.B(n_950),
.C(n_941),
.Y(n_4766)
);

INVxp67_ASAP7_75t_L g4767 ( 
.A(n_4291),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4278),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4282),
.Y(n_4769)
);

OAI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4236),
.A2(n_2856),
.B(n_2852),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_SL g4771 ( 
.A(n_4469),
.B(n_3320),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_SL g4772 ( 
.A(n_4267),
.B(n_2938),
.Y(n_4772)
);

AOI21xp33_ASAP7_75t_L g4773 ( 
.A1(n_4236),
.A2(n_2791),
.B(n_2700),
.Y(n_4773)
);

BUFx3_ASAP7_75t_L g4774 ( 
.A(n_4169),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4223),
.B(n_3157),
.Y(n_4775)
);

NAND2x1p5_ASAP7_75t_L g4776 ( 
.A(n_4267),
.B(n_3220),
.Y(n_4776)
);

AOI21xp5_ASAP7_75t_L g4777 ( 
.A1(n_4281),
.A2(n_3339),
.B(n_3320),
.Y(n_4777)
);

BUFx12f_ASAP7_75t_L g4778 ( 
.A(n_4307),
.Y(n_4778)
);

A2O1A1Ixp33_ASAP7_75t_L g4779 ( 
.A1(n_4467),
.A2(n_950),
.B(n_951),
.C(n_948),
.Y(n_4779)
);

O2A1O1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4162),
.A2(n_955),
.B(n_960),
.C(n_956),
.Y(n_4780)
);

NOR2xp33_ASAP7_75t_L g4781 ( 
.A(n_4171),
.B(n_1622),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4369),
.B(n_3160),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_SL g4783 ( 
.A(n_4469),
.B(n_3320),
.Y(n_4783)
);

OAI21xp33_ASAP7_75t_L g4784 ( 
.A1(n_4471),
.A2(n_955),
.B(n_951),
.Y(n_4784)
);

AND2x6_ASAP7_75t_L g4785 ( 
.A(n_4464),
.B(n_2921),
.Y(n_4785)
);

NOR2xp33_ASAP7_75t_L g4786 ( 
.A(n_4138),
.B(n_1628),
.Y(n_4786)
);

INVx3_ASAP7_75t_L g4787 ( 
.A(n_4227),
.Y(n_4787)
);

AOI22x1_ASAP7_75t_L g4788 ( 
.A1(n_4200),
.A2(n_1635),
.B1(n_1639),
.B2(n_1633),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4318),
.A2(n_3339),
.B(n_3320),
.Y(n_4789)
);

NAND3xp33_ASAP7_75t_L g4790 ( 
.A(n_4462),
.B(n_969),
.C(n_956),
.Y(n_4790)
);

NOR2x1_ASAP7_75t_L g4791 ( 
.A(n_4345),
.B(n_2938),
.Y(n_4791)
);

AOI21xp5_ASAP7_75t_L g4792 ( 
.A1(n_4467),
.A2(n_3346),
.B(n_3339),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4237),
.B(n_3160),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4227),
.B(n_960),
.Y(n_4794)
);

AOI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4468),
.A2(n_3346),
.B(n_3339),
.Y(n_4795)
);

NOR2xp33_ASAP7_75t_L g4796 ( 
.A(n_4138),
.B(n_1633),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4138),
.B(n_1635),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4238),
.B(n_1639),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4468),
.A2(n_3348),
.B(n_3346),
.Y(n_4799)
);

HB1xp67_ASAP7_75t_L g4800 ( 
.A(n_4286),
.Y(n_4800)
);

O2A1O1Ixp5_ASAP7_75t_L g4801 ( 
.A1(n_4348),
.A2(n_2856),
.B(n_2859),
.C(n_2858),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4237),
.B(n_3172),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4293),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4239),
.B(n_3172),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4239),
.B(n_3179),
.Y(n_4805)
);

BUFx4f_ASAP7_75t_L g4806 ( 
.A(n_4307),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_4224),
.B(n_1640),
.Y(n_4807)
);

AOI22xp33_ASAP7_75t_L g4808 ( 
.A1(n_4183),
.A2(n_2858),
.B1(n_2862),
.B2(n_2859),
.Y(n_4808)
);

AOI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4246),
.A2(n_3348),
.B(n_3346),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4246),
.A2(n_3348),
.B(n_3346),
.Y(n_4810)
);

NOR2xp67_ASAP7_75t_L g4811 ( 
.A(n_4324),
.B(n_2938),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4473),
.B(n_3179),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4473),
.B(n_3180),
.Y(n_4813)
);

BUFx2_ASAP7_75t_L g4814 ( 
.A(n_4353),
.Y(n_4814)
);

NAND2x1p5_ASAP7_75t_L g4815 ( 
.A(n_4324),
.B(n_3253),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4480),
.B(n_3180),
.Y(n_4816)
);

AO22x1_ASAP7_75t_L g4817 ( 
.A1(n_4217),
.A2(n_973),
.B1(n_991),
.B2(n_969),
.Y(n_4817)
);

OR2x6_ASAP7_75t_SL g4818 ( 
.A(n_4480),
.B(n_880),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4376),
.B(n_1640),
.Y(n_4819)
);

OR2x6_ASAP7_75t_SL g4820 ( 
.A(n_4483),
.B(n_4510),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4483),
.B(n_3182),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4297),
.Y(n_4822)
);

NOR2xp67_ASAP7_75t_L g4823 ( 
.A(n_4501),
.B(n_3044),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4497),
.B(n_3352),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4510),
.B(n_3182),
.Y(n_4825)
);

BUFx8_ASAP7_75t_L g4826 ( 
.A(n_4356),
.Y(n_4826)
);

NOR2xp67_ASAP7_75t_SL g4827 ( 
.A(n_4200),
.B(n_3253),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4304),
.B(n_3185),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4511),
.A2(n_3368),
.B(n_3352),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4309),
.Y(n_4830)
);

OAI21xp33_ASAP7_75t_L g4831 ( 
.A1(n_4471),
.A2(n_991),
.B(n_973),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4511),
.A2(n_3368),
.B(n_3352),
.Y(n_4832)
);

NAND3xp33_ASAP7_75t_L g4833 ( 
.A(n_4462),
.B(n_1033),
.C(n_1018),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_L g4834 ( 
.A1(n_4290),
.A2(n_999),
.B(n_1001),
.C(n_993),
.Y(n_4834)
);

A2O1A1Ixp33_ASAP7_75t_L g4835 ( 
.A1(n_4315),
.A2(n_999),
.B(n_1001),
.C(n_993),
.Y(n_4835)
);

AOI21xp5_ASAP7_75t_L g4836 ( 
.A1(n_4300),
.A2(n_3368),
.B(n_3154),
.Y(n_4836)
);

OAI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_4429),
.A2(n_2864),
.B(n_2862),
.Y(n_4837)
);

NOR2xp33_ASAP7_75t_L g4838 ( 
.A(n_4486),
.B(n_1642),
.Y(n_4838)
);

HB1xp67_ASAP7_75t_L g4839 ( 
.A(n_4344),
.Y(n_4839)
);

AOI21xp5_ASAP7_75t_L g4840 ( 
.A1(n_4300),
.A2(n_3154),
.B(n_3044),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4357),
.B(n_4360),
.Y(n_4841)
);

A2O1A1Ixp33_ASAP7_75t_L g4842 ( 
.A1(n_4453),
.A2(n_1013),
.B(n_1014),
.C(n_1007),
.Y(n_4842)
);

AOI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4472),
.A2(n_3154),
.B(n_3044),
.Y(n_4843)
);

AOI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4472),
.A2(n_3267),
.B(n_3224),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4370),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4147),
.Y(n_4846)
);

AOI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4234),
.A2(n_3267),
.B(n_3224),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4148),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4234),
.B(n_1007),
.Y(n_4849)
);

AOI22xp5_ASAP7_75t_L g4850 ( 
.A1(n_4395),
.A2(n_4453),
.B1(n_4292),
.B2(n_4319),
.Y(n_4850)
);

NOR3xp33_ASAP7_75t_L g4851 ( 
.A(n_4337),
.B(n_1014),
.C(n_1013),
.Y(n_4851)
);

OAI21x1_ASAP7_75t_L g4852 ( 
.A1(n_4501),
.A2(n_3262),
.B(n_3259),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4262),
.B(n_3190),
.Y(n_4853)
);

NOR2xp33_ASAP7_75t_L g4854 ( 
.A(n_4448),
.B(n_1643),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4380),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4262),
.B(n_3190),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4268),
.B(n_3194),
.Y(n_4857)
);

OAI22xp5_ASAP7_75t_L g4858 ( 
.A1(n_4339),
.A2(n_4420),
.B1(n_4272),
.B2(n_4285),
.Y(n_4858)
);

OAI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4268),
.A2(n_2866),
.B(n_2864),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4156),
.Y(n_4860)
);

AOI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_4292),
.A2(n_1648),
.B1(n_1651),
.B2(n_1643),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4448),
.B(n_1648),
.Y(n_4862)
);

NOR2xp33_ASAP7_75t_R g4863 ( 
.A(n_4222),
.B(n_3253),
.Y(n_4863)
);

AOI21x1_ASAP7_75t_L g4864 ( 
.A1(n_4389),
.A2(n_3264),
.B(n_3262),
.Y(n_4864)
);

AOI22xp5_ASAP7_75t_L g4865 ( 
.A1(n_4292),
.A2(n_1652),
.B1(n_1659),
.B2(n_1651),
.Y(n_4865)
);

AND2x4_ASAP7_75t_L g4866 ( 
.A(n_4319),
.B(n_3277),
.Y(n_4866)
);

BUFx2_ASAP7_75t_SL g4867 ( 
.A(n_4405),
.Y(n_4867)
);

OAI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_4272),
.A2(n_2914),
.B(n_2866),
.Y(n_4868)
);

AOI21xp5_ASAP7_75t_L g4869 ( 
.A1(n_4285),
.A2(n_3267),
.B(n_3224),
.Y(n_4869)
);

AOI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_4319),
.A2(n_1659),
.B1(n_1652),
.B2(n_2967),
.Y(n_4870)
);

AOI21xp5_ASAP7_75t_L g4871 ( 
.A1(n_4303),
.A2(n_3267),
.B(n_3224),
.Y(n_4871)
);

AOI21xp5_ASAP7_75t_L g4872 ( 
.A1(n_4303),
.A2(n_2924),
.B(n_2921),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_L g4873 ( 
.A(n_4481),
.B(n_882),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4306),
.B(n_3195),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4310),
.B(n_3195),
.Y(n_4875)
);

NOR2xp33_ASAP7_75t_L g4876 ( 
.A(n_4481),
.B(n_883),
.Y(n_4876)
);

CKINVDCx10_ASAP7_75t_R g4877 ( 
.A(n_4172),
.Y(n_4877)
);

A2O1A1Ixp33_ASAP7_75t_L g4878 ( 
.A1(n_4310),
.A2(n_1023),
.B(n_1025),
.C(n_1018),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_SL g4879 ( 
.A(n_4497),
.B(n_2967),
.Y(n_4879)
);

AOI22x1_ASAP7_75t_L g4880 ( 
.A1(n_4222),
.A2(n_913),
.B1(n_915),
.B2(n_890),
.Y(n_4880)
);

NOR2xp33_ASAP7_75t_L g4881 ( 
.A(n_4307),
.B(n_917),
.Y(n_4881)
);

BUFx2_ASAP7_75t_L g4882 ( 
.A(n_4414),
.Y(n_4882)
);

NOR2xp33_ASAP7_75t_L g4883 ( 
.A(n_4341),
.B(n_921),
.Y(n_4883)
);

CKINVDCx10_ASAP7_75t_R g4884 ( 
.A(n_4207),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4326),
.B(n_3196),
.Y(n_4885)
);

INVx3_ASAP7_75t_L g4886 ( 
.A(n_4341),
.Y(n_4886)
);

O2A1O1Ixp33_ASAP7_75t_L g4887 ( 
.A1(n_4326),
.A2(n_1025),
.B(n_1033),
.C(n_1023),
.Y(n_4887)
);

BUFx6f_ASAP7_75t_L g4888 ( 
.A(n_4341),
.Y(n_4888)
);

NAND2x1p5_ASAP7_75t_L g4889 ( 
.A(n_4441),
.B(n_3277),
.Y(n_4889)
);

NOR2x1p5_ASAP7_75t_L g4890 ( 
.A(n_4413),
.B(n_1034),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_L g4891 ( 
.A1(n_4144),
.A2(n_2914),
.B1(n_2273),
.B2(n_2235),
.Y(n_4891)
);

O2A1O1Ixp33_ASAP7_75t_L g4892 ( 
.A1(n_4329),
.A2(n_1039),
.B(n_1052),
.C(n_1041),
.Y(n_4892)
);

O2A1O1Ixp33_ASAP7_75t_L g4893 ( 
.A1(n_4329),
.A2(n_1039),
.B(n_1052),
.C(n_1041),
.Y(n_4893)
);

OR2x6_ASAP7_75t_L g4894 ( 
.A(n_4264),
.B(n_3000),
.Y(n_4894)
);

AOI21x1_ASAP7_75t_L g4895 ( 
.A1(n_4331),
.A2(n_3266),
.B(n_3264),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4331),
.B(n_3196),
.Y(n_4896)
);

A2O1A1Ixp33_ASAP7_75t_L g4897 ( 
.A1(n_4333),
.A2(n_1055),
.B(n_1058),
.C(n_1034),
.Y(n_4897)
);

INVx2_ASAP7_75t_SL g4898 ( 
.A(n_4354),
.Y(n_4898)
);

A2O1A1Ixp33_ASAP7_75t_L g4899 ( 
.A1(n_4333),
.A2(n_1058),
.B(n_1062),
.C(n_1055),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_L g4900 ( 
.A(n_4338),
.B(n_3202),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4338),
.B(n_3202),
.Y(n_4901)
);

A2O1A1Ixp33_ASAP7_75t_L g4902 ( 
.A1(n_4575),
.A2(n_1069),
.B(n_1070),
.C(n_1062),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_SL g4903 ( 
.A(n_4575),
.B(n_4354),
.Y(n_4903)
);

OAI21x1_ASAP7_75t_L g4904 ( 
.A1(n_4620),
.A2(n_4441),
.B(n_4265),
.Y(n_4904)
);

OAI22x1_ASAP7_75t_L g4905 ( 
.A1(n_4540),
.A2(n_4527),
.B1(n_4890),
.B2(n_4534),
.Y(n_4905)
);

OAI21xp5_ASAP7_75t_L g4906 ( 
.A1(n_4525),
.A2(n_4367),
.B(n_4359),
.Y(n_4906)
);

INVx3_ASAP7_75t_L g4907 ( 
.A(n_4716),
.Y(n_4907)
);

OAI22xp5_ASAP7_75t_L g4908 ( 
.A1(n_4531),
.A2(n_4567),
.B1(n_4537),
.B2(n_4525),
.Y(n_4908)
);

AOI21x1_ASAP7_75t_L g4909 ( 
.A1(n_4730),
.A2(n_4367),
.B(n_4359),
.Y(n_4909)
);

BUFx2_ASAP7_75t_L g4910 ( 
.A(n_4759),
.Y(n_4910)
);

AOI21xp5_ASAP7_75t_L g4911 ( 
.A1(n_4591),
.A2(n_4264),
.B(n_4219),
.Y(n_4911)
);

OAI21x1_ASAP7_75t_L g4912 ( 
.A1(n_4619),
.A2(n_4265),
.B(n_4263),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4800),
.Y(n_4913)
);

AND2x2_ASAP7_75t_L g4914 ( 
.A(n_4814),
.B(n_4142),
.Y(n_4914)
);

NAND3xp33_ASAP7_75t_L g4915 ( 
.A(n_4581),
.B(n_1070),
.C(n_1069),
.Y(n_4915)
);

A2O1A1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_4553),
.A2(n_1081),
.B(n_1092),
.C(n_1080),
.Y(n_4916)
);

OAI22x1_ASAP7_75t_L g4917 ( 
.A1(n_4646),
.A2(n_4160),
.B1(n_4161),
.B2(n_4159),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4820),
.B(n_4167),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4542),
.B(n_4240),
.Y(n_4919)
);

AO31x2_ASAP7_75t_L g4920 ( 
.A1(n_4763),
.A2(n_4173),
.A3(n_4174),
.B(n_4168),
.Y(n_4920)
);

AOI21x1_ASAP7_75t_L g4921 ( 
.A1(n_4817),
.A2(n_4628),
.B(n_4556),
.Y(n_4921)
);

A2O1A1Ixp33_ASAP7_75t_L g4922 ( 
.A1(n_4569),
.A2(n_1081),
.B(n_1092),
.C(n_1080),
.Y(n_4922)
);

NAND3x1_ASAP7_75t_L g4923 ( 
.A(n_4529),
.B(n_4321),
.C(n_4288),
.Y(n_4923)
);

AOI221xp5_ASAP7_75t_L g4924 ( 
.A1(n_4681),
.A2(n_4599),
.B1(n_4700),
.B2(n_4734),
.C(n_4608),
.Y(n_4924)
);

AOI21xp33_ASAP7_75t_L g4925 ( 
.A1(n_4750),
.A2(n_4752),
.B(n_4763),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_SL g4926 ( 
.A(n_4716),
.B(n_4354),
.Y(n_4926)
);

OAI21x1_ASAP7_75t_SL g4927 ( 
.A1(n_4684),
.A2(n_4466),
.B(n_4409),
.Y(n_4927)
);

OAI222xp33_ASAP7_75t_L g4928 ( 
.A1(n_4750),
.A2(n_4185),
.B1(n_4176),
.B2(n_4189),
.C1(n_4178),
.C2(n_4175),
.Y(n_4928)
);

NAND2x1p5_ASAP7_75t_L g4929 ( 
.A(n_4716),
.B(n_4271),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4716),
.B(n_4373),
.Y(n_4930)
);

AND2x2_ASAP7_75t_L g4931 ( 
.A(n_4542),
.B(n_4335),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4803),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4839),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4615),
.B(n_4374),
.Y(n_4934)
);

AND2x2_ASAP7_75t_L g4935 ( 
.A(n_4615),
.B(n_4381),
.Y(n_4935)
);

O2A1O1Ixp5_ASAP7_75t_L g4936 ( 
.A1(n_4557),
.A2(n_4390),
.B(n_1110),
.C(n_1118),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_4578),
.A2(n_4264),
.B(n_4219),
.Y(n_4937)
);

OAI21x1_ASAP7_75t_L g4938 ( 
.A1(n_4637),
.A2(n_4165),
.B(n_3272),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4739),
.B(n_4204),
.Y(n_4939)
);

NOR2x1_ASAP7_75t_SL g4940 ( 
.A(n_4894),
.B(n_4207),
.Y(n_4940)
);

AOI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4624),
.A2(n_4219),
.B(n_4207),
.Y(n_4941)
);

AOI21xp33_ASAP7_75t_L g4942 ( 
.A1(n_4752),
.A2(n_4214),
.B(n_4206),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4744),
.B(n_4216),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4520),
.Y(n_4944)
);

AO31x2_ASAP7_75t_L g4945 ( 
.A1(n_4673),
.A2(n_4230),
.A3(n_4232),
.B(n_4220),
.Y(n_4945)
);

INVx3_ASAP7_75t_L g4946 ( 
.A(n_4633),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4538),
.Y(n_4947)
);

OAI21x1_ASAP7_75t_L g4948 ( 
.A1(n_4792),
.A2(n_3272),
.B(n_3266),
.Y(n_4948)
);

OAI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4571),
.A2(n_1119),
.B(n_1108),
.Y(n_4949)
);

OAI22xp5_ASAP7_75t_L g4950 ( 
.A1(n_4573),
.A2(n_4410),
.B1(n_1121),
.B2(n_1123),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4521),
.Y(n_4951)
);

AOI221x1_ASAP7_75t_L g4952 ( 
.A1(n_4689),
.A2(n_4242),
.B1(n_1123),
.B2(n_1124),
.C(n_1121),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4610),
.B(n_4373),
.Y(n_4953)
);

AND2x4_ASAP7_75t_L g4954 ( 
.A(n_4633),
.B(n_4416),
.Y(n_4954)
);

AOI221x1_ASAP7_75t_L g4955 ( 
.A1(n_4627),
.A2(n_4851),
.B1(n_4681),
.B2(n_4684),
.C(n_4543),
.Y(n_4955)
);

INVx3_ASAP7_75t_L g4956 ( 
.A(n_4751),
.Y(n_4956)
);

AO31x2_ASAP7_75t_L g4957 ( 
.A1(n_4673),
.A2(n_4270),
.A3(n_4284),
.B(n_4256),
.Y(n_4957)
);

NOR2x1_ASAP7_75t_L g4958 ( 
.A(n_4545),
.B(n_4416),
.Y(n_4958)
);

OAI21x1_ASAP7_75t_L g4959 ( 
.A1(n_4795),
.A2(n_3279),
.B(n_3273),
.Y(n_4959)
);

NOR2xp33_ASAP7_75t_L g4960 ( 
.A(n_4704),
.B(n_34),
.Y(n_4960)
);

NAND2x1_ASAP7_75t_SL g4961 ( 
.A(n_4685),
.B(n_1119),
.Y(n_4961)
);

INVx1_ASAP7_75t_SL g4962 ( 
.A(n_4709),
.Y(n_4962)
);

AO21x1_ASAP7_75t_L g4963 ( 
.A1(n_4573),
.A2(n_1134),
.B(n_1124),
.Y(n_4963)
);

OAI21x1_ASAP7_75t_L g4964 ( 
.A1(n_4799),
.A2(n_3279),
.B(n_3273),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4818),
.A2(n_1136),
.B1(n_1145),
.B2(n_1134),
.Y(n_4965)
);

OAI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4571),
.A2(n_1145),
.B(n_1136),
.Y(n_4966)
);

AOI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_4643),
.A2(n_4416),
.B(n_3376),
.Y(n_4967)
);

AOI21xp5_ASAP7_75t_L g4968 ( 
.A1(n_4653),
.A2(n_3376),
.B(n_3373),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_SL g4969 ( 
.A(n_4863),
.B(n_4497),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4551),
.A2(n_1158),
.B(n_1155),
.Y(n_4970)
);

CKINVDCx14_ASAP7_75t_R g4971 ( 
.A(n_4524),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_4550),
.Y(n_4972)
);

BUFx6f_ASAP7_75t_L g4973 ( 
.A(n_4541),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4841),
.Y(n_4974)
);

AOI21xp5_ASAP7_75t_L g4975 ( 
.A1(n_4671),
.A2(n_3379),
.B(n_3373),
.Y(n_4975)
);

INVx1_ASAP7_75t_SL g4976 ( 
.A(n_4709),
.Y(n_4976)
);

CKINVDCx16_ASAP7_75t_R g4977 ( 
.A(n_4740),
.Y(n_4977)
);

OAI21x1_ASAP7_75t_L g4978 ( 
.A1(n_4829),
.A2(n_3347),
.B(n_3289),
.Y(n_4978)
);

OAI21x1_ASAP7_75t_L g4979 ( 
.A1(n_4832),
.A2(n_4666),
.B(n_4634),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4672),
.A2(n_3386),
.B(n_3379),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4654),
.Y(n_4981)
);

HB1xp67_ASAP7_75t_L g4982 ( 
.A(n_4579),
.Y(n_4982)
);

OAI21x1_ASAP7_75t_L g4983 ( 
.A1(n_4864),
.A2(n_3347),
.B(n_3289),
.Y(n_4983)
);

BUFx2_ASAP7_75t_L g4984 ( 
.A(n_4855),
.Y(n_4984)
);

OAI21x1_ASAP7_75t_L g4985 ( 
.A1(n_4661),
.A2(n_4535),
.B(n_4809),
.Y(n_4985)
);

AOI22xp33_ASAP7_75t_L g4986 ( 
.A1(n_4711),
.A2(n_4295),
.B1(n_4323),
.B2(n_4312),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_4677),
.A2(n_3388),
.B(n_3386),
.Y(n_4987)
);

AO31x2_ASAP7_75t_L g4988 ( 
.A1(n_4858),
.A2(n_4340),
.A3(n_4349),
.B(n_4327),
.Y(n_4988)
);

OAI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_4533),
.A2(n_1158),
.B(n_1155),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4528),
.B(n_1161),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_L g4991 ( 
.A1(n_4683),
.A2(n_3388),
.B(n_2924),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4552),
.A2(n_2924),
.B(n_2921),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4533),
.A2(n_4766),
.B(n_4565),
.Y(n_4993)
);

A2O1A1Ixp33_ASAP7_75t_L g4994 ( 
.A1(n_4707),
.A2(n_1164),
.B(n_1170),
.C(n_1161),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4560),
.A2(n_2934),
.B(n_2924),
.Y(n_4995)
);

OR2x2_ASAP7_75t_L g4996 ( 
.A(n_4548),
.B(n_1164),
.Y(n_4996)
);

OAI21x1_ASAP7_75t_L g4997 ( 
.A1(n_4810),
.A2(n_3351),
.B(n_3350),
.Y(n_4997)
);

AOI21xp33_ASAP7_75t_L g4998 ( 
.A1(n_4630),
.A2(n_1181),
.B(n_1170),
.Y(n_4998)
);

AND2x4_ASAP7_75t_L g4999 ( 
.A(n_4751),
.B(n_2934),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4546),
.B(n_1181),
.Y(n_5000)
);

OAI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_4630),
.A2(n_4779),
.B(n_4887),
.Y(n_5001)
);

A2O1A1Ixp33_ASAP7_75t_L g5002 ( 
.A1(n_4711),
.A2(n_1187),
.B(n_925),
.C(n_927),
.Y(n_5002)
);

OAI22xp5_ASAP7_75t_L g5003 ( 
.A1(n_4605),
.A2(n_1187),
.B1(n_819),
.B2(n_970),
.Y(n_5003)
);

OAI21x1_ASAP7_75t_L g5004 ( 
.A1(n_4713),
.A2(n_3357),
.B(n_3353),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_SL g5005 ( 
.A(n_4517),
.B(n_2235),
.Y(n_5005)
);

OAI21x1_ASAP7_75t_L g5006 ( 
.A1(n_4727),
.A2(n_3357),
.B(n_3353),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4549),
.B(n_911),
.Y(n_5007)
);

OAI22xp5_ASAP7_75t_L g5008 ( 
.A1(n_4640),
.A2(n_4554),
.B1(n_4539),
.B2(n_4641),
.Y(n_5008)
);

OAI22x1_ASAP7_75t_L g5009 ( 
.A1(n_4850),
.A2(n_923),
.B1(n_929),
.B2(n_922),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4566),
.B(n_911),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4592),
.B(n_911),
.Y(n_5011)
);

CKINVDCx11_ASAP7_75t_R g5012 ( 
.A(n_4588),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4598),
.B(n_911),
.Y(n_5013)
);

INVx1_ASAP7_75t_SL g5014 ( 
.A(n_4882),
.Y(n_5014)
);

INVx3_ASAP7_75t_L g5015 ( 
.A(n_4787),
.Y(n_5015)
);

OR2x2_ASAP7_75t_L g5016 ( 
.A(n_4664),
.B(n_911),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4568),
.B(n_911),
.Y(n_5017)
);

NAND3xp33_ASAP7_75t_L g5018 ( 
.A(n_4892),
.B(n_970),
.C(n_911),
.Y(n_5018)
);

AOI221xp5_ASAP7_75t_SL g5019 ( 
.A1(n_4780),
.A2(n_1059),
.B1(n_1065),
.B2(n_987),
.C(n_970),
.Y(n_5019)
);

OAI21x1_ASAP7_75t_L g5020 ( 
.A1(n_4749),
.A2(n_3365),
.B(n_3363),
.Y(n_5020)
);

INVx3_ASAP7_75t_L g5021 ( 
.A(n_4787),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4670),
.Y(n_5022)
);

A2O1A1Ixp33_ASAP7_75t_L g5023 ( 
.A1(n_4893),
.A2(n_930),
.B(n_933),
.C(n_928),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4559),
.B(n_970),
.Y(n_5024)
);

O2A1O1Ixp5_ASAP7_75t_L g5025 ( 
.A1(n_4650),
.A2(n_2235),
.B(n_2283),
.C(n_2270),
.Y(n_5025)
);

AND2x4_ASAP7_75t_L g5026 ( 
.A(n_4618),
.B(n_2934),
.Y(n_5026)
);

AOI21x1_ASAP7_75t_L g5027 ( 
.A1(n_4731),
.A2(n_2290),
.B(n_2286),
.Y(n_5027)
);

OAI21xp5_ASAP7_75t_L g5028 ( 
.A1(n_4612),
.A2(n_2273),
.B(n_2204),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4629),
.B(n_970),
.Y(n_5029)
);

AOI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4691),
.A2(n_2964),
.B(n_2950),
.Y(n_5030)
);

INVxp67_ASAP7_75t_SL g5031 ( 
.A(n_4725),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4626),
.B(n_4694),
.Y(n_5032)
);

OAI21x1_ASAP7_75t_L g5033 ( 
.A1(n_4754),
.A2(n_4764),
.B(n_4582),
.Y(n_5033)
);

INVx3_ASAP7_75t_L g5034 ( 
.A(n_4737),
.Y(n_5034)
);

BUFx2_ASAP7_75t_L g5035 ( 
.A(n_4826),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4746),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4693),
.A2(n_2964),
.B(n_2950),
.Y(n_5037)
);

OAI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4790),
.A2(n_2273),
.B(n_2206),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4812),
.B(n_970),
.Y(n_5039)
);

OAI21x1_ASAP7_75t_L g5040 ( 
.A1(n_4613),
.A2(n_3369),
.B(n_2480),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4753),
.Y(n_5041)
);

AND2x2_ASAP7_75t_L g5042 ( 
.A(n_4561),
.B(n_970),
.Y(n_5042)
);

AOI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4658),
.A2(n_2964),
.B(n_2950),
.Y(n_5043)
);

AOI21xp5_ASAP7_75t_L g5044 ( 
.A1(n_4659),
.A2(n_2966),
.B(n_2964),
.Y(n_5044)
);

A2O1A1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4747),
.A2(n_943),
.B(n_944),
.C(n_935),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4547),
.A2(n_2970),
.B(n_2966),
.Y(n_5046)
);

OAI21x1_ASAP7_75t_L g5047 ( 
.A1(n_4895),
.A2(n_3369),
.B(n_2480),
.Y(n_5047)
);

AOI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4518),
.A2(n_2970),
.B(n_2966),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4846),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4813),
.B(n_987),
.Y(n_5050)
);

INVx5_ASAP7_75t_L g5051 ( 
.A(n_4586),
.Y(n_5051)
);

OAI22xp5_ASAP7_75t_L g5052 ( 
.A1(n_4539),
.A2(n_4641),
.B1(n_4858),
.B2(n_4833),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4816),
.B(n_987),
.Y(n_5053)
);

AOI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4580),
.A2(n_2970),
.B(n_2966),
.Y(n_5054)
);

NAND2x1p5_ASAP7_75t_L g5055 ( 
.A(n_4586),
.B(n_3277),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4768),
.B(n_987),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4769),
.B(n_987),
.Y(n_5057)
);

AND2x6_ASAP7_75t_SL g5058 ( 
.A(n_4708),
.B(n_2270),
.Y(n_5058)
);

BUFx2_ASAP7_75t_L g5059 ( 
.A(n_4826),
.Y(n_5059)
);

BUFx4f_ASAP7_75t_L g5060 ( 
.A(n_4541),
.Y(n_5060)
);

OAI21x1_ASAP7_75t_L g5061 ( 
.A1(n_4574),
.A2(n_2480),
.B(n_3209),
.Y(n_5061)
);

OAI21x1_ASAP7_75t_L g5062 ( 
.A1(n_4755),
.A2(n_3210),
.B(n_3209),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4822),
.B(n_987),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4830),
.B(n_987),
.Y(n_5064)
);

BUFx6f_ASAP7_75t_L g5065 ( 
.A(n_4541),
.Y(n_5065)
);

AND2x2_ASAP7_75t_L g5066 ( 
.A(n_4674),
.B(n_1059),
.Y(n_5066)
);

OAI21x1_ASAP7_75t_L g5067 ( 
.A1(n_4522),
.A2(n_3216),
.B(n_3210),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4679),
.B(n_1059),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4845),
.B(n_1059),
.Y(n_5069)
);

OAI21xp33_ASAP7_75t_L g5070 ( 
.A1(n_4757),
.A2(n_1065),
.B(n_1059),
.Y(n_5070)
);

OAI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_4834),
.A2(n_2273),
.B(n_2184),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_SL g5072 ( 
.A(n_4517),
.B(n_2270),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4848),
.Y(n_5073)
);

AO21x1_ASAP7_75t_L g5074 ( 
.A1(n_4516),
.A2(n_4519),
.B(n_4623),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_SL g5075 ( 
.A(n_4597),
.B(n_2283),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_4821),
.B(n_1059),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4825),
.B(n_1059),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4663),
.B(n_1065),
.Y(n_5078)
);

BUFx6f_ASAP7_75t_L g5079 ( 
.A(n_4597),
.Y(n_5079)
);

AO31x2_ASAP7_75t_L g5080 ( 
.A1(n_4719),
.A2(n_2687),
.A3(n_2684),
.B(n_3290),
.Y(n_5080)
);

OAI21x1_ASAP7_75t_SL g5081 ( 
.A1(n_4648),
.A2(n_4611),
.B(n_4669),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4665),
.B(n_1065),
.Y(n_5082)
);

AO21x1_ASAP7_75t_L g5083 ( 
.A1(n_4687),
.A2(n_2283),
.B(n_2333),
.Y(n_5083)
);

INVx4_ASAP7_75t_L g5084 ( 
.A(n_4778),
.Y(n_5084)
);

OAI21x1_ASAP7_75t_L g5085 ( 
.A1(n_4852),
.A2(n_3226),
.B(n_3221),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4860),
.Y(n_5086)
);

OAI21x1_ASAP7_75t_L g5087 ( 
.A1(n_4660),
.A2(n_4789),
.B(n_4777),
.Y(n_5087)
);

BUFx6f_ASAP7_75t_L g5088 ( 
.A(n_4597),
.Y(n_5088)
);

BUFx3_ASAP7_75t_L g5089 ( 
.A(n_4696),
.Y(n_5089)
);

BUFx4_ASAP7_75t_SL g5090 ( 
.A(n_4562),
.Y(n_5090)
);

AO31x2_ASAP7_75t_L g5091 ( 
.A1(n_4596),
.A2(n_2687),
.A3(n_2684),
.B(n_3290),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4772),
.A2(n_2992),
.B(n_2971),
.Y(n_5092)
);

OAI21xp5_ASAP7_75t_L g5093 ( 
.A1(n_4835),
.A2(n_2368),
.B(n_2246),
.Y(n_5093)
);

NAND3xp33_ASAP7_75t_L g5094 ( 
.A(n_4878),
.B(n_1068),
.C(n_1065),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4712),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4530),
.Y(n_5096)
);

AOI21x1_ASAP7_75t_L g5097 ( 
.A1(n_4827),
.A2(n_2308),
.B(n_2302),
.Y(n_5097)
);

NAND2x1_ASAP7_75t_L g5098 ( 
.A(n_4728),
.B(n_3119),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4595),
.Y(n_5099)
);

OAI22xp5_ASAP7_75t_SL g5100 ( 
.A1(n_4555),
.A2(n_949),
.B1(n_957),
.B2(n_947),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4616),
.Y(n_5101)
);

OAI21xp5_ASAP7_75t_L g5102 ( 
.A1(n_4676),
.A2(n_4831),
.B(n_4784),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4775),
.B(n_1065),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4729),
.B(n_1065),
.Y(n_5104)
);

NAND3xp33_ASAP7_75t_L g5105 ( 
.A(n_4897),
.B(n_1097),
.C(n_1068),
.Y(n_5105)
);

INVxp67_ASAP7_75t_L g5106 ( 
.A(n_4690),
.Y(n_5106)
);

NOR2xp33_ASAP7_75t_L g5107 ( 
.A(n_4732),
.B(n_35),
.Y(n_5107)
);

OAI21xp5_ASAP7_75t_L g5108 ( 
.A1(n_4842),
.A2(n_2368),
.B(n_2269),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4621),
.Y(n_5109)
);

INVx4_ASAP7_75t_L g5110 ( 
.A(n_4604),
.Y(n_5110)
);

BUFx4_ASAP7_75t_SL g5111 ( 
.A(n_4774),
.Y(n_5111)
);

INVx1_ASAP7_75t_SL g5112 ( 
.A(n_4867),
.Y(n_5112)
);

INVx4_ASAP7_75t_L g5113 ( 
.A(n_4604),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_SL g5114 ( 
.A(n_4806),
.B(n_2992),
.Y(n_5114)
);

OAI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_4899),
.A2(n_2368),
.B(n_2274),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_4721),
.B(n_1068),
.Y(n_5116)
);

INVx5_ASAP7_75t_L g5117 ( 
.A(n_4586),
.Y(n_5117)
);

OAI21x1_ASAP7_75t_L g5118 ( 
.A1(n_4843),
.A2(n_3236),
.B(n_2612),
.Y(n_5118)
);

OAI21x1_ASAP7_75t_L g5119 ( 
.A1(n_4844),
.A2(n_2612),
.B(n_2605),
.Y(n_5119)
);

AOI22xp33_ASAP7_75t_L g5120 ( 
.A1(n_4526),
.A2(n_2076),
.B1(n_2932),
.B2(n_2922),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4794),
.B(n_1068),
.Y(n_5121)
);

A2O1A1Ixp33_ASAP7_75t_L g5122 ( 
.A1(n_4631),
.A2(n_959),
.B(n_962),
.C(n_958),
.Y(n_5122)
);

AOI21x1_ASAP7_75t_L g5123 ( 
.A1(n_4636),
.A2(n_2315),
.B(n_2312),
.Y(n_5123)
);

AOI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_4564),
.A2(n_2996),
.B(n_2994),
.Y(n_5124)
);

AOI21xp5_ASAP7_75t_L g5125 ( 
.A1(n_4564),
.A2(n_2996),
.B(n_2994),
.Y(n_5125)
);

A2O1A1Ixp33_ASAP7_75t_L g5126 ( 
.A1(n_4798),
.A2(n_968),
.B(n_971),
.C(n_964),
.Y(n_5126)
);

AOI221xp5_ASAP7_75t_SL g5127 ( 
.A1(n_4622),
.A2(n_1102),
.B1(n_1131),
.B2(n_1097),
.C(n_1068),
.Y(n_5127)
);

INVx4_ASAP7_75t_L g5128 ( 
.A(n_4604),
.Y(n_5128)
);

AOI221xp5_ASAP7_75t_SL g5129 ( 
.A1(n_4807),
.A2(n_1102),
.B1(n_1131),
.B2(n_1097),
.C(n_1068),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4625),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_L g5131 ( 
.A(n_4638),
.B(n_4733),
.Y(n_5131)
);

INVx2_ASAP7_75t_SL g5132 ( 
.A(n_4583),
.Y(n_5132)
);

OAI21xp5_ASAP7_75t_L g5133 ( 
.A1(n_4801),
.A2(n_2292),
.B(n_2219),
.Y(n_5133)
);

O2A1O1Ixp5_ASAP7_75t_L g5134 ( 
.A1(n_4714),
.A2(n_2315),
.B(n_2312),
.C(n_2996),
.Y(n_5134)
);

A2O1A1Ixp33_ASAP7_75t_L g5135 ( 
.A1(n_4861),
.A2(n_974),
.B(n_976),
.C(n_972),
.Y(n_5135)
);

CKINVDCx5p33_ASAP7_75t_R g5136 ( 
.A(n_4550),
.Y(n_5136)
);

OAI21x1_ASAP7_75t_SL g5137 ( 
.A1(n_4590),
.A2(n_2317),
.B(n_2074),
.Y(n_5137)
);

AOI21xp5_ASAP7_75t_L g5138 ( 
.A1(n_4656),
.A2(n_3028),
.B(n_3021),
.Y(n_5138)
);

NOR2xp33_ASAP7_75t_L g5139 ( 
.A(n_4781),
.B(n_35),
.Y(n_5139)
);

NAND3xp33_ASAP7_75t_L g5140 ( 
.A(n_4870),
.B(n_1097),
.C(n_1068),
.Y(n_5140)
);

AO21x2_ASAP7_75t_L g5141 ( 
.A1(n_4773),
.A2(n_2677),
.B(n_2672),
.Y(n_5141)
);

OAI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_4756),
.A2(n_2076),
.B(n_2768),
.Y(n_5142)
);

AND2x4_ASAP7_75t_L g5143 ( 
.A(n_4572),
.B(n_3021),
.Y(n_5143)
);

OAI21x1_ASAP7_75t_L g5144 ( 
.A1(n_4869),
.A2(n_2652),
.B(n_2648),
.Y(n_5144)
);

A2O1A1Ixp33_ASAP7_75t_L g5145 ( 
.A1(n_4865),
.A2(n_980),
.B(n_981),
.C(n_979),
.Y(n_5145)
);

BUFx2_ASAP7_75t_L g5146 ( 
.A(n_4682),
.Y(n_5146)
);

OAI21x1_ASAP7_75t_L g5147 ( 
.A1(n_4871),
.A2(n_2652),
.B(n_2648),
.Y(n_5147)
);

A2O1A1Ixp33_ASAP7_75t_L g5148 ( 
.A1(n_4536),
.A2(n_983),
.B(n_984),
.C(n_982),
.Y(n_5148)
);

AOI21xp5_ASAP7_75t_L g5149 ( 
.A1(n_4836),
.A2(n_3028),
.B(n_3021),
.Y(n_5149)
);

OAI22xp5_ASAP7_75t_L g5150 ( 
.A1(n_4686),
.A2(n_1102),
.B1(n_1131),
.B2(n_1097),
.Y(n_5150)
);

OAI21x1_ASAP7_75t_L g5151 ( 
.A1(n_4606),
.A2(n_4577),
.B(n_4576),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_4617),
.B(n_1097),
.Y(n_5152)
);

AND2x2_ASAP7_75t_L g5153 ( 
.A(n_4849),
.B(n_1097),
.Y(n_5153)
);

OAI21xp33_ASAP7_75t_SL g5154 ( 
.A1(n_4717),
.A2(n_4688),
.B(n_4854),
.Y(n_5154)
);

AO31x2_ASAP7_75t_L g5155 ( 
.A1(n_4678),
.A2(n_3308),
.A3(n_3313),
.B(n_3292),
.Y(n_5155)
);

BUFx6f_ASAP7_75t_L g5156 ( 
.A(n_4806),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4662),
.Y(n_5157)
);

CKINVDCx16_ASAP7_75t_R g5158 ( 
.A(n_4786),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4738),
.B(n_1102),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_4523),
.Y(n_5160)
);

CKINVDCx11_ASAP7_75t_R g5161 ( 
.A(n_4607),
.Y(n_5161)
);

A2O1A1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_4705),
.A2(n_986),
.B(n_988),
.C(n_985),
.Y(n_5162)
);

OAI21xp5_ASAP7_75t_L g5163 ( 
.A1(n_4756),
.A2(n_2076),
.B(n_2768),
.Y(n_5163)
);

AOI221x1_ASAP7_75t_L g5164 ( 
.A1(n_4873),
.A2(n_1152),
.B1(n_1191),
.B2(n_1131),
.C(n_1102),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4675),
.Y(n_5165)
);

AOI21x1_ASAP7_75t_SL g5166 ( 
.A1(n_4877),
.A2(n_2222),
.B(n_7),
.Y(n_5166)
);

OAI22xp5_ASAP7_75t_L g5167 ( 
.A1(n_4891),
.A2(n_1131),
.B1(n_1152),
.B2(n_1102),
.Y(n_5167)
);

AND2x6_ASAP7_75t_L g5168 ( 
.A(n_4572),
.B(n_3031),
.Y(n_5168)
);

INVx8_ASAP7_75t_L g5169 ( 
.A(n_4728),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_4748),
.B(n_1131),
.Y(n_5170)
);

NOR2x1p5_ASAP7_75t_SL g5171 ( 
.A(n_4632),
.B(n_2659),
.Y(n_5171)
);

AOI21x1_ASAP7_75t_L g5172 ( 
.A1(n_4762),
.A2(n_2075),
.B(n_2073),
.Y(n_5172)
);

OAI21x1_ASAP7_75t_SL g5173 ( 
.A1(n_4872),
.A2(n_2079),
.B(n_2078),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4699),
.Y(n_5174)
);

BUFx2_ASAP7_75t_L g5175 ( 
.A(n_4743),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4853),
.B(n_1131),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_L g5177 ( 
.A1(n_4770),
.A2(n_2659),
.B(n_3031),
.Y(n_5177)
);

OAI21x1_ASAP7_75t_L g5178 ( 
.A1(n_4770),
.A2(n_3086),
.B(n_3031),
.Y(n_5178)
);

OAI21x1_ASAP7_75t_L g5179 ( 
.A1(n_4859),
.A2(n_3086),
.B(n_3031),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_SL g5180 ( 
.A(n_4642),
.B(n_3086),
.Y(n_5180)
);

AOI21x1_ASAP7_75t_L g5181 ( 
.A1(n_4879),
.A2(n_4735),
.B(n_4771),
.Y(n_5181)
);

OA22x2_ASAP7_75t_L g5182 ( 
.A1(n_4532),
.A2(n_3068),
.B1(n_3128),
.B2(n_3000),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_SL g5183 ( 
.A1(n_4600),
.A2(n_3128),
.B(n_3068),
.Y(n_5183)
);

AO221x2_ASAP7_75t_L g5184 ( 
.A1(n_4698),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.C(n_11),
.Y(n_5184)
);

O2A1O1Ixp5_ASAP7_75t_L g5185 ( 
.A1(n_4862),
.A2(n_3110),
.B(n_3133),
.C(n_3086),
.Y(n_5185)
);

OAI21x1_ASAP7_75t_L g5186 ( 
.A1(n_4859),
.A2(n_3133),
.B(n_3110),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_SL g5187 ( 
.A1(n_4563),
.A2(n_2777),
.B(n_2776),
.Y(n_5187)
);

AOI21x1_ASAP7_75t_SL g5188 ( 
.A1(n_4639),
.A2(n_2222),
.B(n_9),
.Y(n_5188)
);

BUFx6f_ASAP7_75t_L g5189 ( 
.A(n_4642),
.Y(n_5189)
);

AOI21xp5_ASAP7_75t_L g5190 ( 
.A1(n_4840),
.A2(n_3133),
.B(n_3110),
.Y(n_5190)
);

OAI21x1_ASAP7_75t_SL g5191 ( 
.A1(n_4722),
.A2(n_2091),
.B(n_2087),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_4736),
.Y(n_5192)
);

AOI221x1_ASAP7_75t_L g5193 ( 
.A1(n_4876),
.A2(n_1191),
.B1(n_1152),
.B2(n_3133),
.C(n_3110),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_4745),
.Y(n_5194)
);

A2O1A1Ixp33_ASAP7_75t_L g5195 ( 
.A1(n_4649),
.A2(n_990),
.B(n_992),
.C(n_989),
.Y(n_5195)
);

HB1xp67_ASAP7_75t_L g5196 ( 
.A(n_4782),
.Y(n_5196)
);

AOI21x1_ASAP7_75t_L g5197 ( 
.A1(n_4783),
.A2(n_2100),
.B(n_2096),
.Y(n_5197)
);

AO21x2_ASAP7_75t_L g5198 ( 
.A1(n_4695),
.A2(n_2677),
.B(n_2672),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_4856),
.B(n_1152),
.Y(n_5199)
);

AOI21xp5_ASAP7_75t_L g5200 ( 
.A1(n_4668),
.A2(n_3199),
.B(n_3137),
.Y(n_5200)
);

INVxp67_ASAP7_75t_L g5201 ( 
.A(n_4819),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_4761),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4857),
.B(n_1152),
.Y(n_5203)
);

AND2x4_ASAP7_75t_L g5204 ( 
.A(n_4866),
.B(n_3137),
.Y(n_5204)
);

OAI21x1_ASAP7_75t_L g5205 ( 
.A1(n_4868),
.A2(n_3199),
.B(n_3137),
.Y(n_5205)
);

AOI21xp5_ASAP7_75t_L g5206 ( 
.A1(n_4697),
.A2(n_4710),
.B(n_4847),
.Y(n_5206)
);

OAI22xp5_ASAP7_75t_L g5207 ( 
.A1(n_4767),
.A2(n_1191),
.B1(n_1152),
.B2(n_997),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_4874),
.B(n_11),
.Y(n_5208)
);

OAI21x1_ASAP7_75t_L g5209 ( 
.A1(n_4868),
.A2(n_3206),
.B(n_3199),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_4886),
.B(n_789),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_4886),
.B(n_789),
.Y(n_5211)
);

NOR2xp33_ASAP7_75t_L g5212 ( 
.A(n_4838),
.B(n_36),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_4828),
.Y(n_5213)
);

BUFx3_ASAP7_75t_L g5214 ( 
.A(n_4639),
.Y(n_5214)
);

AOI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_4558),
.A2(n_3206),
.B(n_3199),
.Y(n_5215)
);

AO31x2_ASAP7_75t_L g5216 ( 
.A1(n_4680),
.A2(n_3308),
.A3(n_3313),
.B(n_3292),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_4875),
.B(n_996),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_4898),
.B(n_789),
.Y(n_5218)
);

OAI21xp5_ASAP7_75t_L g5219 ( 
.A1(n_4720),
.A2(n_2076),
.B(n_2776),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_4885),
.B(n_998),
.Y(n_5220)
);

INVx5_ASAP7_75t_L g5221 ( 
.A(n_4728),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4718),
.Y(n_5222)
);

INVx2_ASAP7_75t_SL g5223 ( 
.A(n_4724),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4896),
.B(n_12),
.Y(n_5224)
);

AOI21xp5_ASAP7_75t_L g5225 ( 
.A1(n_4824),
.A2(n_3249),
.B(n_3240),
.Y(n_5225)
);

BUFx6f_ASAP7_75t_L g5226 ( 
.A(n_4647),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_4900),
.B(n_1002),
.Y(n_5227)
);

OA21x2_ASAP7_75t_L g5228 ( 
.A1(n_4594),
.A2(n_3323),
.B(n_3316),
.Y(n_5228)
);

BUFx12f_ASAP7_75t_L g5229 ( 
.A(n_4726),
.Y(n_5229)
);

NAND2x1p5_ASAP7_75t_L g5230 ( 
.A(n_4645),
.B(n_3249),
.Y(n_5230)
);

AOI21xp5_ASAP7_75t_L g5231 ( 
.A1(n_4823),
.A2(n_3281),
.B(n_3249),
.Y(n_5231)
);

OR2x2_ASAP7_75t_L g5232 ( 
.A(n_4667),
.B(n_13),
.Y(n_5232)
);

AND2x4_ASAP7_75t_L g5233 ( 
.A(n_4866),
.B(n_3281),
.Y(n_5233)
);

OAI21x1_ASAP7_75t_L g5234 ( 
.A1(n_4741),
.A2(n_3304),
.B(n_3281),
.Y(n_5234)
);

AOI21x1_ASAP7_75t_L g5235 ( 
.A1(n_4584),
.A2(n_2110),
.B(n_2105),
.Y(n_5235)
);

OAI21xp5_ASAP7_75t_L g5236 ( 
.A1(n_4602),
.A2(n_2076),
.B(n_2777),
.Y(n_5236)
);

INVx3_ASAP7_75t_L g5237 ( 
.A(n_4726),
.Y(n_5237)
);

AOI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_4692),
.A2(n_4837),
.B(n_4614),
.Y(n_5238)
);

AO31x2_ASAP7_75t_L g5239 ( 
.A1(n_4793),
.A2(n_3323),
.A3(n_3324),
.B(n_3316),
.Y(n_5239)
);

AND2x2_ASAP7_75t_L g5240 ( 
.A(n_4726),
.B(n_888),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_SL g5241 ( 
.A(n_4888),
.B(n_3304),
.Y(n_5241)
);

AOI21xp5_ASAP7_75t_L g5242 ( 
.A1(n_4692),
.A2(n_3306),
.B(n_3304),
.Y(n_5242)
);

INVx3_ASAP7_75t_L g5243 ( 
.A(n_4888),
.Y(n_5243)
);

BUFx2_ASAP7_75t_L g5244 ( 
.A(n_4743),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_4765),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_4837),
.A2(n_3306),
.B(n_3304),
.Y(n_5246)
);

AOI21xp5_ASAP7_75t_L g5247 ( 
.A1(n_4894),
.A2(n_3360),
.B(n_3306),
.Y(n_5247)
);

INVxp67_ASAP7_75t_SL g5248 ( 
.A(n_4901),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_4742),
.A2(n_2783),
.B(n_2781),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4802),
.B(n_1003),
.Y(n_5250)
);

NOR2xp33_ASAP7_75t_L g5251 ( 
.A(n_4715),
.B(n_36),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_4635),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4760),
.B(n_13),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_4804),
.B(n_15),
.Y(n_5254)
);

NAND2x1_ASAP7_75t_L g5255 ( 
.A(n_4728),
.B(n_3119),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_4570),
.Y(n_5256)
);

AOI21xp5_ASAP7_75t_L g5257 ( 
.A1(n_4894),
.A2(n_3384),
.B(n_3360),
.Y(n_5257)
);

NAND2xp5_ASAP7_75t_L g5258 ( 
.A(n_4805),
.B(n_15),
.Y(n_5258)
);

INVx3_ASAP7_75t_L g5259 ( 
.A(n_4888),
.Y(n_5259)
);

AOI21xp5_ASAP7_75t_L g5260 ( 
.A1(n_4791),
.A2(n_3384),
.B(n_3360),
.Y(n_5260)
);

OAI21x1_ASAP7_75t_L g5261 ( 
.A1(n_4544),
.A2(n_3384),
.B(n_2669),
.Y(n_5261)
);

OAI22xp5_ASAP7_75t_L g5262 ( 
.A1(n_4593),
.A2(n_1009),
.B1(n_1012),
.B2(n_1011),
.Y(n_5262)
);

NOR3xp33_ASAP7_75t_L g5263 ( 
.A(n_4723),
.B(n_1016),
.C(n_1015),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4603),
.B(n_16),
.Y(n_5264)
);

AOI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_4601),
.A2(n_3384),
.B(n_2801),
.Y(n_5265)
);

OAI21xp5_ASAP7_75t_L g5266 ( 
.A1(n_4796),
.A2(n_2783),
.B(n_2781),
.Y(n_5266)
);

AND2x2_ASAP7_75t_L g5267 ( 
.A(n_4797),
.B(n_888),
.Y(n_5267)
);

INVx2_ASAP7_75t_L g5268 ( 
.A(n_4585),
.Y(n_5268)
);

OA21x2_ASAP7_75t_L g5269 ( 
.A1(n_5087),
.A2(n_4609),
.B(n_4701),
.Y(n_5269)
);

OAI21x1_ASAP7_75t_L g5270 ( 
.A1(n_4909),
.A2(n_4889),
.B(n_4703),
.Y(n_5270)
);

OAI21x1_ASAP7_75t_L g5271 ( 
.A1(n_5206),
.A2(n_4889),
.B(n_4702),
.Y(n_5271)
);

INVxp67_ASAP7_75t_L g5272 ( 
.A(n_4982),
.Y(n_5272)
);

AOI22xp5_ASAP7_75t_L g5273 ( 
.A1(n_4908),
.A2(n_4651),
.B1(n_4587),
.B2(n_4881),
.Y(n_5273)
);

OAI22xp5_ASAP7_75t_L g5274 ( 
.A1(n_4908),
.A2(n_4655),
.B1(n_4883),
.B2(n_4788),
.Y(n_5274)
);

BUFx8_ASAP7_75t_L g5275 ( 
.A(n_5132),
.Y(n_5275)
);

AO22x1_ASAP7_75t_L g5276 ( 
.A1(n_5112),
.A2(n_4785),
.B1(n_4884),
.B2(n_4645),
.Y(n_5276)
);

OAI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_4915),
.A2(n_4644),
.B(n_4589),
.Y(n_5277)
);

OR2x2_ASAP7_75t_L g5278 ( 
.A(n_5014),
.B(n_4758),
.Y(n_5278)
);

INVx2_ASAP7_75t_L g5279 ( 
.A(n_5049),
.Y(n_5279)
);

AND2x4_ASAP7_75t_L g5280 ( 
.A(n_4984),
.B(n_4811),
.Y(n_5280)
);

AO21x2_ASAP7_75t_L g5281 ( 
.A1(n_4949),
.A2(n_4657),
.B(n_2198),
.Y(n_5281)
);

AOI22xp5_ASAP7_75t_L g5282 ( 
.A1(n_5052),
.A2(n_4808),
.B1(n_4785),
.B2(n_4776),
.Y(n_5282)
);

OAI21x1_ASAP7_75t_L g5283 ( 
.A1(n_5151),
.A2(n_4815),
.B(n_4776),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_5052),
.A2(n_4706),
.B(n_4815),
.Y(n_5284)
);

AOI21xp5_ASAP7_75t_L g5285 ( 
.A1(n_4949),
.A2(n_4706),
.B(n_2797),
.Y(n_5285)
);

AND2x4_ASAP7_75t_L g5286 ( 
.A(n_4910),
.B(n_4785),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_5014),
.B(n_16),
.Y(n_5287)
);

INVxp67_ASAP7_75t_L g5288 ( 
.A(n_4918),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4913),
.Y(n_5289)
);

NAND3xp33_ASAP7_75t_L g5290 ( 
.A(n_4955),
.B(n_4652),
.C(n_4880),
.Y(n_5290)
);

INVxp67_ASAP7_75t_SL g5291 ( 
.A(n_5074),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4932),
.Y(n_5292)
);

AOI21x1_ASAP7_75t_L g5293 ( 
.A1(n_5017),
.A2(n_2200),
.B(n_2114),
.Y(n_5293)
);

OR2x2_ASAP7_75t_L g5294 ( 
.A(n_4933),
.B(n_16),
.Y(n_5294)
);

AOI21xp5_ASAP7_75t_L g5295 ( 
.A1(n_4966),
.A2(n_2797),
.B(n_2786),
.Y(n_5295)
);

OAI21x1_ASAP7_75t_L g5296 ( 
.A1(n_5033),
.A2(n_2640),
.B(n_2483),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4962),
.B(n_1017),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4966),
.A2(n_2803),
.B(n_2786),
.Y(n_5298)
);

OA21x2_ASAP7_75t_L g5299 ( 
.A1(n_4943),
.A2(n_1020),
.B(n_1019),
.Y(n_5299)
);

OAI21x1_ASAP7_75t_L g5300 ( 
.A1(n_4979),
.A2(n_2640),
.B(n_2483),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_4976),
.B(n_1029),
.Y(n_5301)
);

BUFx4_ASAP7_75t_SL g5302 ( 
.A(n_4972),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_4981),
.Y(n_5303)
);

NOR2xp67_ASAP7_75t_SL g5304 ( 
.A(n_5221),
.B(n_5140),
.Y(n_5304)
);

INVx6_ASAP7_75t_L g5305 ( 
.A(n_4977),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_4976),
.B(n_4906),
.Y(n_5306)
);

AND2x2_ASAP7_75t_L g5307 ( 
.A(n_4914),
.B(n_17),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_4943),
.Y(n_5308)
);

CKINVDCx11_ASAP7_75t_R g5309 ( 
.A(n_5161),
.Y(n_5309)
);

INVx3_ASAP7_75t_L g5310 ( 
.A(n_4946),
.Y(n_5310)
);

AO31x2_ASAP7_75t_L g5311 ( 
.A1(n_4917),
.A2(n_3331),
.A3(n_3332),
.B(n_3324),
.Y(n_5311)
);

OR2x2_ASAP7_75t_L g5312 ( 
.A(n_5196),
.B(n_17),
.Y(n_5312)
);

OAI21x1_ASAP7_75t_L g5313 ( 
.A1(n_5027),
.A2(n_2640),
.B(n_2483),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5022),
.Y(n_5314)
);

OAI21x1_ASAP7_75t_L g5315 ( 
.A1(n_4985),
.A2(n_2485),
.B(n_2471),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_4951),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5036),
.Y(n_5317)
);

HB1xp67_ASAP7_75t_L g5318 ( 
.A(n_4944),
.Y(n_5318)
);

OAI21x1_ASAP7_75t_L g5319 ( 
.A1(n_5137),
.A2(n_2485),
.B(n_2471),
.Y(n_5319)
);

OR2x2_ASAP7_75t_L g5320 ( 
.A(n_5032),
.B(n_18),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_4906),
.B(n_1030),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_L g5322 ( 
.A(n_5131),
.B(n_37),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_4974),
.B(n_1035),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_4946),
.B(n_18),
.Y(n_5324)
);

AO31x2_ASAP7_75t_L g5325 ( 
.A1(n_4940),
.A2(n_3332),
.A3(n_3335),
.B(n_3331),
.Y(n_5325)
);

NOR2xp33_ASAP7_75t_L g5326 ( 
.A(n_4971),
.B(n_37),
.Y(n_5326)
);

INVx1_ASAP7_75t_SL g5327 ( 
.A(n_5111),
.Y(n_5327)
);

NOR2xp33_ASAP7_75t_R g5328 ( 
.A(n_5136),
.B(n_40),
.Y(n_5328)
);

AOI21xp5_ASAP7_75t_L g5329 ( 
.A1(n_5008),
.A2(n_2804),
.B(n_2803),
.Y(n_5329)
);

O2A1O1Ixp5_ASAP7_75t_L g5330 ( 
.A1(n_4903),
.A2(n_2804),
.B(n_2811),
.C(n_2807),
.Y(n_5330)
);

NAND3x1_ASAP7_75t_L g5331 ( 
.A(n_4960),
.B(n_2236),
.C(n_2233),
.Y(n_5331)
);

BUFx6f_ASAP7_75t_L g5332 ( 
.A(n_5229),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_4956),
.B(n_5015),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_5031),
.B(n_1038),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_5041),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_5073),
.Y(n_5336)
);

CKINVDCx20_ASAP7_75t_R g5337 ( 
.A(n_5012),
.Y(n_5337)
);

CKINVDCx9p33_ASAP7_75t_R g5338 ( 
.A(n_5035),
.Y(n_5338)
);

INVx3_ASAP7_75t_L g5339 ( 
.A(n_4956),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5086),
.Y(n_5340)
);

BUFx2_ASAP7_75t_L g5341 ( 
.A(n_5146),
.Y(n_5341)
);

AOI21xp5_ASAP7_75t_L g5342 ( 
.A1(n_5008),
.A2(n_2811),
.B(n_2807),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_SL g5343 ( 
.A(n_5221),
.B(n_888),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_4953),
.B(n_1040),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_4947),
.Y(n_5345)
);

OAI21xp5_ASAP7_75t_L g5346 ( 
.A1(n_4915),
.A2(n_1045),
.B(n_1044),
.Y(n_5346)
);

AOI21xp5_ASAP7_75t_L g5347 ( 
.A1(n_5071),
.A2(n_2829),
.B(n_2812),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_4953),
.B(n_1047),
.Y(n_5348)
);

OAI21x1_ASAP7_75t_L g5349 ( 
.A1(n_5185),
.A2(n_2490),
.B(n_2488),
.Y(n_5349)
);

NAND2xp5_ASAP7_75t_SL g5350 ( 
.A(n_5221),
.B(n_888),
.Y(n_5350)
);

OAI21x1_ASAP7_75t_L g5351 ( 
.A1(n_5182),
.A2(n_2490),
.B(n_2488),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_SL g5352 ( 
.A(n_5154),
.B(n_1021),
.Y(n_5352)
);

NOR2xp33_ASAP7_75t_L g5353 ( 
.A(n_5089),
.B(n_38),
.Y(n_5353)
);

AOI221xp5_ASAP7_75t_L g5354 ( 
.A1(n_4965),
.A2(n_1050),
.B1(n_1060),
.B2(n_1056),
.C(n_1048),
.Y(n_5354)
);

NOR2x1_ASAP7_75t_L g5355 ( 
.A(n_5112),
.B(n_2663),
.Y(n_5355)
);

OAI21x1_ASAP7_75t_L g5356 ( 
.A1(n_5182),
.A2(n_4937),
.B(n_4904),
.Y(n_5356)
);

INVx5_ASAP7_75t_L g5357 ( 
.A(n_5059),
.Y(n_5357)
);

NAND2xp5_ASAP7_75t_L g5358 ( 
.A(n_5248),
.B(n_1061),
.Y(n_5358)
);

OAI21xp5_ASAP7_75t_L g5359 ( 
.A1(n_5002),
.A2(n_1066),
.B(n_1063),
.Y(n_5359)
);

OAI21xp5_ASAP7_75t_L g5360 ( 
.A1(n_4902),
.A2(n_1078),
.B(n_1071),
.Y(n_5360)
);

OAI21x1_ASAP7_75t_L g5361 ( 
.A1(n_5181),
.A2(n_2504),
.B(n_2678),
.Y(n_5361)
);

NAND2xp33_ASAP7_75t_L g5362 ( 
.A(n_5169),
.B(n_1082),
.Y(n_5362)
);

AOI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_4924),
.A2(n_4925),
.B1(n_5184),
.B2(n_5070),
.Y(n_5363)
);

BUFx10_ASAP7_75t_L g5364 ( 
.A(n_5160),
.Y(n_5364)
);

AOI21xp33_ASAP7_75t_L g5365 ( 
.A1(n_4905),
.A2(n_1084),
.B(n_1083),
.Y(n_5365)
);

AOI21xp5_ASAP7_75t_L g5366 ( 
.A1(n_5071),
.A2(n_2829),
.B(n_2812),
.Y(n_5366)
);

INVx3_ASAP7_75t_L g5367 ( 
.A(n_5021),
.Y(n_5367)
);

AOI21x1_ASAP7_75t_SL g5368 ( 
.A1(n_5264),
.A2(n_19),
.B(n_20),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_SL g5369 ( 
.A(n_4958),
.B(n_1021),
.Y(n_5369)
);

AOI221x1_ASAP7_75t_L g5370 ( 
.A1(n_4965),
.A2(n_1362),
.B1(n_1447),
.B2(n_1267),
.C(n_1229),
.Y(n_5370)
);

BUFx6f_ASAP7_75t_SL g5371 ( 
.A(n_5214),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_SL g5372 ( 
.A(n_5034),
.B(n_1021),
.Y(n_5372)
);

OAI21x1_ASAP7_75t_L g5373 ( 
.A1(n_4927),
.A2(n_2504),
.B(n_2686),
.Y(n_5373)
);

AO22x2_ASAP7_75t_L g5374 ( 
.A1(n_5222),
.A2(n_5245),
.B1(n_5096),
.B2(n_5095),
.Y(n_5374)
);

OAI21x1_ASAP7_75t_L g5375 ( 
.A1(n_4923),
.A2(n_2504),
.B(n_2686),
.Y(n_5375)
);

AOI22xp5_ASAP7_75t_L g5376 ( 
.A1(n_4925),
.A2(n_1073),
.B1(n_1093),
.B2(n_1021),
.Y(n_5376)
);

OAI21x1_ASAP7_75t_SL g5377 ( 
.A1(n_5081),
.A2(n_19),
.B(n_21),
.Y(n_5377)
);

OAI21xp5_ASAP7_75t_L g5378 ( 
.A1(n_5251),
.A2(n_1087),
.B(n_1086),
.Y(n_5378)
);

AOI21xp5_ASAP7_75t_L g5379 ( 
.A1(n_4993),
.A2(n_2833),
.B(n_2830),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_4921),
.A2(n_2935),
.B(n_2932),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5213),
.Y(n_5381)
);

OAI21x1_ASAP7_75t_L g5382 ( 
.A1(n_4941),
.A2(n_2937),
.B(n_2935),
.Y(n_5382)
);

NAND2xp5_ASAP7_75t_SL g5383 ( 
.A(n_5034),
.B(n_1021),
.Y(n_5383)
);

AOI221xp5_ASAP7_75t_SL g5384 ( 
.A1(n_5107),
.A2(n_5212),
.B1(n_5139),
.B2(n_5148),
.C(n_4922),
.Y(n_5384)
);

OAI21xp5_ASAP7_75t_L g5385 ( 
.A1(n_5140),
.A2(n_1094),
.B(n_1089),
.Y(n_5385)
);

OAI21x1_ASAP7_75t_L g5386 ( 
.A1(n_4911),
.A2(n_2941),
.B(n_2937),
.Y(n_5386)
);

BUFx6f_ASAP7_75t_L g5387 ( 
.A(n_5189),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_5252),
.Y(n_5388)
);

NAND2xp5_ASAP7_75t_SL g5389 ( 
.A(n_4973),
.B(n_1073),
.Y(n_5389)
);

NOR2xp33_ASAP7_75t_L g5390 ( 
.A(n_5201),
.B(n_39),
.Y(n_5390)
);

AND2x4_ASAP7_75t_L g5391 ( 
.A(n_4919),
.B(n_19),
.Y(n_5391)
);

NOR2xp33_ASAP7_75t_L g5392 ( 
.A(n_5223),
.B(n_39),
.Y(n_5392)
);

AO31x2_ASAP7_75t_L g5393 ( 
.A1(n_5083),
.A2(n_3336),
.A3(n_3337),
.B(n_3335),
.Y(n_5393)
);

NOR2x1_ASAP7_75t_SL g5394 ( 
.A(n_5051),
.B(n_2830),
.Y(n_5394)
);

AND2x4_ASAP7_75t_L g5395 ( 
.A(n_4931),
.B(n_21),
.Y(n_5395)
);

OR2x2_ASAP7_75t_L g5396 ( 
.A(n_5106),
.B(n_23),
.Y(n_5396)
);

INVxp67_ASAP7_75t_L g5397 ( 
.A(n_4990),
.Y(n_5397)
);

AOI21xp5_ASAP7_75t_L g5398 ( 
.A1(n_4993),
.A2(n_2835),
.B(n_2833),
.Y(n_5398)
);

NOR4xp25_ASAP7_75t_L g5399 ( 
.A(n_5000),
.B(n_1093),
.C(n_1073),
.D(n_25),
.Y(n_5399)
);

CKINVDCx14_ASAP7_75t_R g5400 ( 
.A(n_5090),
.Y(n_5400)
);

AND2x2_ASAP7_75t_L g5401 ( 
.A(n_4934),
.B(n_23),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4939),
.Y(n_5402)
);

OA21x2_ASAP7_75t_L g5403 ( 
.A1(n_5024),
.A2(n_1103),
.B(n_1096),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5010),
.B(n_1107),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_5038),
.A2(n_2836),
.B(n_2835),
.Y(n_5405)
);

NAND3x1_ASAP7_75t_L g5406 ( 
.A(n_4907),
.B(n_23),
.C(n_24),
.Y(n_5406)
);

NOR2xp33_ASAP7_75t_L g5407 ( 
.A(n_5158),
.B(n_41),
.Y(n_5407)
);

NAND2xp5_ASAP7_75t_L g5408 ( 
.A(n_5011),
.B(n_1109),
.Y(n_5408)
);

AOI21xp5_ASAP7_75t_L g5409 ( 
.A1(n_5038),
.A2(n_2843),
.B(n_2836),
.Y(n_5409)
);

NOR2x1_ASAP7_75t_L g5410 ( 
.A(n_5029),
.B(n_2663),
.Y(n_5410)
);

AOI21xp5_ASAP7_75t_L g5411 ( 
.A1(n_5028),
.A2(n_2845),
.B(n_2843),
.Y(n_5411)
);

OAI21x1_ASAP7_75t_L g5412 ( 
.A1(n_4948),
.A2(n_2942),
.B(n_2941),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_5013),
.B(n_1111),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_4945),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5099),
.Y(n_5415)
);

OAI22xp5_ASAP7_75t_L g5416 ( 
.A1(n_5001),
.A2(n_4950),
.B1(n_5028),
.B2(n_5249),
.Y(n_5416)
);

AO31x2_ASAP7_75t_L g5417 ( 
.A1(n_5056),
.A2(n_3337),
.A3(n_3336),
.B(n_2944),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_L g5418 ( 
.A(n_5057),
.B(n_5063),
.Y(n_5418)
);

OAI21x1_ASAP7_75t_L g5419 ( 
.A1(n_4959),
.A2(n_2944),
.B(n_2942),
.Y(n_5419)
);

INVx2_ASAP7_75t_SL g5420 ( 
.A(n_4935),
.Y(n_5420)
);

BUFx6f_ASAP7_75t_L g5421 ( 
.A(n_5189),
.Y(n_5421)
);

AOI21xp5_ASAP7_75t_L g5422 ( 
.A1(n_5098),
.A2(n_2854),
.B(n_2845),
.Y(n_5422)
);

BUFx6f_ASAP7_75t_L g5423 ( 
.A(n_5189),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5101),
.Y(n_5424)
);

BUFx6f_ASAP7_75t_L g5425 ( 
.A(n_5226),
.Y(n_5425)
);

OAI21x1_ASAP7_75t_L g5426 ( 
.A1(n_4964),
.A2(n_2948),
.B(n_2945),
.Y(n_5426)
);

NAND3xp33_ASAP7_75t_SL g5427 ( 
.A(n_4963),
.B(n_1114),
.C(n_1113),
.Y(n_5427)
);

OAI21xp5_ASAP7_75t_L g5428 ( 
.A1(n_4970),
.A2(n_1116),
.B(n_1115),
.Y(n_5428)
);

AOI221x1_ASAP7_75t_L g5429 ( 
.A1(n_5009),
.A2(n_1362),
.B1(n_1447),
.B2(n_1267),
.C(n_1229),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_5064),
.B(n_1117),
.Y(n_5430)
);

A2O1A1Ixp33_ASAP7_75t_L g5431 ( 
.A1(n_5001),
.A2(n_1125),
.B(n_1150),
.C(n_1140),
.Y(n_5431)
);

OAI21x1_ASAP7_75t_L g5432 ( 
.A1(n_4978),
.A2(n_2948),
.B(n_2945),
.Y(n_5432)
);

NOR2x1_ASAP7_75t_SL g5433 ( 
.A(n_5051),
.B(n_2854),
.Y(n_5433)
);

OAI21xp5_ASAP7_75t_L g5434 ( 
.A1(n_4970),
.A2(n_1127),
.B(n_1120),
.Y(n_5434)
);

OAI21x1_ASAP7_75t_L g5435 ( 
.A1(n_5123),
.A2(n_5067),
.B(n_5238),
.Y(n_5435)
);

AOI21x1_ASAP7_75t_SL g5436 ( 
.A1(n_5208),
.A2(n_25),
.B(n_26),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_5184),
.A2(n_1093),
.B1(n_1073),
.B2(n_2222),
.Y(n_5437)
);

A2O1A1Ixp33_ASAP7_75t_L g5438 ( 
.A1(n_5129),
.A2(n_1146),
.B(n_1163),
.C(n_1130),
.Y(n_5438)
);

AOI221xp5_ASAP7_75t_SL g5439 ( 
.A1(n_5126),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_5439)
);

AND2x4_ASAP7_75t_L g5440 ( 
.A(n_4954),
.B(n_26),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5109),
.Y(n_5441)
);

AOI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_5129),
.A2(n_1093),
.B1(n_1073),
.B2(n_2307),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_5255),
.A2(n_4995),
.B(n_4992),
.Y(n_5443)
);

OAI21x1_ASAP7_75t_L g5444 ( 
.A1(n_4912),
.A2(n_2959),
.B(n_2949),
.Y(n_5444)
);

OAI21x1_ASAP7_75t_L g5445 ( 
.A1(n_5118),
.A2(n_2959),
.B(n_2949),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_L g5446 ( 
.A(n_5069),
.B(n_1128),
.Y(n_5446)
);

OAI21x1_ASAP7_75t_L g5447 ( 
.A1(n_5124),
.A2(n_2961),
.B(n_2960),
.Y(n_5447)
);

AOI21x1_ASAP7_75t_SL g5448 ( 
.A1(n_5224),
.A2(n_28),
.B(n_30),
.Y(n_5448)
);

AO31x2_ASAP7_75t_L g5449 ( 
.A1(n_5193),
.A2(n_2961),
.A3(n_2965),
.B(n_2960),
.Y(n_5449)
);

HB1xp67_ASAP7_75t_L g5450 ( 
.A(n_5016),
.Y(n_5450)
);

OAI22xp5_ASAP7_75t_L g5451 ( 
.A1(n_4950),
.A2(n_1129),
.B1(n_1137),
.B2(n_1135),
.Y(n_5451)
);

INVx3_ASAP7_75t_L g5452 ( 
.A(n_5051),
.Y(n_5452)
);

NOR2xp33_ASAP7_75t_R g5453 ( 
.A(n_5060),
.B(n_5156),
.Y(n_5453)
);

OAI21x1_ASAP7_75t_L g5454 ( 
.A1(n_5125),
.A2(n_2972),
.B(n_2965),
.Y(n_5454)
);

AO31x2_ASAP7_75t_L g5455 ( 
.A1(n_5150),
.A2(n_2974),
.A3(n_2983),
.B(n_2972),
.Y(n_5455)
);

AOI21xp5_ASAP7_75t_L g5456 ( 
.A1(n_5169),
.A2(n_2863),
.B(n_2857),
.Y(n_5456)
);

HB1xp67_ASAP7_75t_L g5457 ( 
.A(n_5175),
.Y(n_5457)
);

BUFx2_ASAP7_75t_L g5458 ( 
.A(n_5244),
.Y(n_5458)
);

CKINVDCx11_ASAP7_75t_R g5459 ( 
.A(n_5084),
.Y(n_5459)
);

O2A1O1Ixp33_ASAP7_75t_L g5460 ( 
.A1(n_4916),
.A2(n_2245),
.B(n_2254),
.C(n_2247),
.Y(n_5460)
);

BUFx5_ASAP7_75t_L g5461 ( 
.A(n_5168),
.Y(n_5461)
);

NOR2x1_ASAP7_75t_SL g5462 ( 
.A(n_5051),
.B(n_2857),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_5232),
.B(n_1138),
.Y(n_5463)
);

AO31x2_ASAP7_75t_L g5464 ( 
.A1(n_5150),
.A2(n_2983),
.A3(n_2989),
.B(n_2974),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_5007),
.B(n_1141),
.Y(n_5465)
);

OA22x2_ASAP7_75t_L g5466 ( 
.A1(n_5042),
.A2(n_1142),
.B1(n_1144),
.B2(n_1143),
.Y(n_5466)
);

INVx1_ASAP7_75t_SL g5467 ( 
.A(n_4961),
.Y(n_5467)
);

OA21x2_ASAP7_75t_L g5468 ( 
.A1(n_5039),
.A2(n_1148),
.B(n_1147),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_4945),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5157),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5165),
.Y(n_5471)
);

AOI21xp5_ASAP7_75t_L g5472 ( 
.A1(n_5169),
.A2(n_2865),
.B(n_2863),
.Y(n_5472)
);

AOI211x1_ASAP7_75t_L g5473 ( 
.A1(n_4998),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_5473)
);

AOI221x1_ASAP7_75t_L g5474 ( 
.A1(n_5253),
.A2(n_1267),
.B1(n_1470),
.B2(n_1447),
.C(n_1362),
.Y(n_5474)
);

NAND2xp5_ASAP7_75t_L g5475 ( 
.A(n_5254),
.B(n_1151),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5258),
.B(n_1154),
.Y(n_5476)
);

O2A1O1Ixp5_ASAP7_75t_L g5477 ( 
.A1(n_5207),
.A2(n_2868),
.B(n_2869),
.C(n_2865),
.Y(n_5477)
);

OAI21x1_ASAP7_75t_L g5478 ( 
.A1(n_4997),
.A2(n_2993),
.B(n_2989),
.Y(n_5478)
);

OR2x2_ASAP7_75t_L g5479 ( 
.A(n_4996),
.B(n_32),
.Y(n_5479)
);

OAI22xp5_ASAP7_75t_L g5480 ( 
.A1(n_5249),
.A2(n_1156),
.B1(n_1162),
.B2(n_1159),
.Y(n_5480)
);

AOI21xp5_ASAP7_75t_L g5481 ( 
.A1(n_4926),
.A2(n_2869),
.B(n_2868),
.Y(n_5481)
);

AOI21xp5_ASAP7_75t_L g5482 ( 
.A1(n_4930),
.A2(n_2881),
.B(n_2876),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5004),
.A2(n_2995),
.B(n_2993),
.Y(n_5483)
);

OA21x2_ASAP7_75t_L g5484 ( 
.A1(n_5039),
.A2(n_1169),
.B(n_1165),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_L g5485 ( 
.A(n_5050),
.B(n_1171),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_L g5486 ( 
.A1(n_5046),
.A2(n_2881),
.B(n_2876),
.Y(n_5486)
);

OAI22xp5_ASAP7_75t_L g5487 ( 
.A1(n_5018),
.A2(n_1172),
.B1(n_1174),
.B2(n_1173),
.Y(n_5487)
);

INVx3_ASAP7_75t_SL g5488 ( 
.A(n_5084),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5174),
.Y(n_5489)
);

AOI21x1_ASAP7_75t_L g5490 ( 
.A1(n_5078),
.A2(n_2256),
.B(n_2901),
.Y(n_5490)
);

OAI21x1_ASAP7_75t_L g5491 ( 
.A1(n_5006),
.A2(n_3002),
.B(n_2995),
.Y(n_5491)
);

INVx5_ASAP7_75t_L g5492 ( 
.A(n_5226),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5130),
.Y(n_5493)
);

AOI21xp5_ASAP7_75t_SL g5494 ( 
.A1(n_4969),
.A2(n_1178),
.B(n_1175),
.Y(n_5494)
);

INVx1_ASAP7_75t_SL g5495 ( 
.A(n_4954),
.Y(n_5495)
);

AOI22xp5_ASAP7_75t_L g5496 ( 
.A1(n_5102),
.A2(n_1093),
.B1(n_2313),
.B2(n_2307),
.Y(n_5496)
);

INVx5_ASAP7_75t_L g5497 ( 
.A(n_5226),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_4945),
.Y(n_5498)
);

AOI21xp5_ASAP7_75t_L g5499 ( 
.A1(n_5048),
.A2(n_2902),
.B(n_2901),
.Y(n_5499)
);

AOI211x1_ASAP7_75t_L g5500 ( 
.A1(n_4998),
.A2(n_32),
.B(n_33),
.C(n_42),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5050),
.B(n_1182),
.Y(n_5501)
);

OAI21x1_ASAP7_75t_L g5502 ( 
.A1(n_5020),
.A2(n_3013),
.B(n_3003),
.Y(n_5502)
);

BUFx3_ASAP7_75t_L g5503 ( 
.A(n_5060),
.Y(n_5503)
);

AOI21xp5_ASAP7_75t_L g5504 ( 
.A1(n_5092),
.A2(n_2906),
.B(n_2902),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_5192),
.Y(n_5505)
);

OAI21x1_ASAP7_75t_L g5506 ( 
.A1(n_4967),
.A2(n_3014),
.B(n_3013),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5202),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5053),
.B(n_1183),
.Y(n_5508)
);

AOI211x1_ASAP7_75t_L g5509 ( 
.A1(n_5207),
.A2(n_47),
.B(n_44),
.C(n_45),
.Y(n_5509)
);

A2O1A1Ixp33_ASAP7_75t_L g5510 ( 
.A1(n_5127),
.A2(n_1185),
.B(n_1184),
.C(n_2249),
.Y(n_5510)
);

AOI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_5102),
.A2(n_2307),
.B1(n_2328),
.B2(n_2313),
.Y(n_5511)
);

AO21x1_ASAP7_75t_L g5512 ( 
.A1(n_5217),
.A2(n_44),
.B(n_48),
.Y(n_5512)
);

NAND2x1p5_ASAP7_75t_L g5513 ( 
.A(n_5156),
.B(n_2473),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5194),
.Y(n_5514)
);

INVxp67_ASAP7_75t_L g5515 ( 
.A(n_5066),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_L g5516 ( 
.A(n_5104),
.B(n_5026),
.Y(n_5516)
);

OAI21xp5_ASAP7_75t_L g5517 ( 
.A1(n_5127),
.A2(n_2910),
.B(n_2907),
.Y(n_5517)
);

AO21x2_ASAP7_75t_L g5518 ( 
.A1(n_5082),
.A2(n_3079),
.B(n_3075),
.Y(n_5518)
);

BUFx2_ASAP7_75t_L g5519 ( 
.A(n_5237),
.Y(n_5519)
);

NOR2x1_ASAP7_75t_SL g5520 ( 
.A(n_5117),
.B(n_2915),
.Y(n_5520)
);

OAI21x1_ASAP7_75t_L g5521 ( 
.A1(n_5144),
.A2(n_3018),
.B(n_3014),
.Y(n_5521)
);

AOI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5187),
.A2(n_2917),
.B(n_2541),
.Y(n_5522)
);

NOR4xp25_ASAP7_75t_L g5523 ( 
.A(n_5250),
.B(n_52),
.C(n_49),
.D(n_51),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5026),
.B(n_49),
.Y(n_5524)
);

NAND2x1p5_ASAP7_75t_L g5525 ( 
.A(n_5156),
.B(n_2473),
.Y(n_5525)
);

AND2x2_ASAP7_75t_L g5526 ( 
.A(n_5110),
.B(n_5113),
.Y(n_5526)
);

NOR2xp33_ASAP7_75t_SL g5527 ( 
.A(n_5110),
.B(n_2917),
.Y(n_5527)
);

INVx4_ASAP7_75t_L g5528 ( 
.A(n_4973),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5256),
.B(n_51),
.Y(n_5529)
);

AOI21xp5_ASAP7_75t_L g5530 ( 
.A1(n_5054),
.A2(n_2801),
.B(n_2773),
.Y(n_5530)
);

BUFx6f_ASAP7_75t_L g5531 ( 
.A(n_4973),
.Y(n_5531)
);

HB1xp67_ASAP7_75t_L g5532 ( 
.A(n_4988),
.Y(n_5532)
);

OAI21xp5_ASAP7_75t_L g5533 ( 
.A1(n_5018),
.A2(n_2647),
.B(n_2644),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_4988),
.Y(n_5534)
);

OA21x2_ASAP7_75t_L g5535 ( 
.A1(n_5076),
.A2(n_5159),
.B(n_5077),
.Y(n_5535)
);

CKINVDCx5p33_ASAP7_75t_R g5536 ( 
.A(n_5065),
.Y(n_5536)
);

OAI21x1_ASAP7_75t_L g5537 ( 
.A1(n_5147),
.A2(n_3022),
.B(n_3018),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_4988),
.Y(n_5538)
);

OAI21x1_ASAP7_75t_L g5539 ( 
.A1(n_5119),
.A2(n_3024),
.B(n_3022),
.Y(n_5539)
);

BUFx6f_ASAP7_75t_L g5540 ( 
.A(n_5065),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_L g5541 ( 
.A(n_5268),
.B(n_52),
.Y(n_5541)
);

OAI21xp5_ASAP7_75t_L g5542 ( 
.A1(n_4952),
.A2(n_2647),
.B(n_2644),
.Y(n_5542)
);

AOI21xp5_ASAP7_75t_L g5543 ( 
.A1(n_5043),
.A2(n_2806),
.B(n_2801),
.Y(n_5543)
);

AND2x4_ASAP7_75t_L g5544 ( 
.A(n_4907),
.B(n_54),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_5250),
.B(n_55),
.Y(n_5545)
);

BUFx6f_ASAP7_75t_L g5546 ( 
.A(n_5079),
.Y(n_5546)
);

AOI21xp33_ASAP7_75t_L g5547 ( 
.A1(n_5152),
.A2(n_55),
.B(n_56),
.Y(n_5547)
);

AOI21xp5_ASAP7_75t_L g5548 ( 
.A1(n_5044),
.A2(n_2806),
.B(n_2801),
.Y(n_5548)
);

OAI21x1_ASAP7_75t_L g5549 ( 
.A1(n_5062),
.A2(n_3027),
.B(n_3024),
.Y(n_5549)
);

NOR3xp33_ASAP7_75t_L g5550 ( 
.A(n_4936),
.B(n_2680),
.C(n_2663),
.Y(n_5550)
);

INVx6_ASAP7_75t_L g5551 ( 
.A(n_5079),
.Y(n_5551)
);

NAND2xp5_ASAP7_75t_L g5552 ( 
.A(n_5217),
.B(n_57),
.Y(n_5552)
);

OAI22xp5_ASAP7_75t_L g5553 ( 
.A1(n_5023),
.A2(n_2655),
.B1(n_2658),
.B2(n_2654),
.Y(n_5553)
);

OAI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5045),
.A2(n_2655),
.B(n_2654),
.Y(n_5554)
);

OAI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_5122),
.A2(n_2662),
.B1(n_2665),
.B2(n_2658),
.Y(n_5555)
);

BUFx6f_ASAP7_75t_L g5556 ( 
.A(n_5079),
.Y(n_5556)
);

AO31x2_ASAP7_75t_L g5557 ( 
.A1(n_5164),
.A2(n_3035),
.A3(n_3036),
.B(n_3033),
.Y(n_5557)
);

OAI21x1_ASAP7_75t_L g5558 ( 
.A1(n_5178),
.A2(n_3036),
.B(n_3035),
.Y(n_5558)
);

AOI21xp5_ASAP7_75t_L g5559 ( 
.A1(n_5142),
.A2(n_2806),
.B(n_2801),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4957),
.Y(n_5560)
);

OAI21x1_ASAP7_75t_L g5561 ( 
.A1(n_5179),
.A2(n_3042),
.B(n_3040),
.Y(n_5561)
);

AOI21xp5_ASAP7_75t_L g5562 ( 
.A1(n_5142),
.A2(n_2817),
.B(n_2806),
.Y(n_5562)
);

INVx2_ASAP7_75t_SL g5563 ( 
.A(n_5088),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_4957),
.Y(n_5564)
);

AND2x2_ASAP7_75t_L g5565 ( 
.A(n_5113),
.B(n_57),
.Y(n_5565)
);

AOI21x1_ASAP7_75t_L g5566 ( 
.A1(n_5170),
.A2(n_2665),
.B(n_2662),
.Y(n_5566)
);

AOI21xp5_ASAP7_75t_L g5567 ( 
.A1(n_5163),
.A2(n_2817),
.B(n_2806),
.Y(n_5567)
);

OAI21xp5_ASAP7_75t_L g5568 ( 
.A1(n_5263),
.A2(n_2668),
.B(n_2667),
.Y(n_5568)
);

NOR2xp33_ASAP7_75t_L g5569 ( 
.A(n_5220),
.B(n_5227),
.Y(n_5569)
);

AO31x2_ASAP7_75t_L g5570 ( 
.A1(n_5103),
.A2(n_3042),
.A3(n_3048),
.B(n_3040),
.Y(n_5570)
);

OAI21x1_ASAP7_75t_L g5571 ( 
.A1(n_5186),
.A2(n_3054),
.B(n_3048),
.Y(n_5571)
);

AND2x4_ASAP7_75t_L g5572 ( 
.A(n_5117),
.B(n_58),
.Y(n_5572)
);

OA21x2_ASAP7_75t_L g5573 ( 
.A1(n_4928),
.A2(n_2661),
.B(n_2660),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_4957),
.Y(n_5574)
);

BUFx2_ASAP7_75t_L g5575 ( 
.A(n_5237),
.Y(n_5575)
);

AOI21xp5_ASAP7_75t_L g5576 ( 
.A1(n_5163),
.A2(n_2817),
.B(n_2806),
.Y(n_5576)
);

OR2x2_ASAP7_75t_L g5577 ( 
.A(n_5176),
.B(n_59),
.Y(n_5577)
);

OAI21x1_ASAP7_75t_L g5578 ( 
.A1(n_5205),
.A2(n_3071),
.B(n_3054),
.Y(n_5578)
);

O2A1O1Ixp33_ASAP7_75t_L g5579 ( 
.A1(n_5135),
.A2(n_2249),
.B(n_62),
.C(n_60),
.Y(n_5579)
);

A2O1A1Ixp33_ASAP7_75t_L g5580 ( 
.A1(n_5267),
.A2(n_2313),
.B(n_2328),
.C(n_2307),
.Y(n_5580)
);

OAI21x1_ASAP7_75t_L g5581 ( 
.A1(n_5209),
.A2(n_3074),
.B(n_3071),
.Y(n_5581)
);

AOI21xp5_ASAP7_75t_L g5582 ( 
.A1(n_5236),
.A2(n_2819),
.B(n_2817),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5227),
.B(n_60),
.Y(n_5583)
);

AND2x2_ASAP7_75t_L g5584 ( 
.A(n_5128),
.B(n_61),
.Y(n_5584)
);

AND3x4_ASAP7_75t_L g5585 ( 
.A(n_5166),
.B(n_63),
.C(n_64),
.Y(n_5585)
);

OAI21x1_ASAP7_75t_L g5586 ( 
.A1(n_5235),
.A2(n_3075),
.B(n_3074),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_4920),
.Y(n_5587)
);

OAI21x1_ASAP7_75t_L g5588 ( 
.A1(n_5356),
.A2(n_5203),
.B(n_5199),
.Y(n_5588)
);

AO21x2_ASAP7_75t_L g5589 ( 
.A1(n_5291),
.A2(n_5236),
.B(n_4942),
.Y(n_5589)
);

OAI21x1_ASAP7_75t_L g5590 ( 
.A1(n_5270),
.A2(n_4929),
.B(n_5243),
.Y(n_5590)
);

OAI21x1_ASAP7_75t_L g5591 ( 
.A1(n_5271),
.A2(n_4929),
.B(n_5243),
.Y(n_5591)
);

INVx2_ASAP7_75t_L g5592 ( 
.A(n_5374),
.Y(n_5592)
);

NAND3xp33_ASAP7_75t_L g5593 ( 
.A(n_5299),
.B(n_5019),
.C(n_4994),
.Y(n_5593)
);

OAI21x1_ASAP7_75t_L g5594 ( 
.A1(n_5355),
.A2(n_5259),
.B(n_4938),
.Y(n_5594)
);

AOI22x1_ASAP7_75t_L g5595 ( 
.A1(n_5327),
.A2(n_5128),
.B1(n_5173),
.B2(n_5259),
.Y(n_5595)
);

NOR2xp33_ASAP7_75t_L g5596 ( 
.A(n_5322),
.B(n_5240),
.Y(n_5596)
);

OAI21x1_ASAP7_75t_L g5597 ( 
.A1(n_5435),
.A2(n_4986),
.B(n_5266),
.Y(n_5597)
);

AOI22xp33_ASAP7_75t_L g5598 ( 
.A1(n_5416),
.A2(n_4989),
.B1(n_5105),
.B2(n_5094),
.Y(n_5598)
);

OAI21x1_ASAP7_75t_L g5599 ( 
.A1(n_5315),
.A2(n_5266),
.B(n_4983),
.Y(n_5599)
);

INVx4_ASAP7_75t_L g5600 ( 
.A(n_5309),
.Y(n_5600)
);

INVx2_ASAP7_75t_L g5601 ( 
.A(n_5374),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_5318),
.Y(n_5602)
);

BUFx2_ASAP7_75t_L g5603 ( 
.A(n_5338),
.Y(n_5603)
);

HB1xp67_ASAP7_75t_L g5604 ( 
.A(n_5308),
.Y(n_5604)
);

OA21x2_ASAP7_75t_L g5605 ( 
.A1(n_5587),
.A2(n_4942),
.B(n_5234),
.Y(n_5605)
);

HB1xp67_ASAP7_75t_L g5606 ( 
.A(n_5308),
.Y(n_5606)
);

NOR2xp33_ASAP7_75t_L g5607 ( 
.A(n_5288),
.B(n_5210),
.Y(n_5607)
);

AOI22xp5_ASAP7_75t_L g5608 ( 
.A1(n_5585),
.A2(n_5003),
.B1(n_5072),
.B2(n_5005),
.Y(n_5608)
);

BUFx3_ASAP7_75t_L g5609 ( 
.A(n_5275),
.Y(n_5609)
);

AND2x2_ASAP7_75t_L g5610 ( 
.A(n_5420),
.B(n_4999),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_5279),
.Y(n_5611)
);

NOR2xp33_ASAP7_75t_L g5612 ( 
.A(n_5334),
.B(n_5211),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5340),
.Y(n_5613)
);

OA21x2_ASAP7_75t_L g5614 ( 
.A1(n_5587),
.A2(n_5019),
.B(n_5177),
.Y(n_5614)
);

INVx2_ASAP7_75t_L g5615 ( 
.A(n_5316),
.Y(n_5615)
);

OAI21x1_ASAP7_75t_L g5616 ( 
.A1(n_5283),
.A2(n_5172),
.B(n_5097),
.Y(n_5616)
);

BUFx2_ASAP7_75t_L g5617 ( 
.A(n_5305),
.Y(n_5617)
);

INVx2_ASAP7_75t_SL g5618 ( 
.A(n_5305),
.Y(n_5618)
);

NOR2xp33_ASAP7_75t_L g5619 ( 
.A(n_5306),
.B(n_5058),
.Y(n_5619)
);

BUFx2_ASAP7_75t_R g5620 ( 
.A(n_5488),
.Y(n_5620)
);

NAND2x1p5_ASAP7_75t_L g5621 ( 
.A(n_5492),
.B(n_5117),
.Y(n_5621)
);

AOI21xp5_ASAP7_75t_L g5622 ( 
.A1(n_5443),
.A2(n_5003),
.B(n_5134),
.Y(n_5622)
);

OR2x6_ASAP7_75t_L g5623 ( 
.A(n_5284),
.B(n_5055),
.Y(n_5623)
);

OAI21xp5_ASAP7_75t_L g5624 ( 
.A1(n_5363),
.A2(n_5105),
.B(n_5094),
.Y(n_5624)
);

OAI21x1_ASAP7_75t_L g5625 ( 
.A1(n_5452),
.A2(n_5047),
.B(n_5197),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5388),
.B(n_5171),
.Y(n_5626)
);

CKINVDCx11_ASAP7_75t_R g5627 ( 
.A(n_5337),
.Y(n_5627)
);

OAI21xp5_ASAP7_75t_L g5628 ( 
.A1(n_5523),
.A2(n_4989),
.B(n_5025),
.Y(n_5628)
);

BUFx3_ASAP7_75t_L g5629 ( 
.A(n_5275),
.Y(n_5629)
);

BUFx3_ASAP7_75t_L g5630 ( 
.A(n_5459),
.Y(n_5630)
);

OAI21xp5_ASAP7_75t_L g5631 ( 
.A1(n_5352),
.A2(n_5399),
.B(n_5299),
.Y(n_5631)
);

INVx4_ASAP7_75t_L g5632 ( 
.A(n_5371),
.Y(n_5632)
);

OAI21x1_ASAP7_75t_L g5633 ( 
.A1(n_5452),
.A2(n_5188),
.B(n_5228),
.Y(n_5633)
);

AO21x2_ASAP7_75t_L g5634 ( 
.A1(n_5414),
.A2(n_4968),
.B(n_5068),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5345),
.Y(n_5635)
);

AO21x2_ASAP7_75t_L g5636 ( 
.A1(n_5469),
.A2(n_5116),
.B(n_5121),
.Y(n_5636)
);

INVx3_ASAP7_75t_L g5637 ( 
.A(n_5310),
.Y(n_5637)
);

NOR2xp33_ASAP7_75t_L g5638 ( 
.A(n_5272),
.B(n_5569),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5345),
.Y(n_5639)
);

BUFx4f_ASAP7_75t_L g5640 ( 
.A(n_5572),
.Y(n_5640)
);

AO21x2_ASAP7_75t_L g5641 ( 
.A1(n_5469),
.A2(n_5153),
.B(n_5141),
.Y(n_5641)
);

NAND3xp33_ASAP7_75t_L g5642 ( 
.A(n_5384),
.B(n_5145),
.C(n_5219),
.Y(n_5642)
);

INVxp67_ASAP7_75t_L g5643 ( 
.A(n_5457),
.Y(n_5643)
);

AOI21xp5_ASAP7_75t_L g5644 ( 
.A1(n_5543),
.A2(n_5246),
.B(n_5215),
.Y(n_5644)
);

AO21x2_ASAP7_75t_L g5645 ( 
.A1(n_5498),
.A2(n_5141),
.B(n_4980),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5303),
.Y(n_5646)
);

OR2x6_ASAP7_75t_L g5647 ( 
.A(n_5276),
.B(n_5055),
.Y(n_5647)
);

INVx3_ASAP7_75t_L g5648 ( 
.A(n_5310),
.Y(n_5648)
);

NAND3xp33_ASAP7_75t_L g5649 ( 
.A(n_5321),
.B(n_5219),
.C(n_5162),
.Y(n_5649)
);

NAND2x1p5_ASAP7_75t_L g5650 ( 
.A(n_5492),
.B(n_5088),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_5493),
.Y(n_5651)
);

INVx2_ASAP7_75t_SL g5652 ( 
.A(n_5357),
.Y(n_5652)
);

NOR2xp67_ASAP7_75t_SL g5653 ( 
.A(n_5357),
.B(n_5183),
.Y(n_5653)
);

AO21x2_ASAP7_75t_L g5654 ( 
.A1(n_5534),
.A2(n_4987),
.B(n_4975),
.Y(n_5654)
);

OA21x2_ASAP7_75t_L g5655 ( 
.A1(n_5538),
.A2(n_5061),
.B(n_5085),
.Y(n_5655)
);

OAI21x1_ASAP7_75t_L g5656 ( 
.A1(n_5361),
.A2(n_5228),
.B(n_4991),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_5505),
.Y(n_5657)
);

OA21x2_ASAP7_75t_L g5658 ( 
.A1(n_5560),
.A2(n_5040),
.B(n_5200),
.Y(n_5658)
);

AO21x2_ASAP7_75t_L g5659 ( 
.A1(n_5564),
.A2(n_5574),
.B(n_5532),
.Y(n_5659)
);

CKINVDCx16_ASAP7_75t_R g5660 ( 
.A(n_5400),
.Y(n_5660)
);

OAI21x1_ASAP7_75t_L g5661 ( 
.A1(n_5373),
.A2(n_5190),
.B(n_5149),
.Y(n_5661)
);

OAI21x1_ASAP7_75t_L g5662 ( 
.A1(n_5269),
.A2(n_5257),
.B(n_5247),
.Y(n_5662)
);

OAI21x1_ASAP7_75t_L g5663 ( 
.A1(n_5269),
.A2(n_5260),
.B(n_5230),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5314),
.Y(n_5664)
);

AOI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_5274),
.A2(n_5075),
.B1(n_5218),
.B2(n_5167),
.Y(n_5665)
);

OAI22xp33_ASAP7_75t_L g5666 ( 
.A1(n_5282),
.A2(n_5167),
.B1(n_5108),
.B2(n_5262),
.Y(n_5666)
);

OAI21x1_ASAP7_75t_L g5667 ( 
.A1(n_5382),
.A2(n_5230),
.B(n_5138),
.Y(n_5667)
);

HB1xp67_ASAP7_75t_L g5668 ( 
.A(n_5289),
.Y(n_5668)
);

AO21x2_ASAP7_75t_L g5669 ( 
.A1(n_5377),
.A2(n_5198),
.B(n_5115),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_5512),
.A2(n_5262),
.B1(n_5108),
.B2(n_5115),
.Y(n_5670)
);

AOI21x1_ASAP7_75t_L g5671 ( 
.A1(n_5358),
.A2(n_5304),
.B(n_5344),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_5415),
.Y(n_5672)
);

NAND2xp5_ASAP7_75t_L g5673 ( 
.A(n_5292),
.B(n_4920),
.Y(n_5673)
);

OAI21x1_ASAP7_75t_L g5674 ( 
.A1(n_5319),
.A2(n_5037),
.B(n_5030),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5317),
.Y(n_5675)
);

OAI21x1_ASAP7_75t_SL g5676 ( 
.A1(n_5394),
.A2(n_5462),
.B(n_5433),
.Y(n_5676)
);

AOI21xp33_ASAP7_75t_L g5677 ( 
.A1(n_5468),
.A2(n_5100),
.B(n_5191),
.Y(n_5677)
);

OAI21x1_ASAP7_75t_SL g5678 ( 
.A1(n_5394),
.A2(n_5133),
.B(n_5265),
.Y(n_5678)
);

AOI21xp5_ASAP7_75t_L g5679 ( 
.A1(n_5548),
.A2(n_5093),
.B(n_5242),
.Y(n_5679)
);

OAI21xp5_ASAP7_75t_L g5680 ( 
.A1(n_5406),
.A2(n_5093),
.B(n_5195),
.Y(n_5680)
);

AOI21xp33_ASAP7_75t_L g5681 ( 
.A1(n_5468),
.A2(n_5133),
.B(n_5120),
.Y(n_5681)
);

OR2x6_ASAP7_75t_L g5682 ( 
.A(n_5572),
.B(n_5204),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5335),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5336),
.Y(n_5684)
);

OAI21x1_ASAP7_75t_L g5685 ( 
.A1(n_5490),
.A2(n_5261),
.B(n_5231),
.Y(n_5685)
);

AND2x4_ASAP7_75t_L g5686 ( 
.A(n_5286),
.B(n_4920),
.Y(n_5686)
);

BUFx6f_ASAP7_75t_L g5687 ( 
.A(n_5364),
.Y(n_5687)
);

OAI21x1_ASAP7_75t_L g5688 ( 
.A1(n_5530),
.A2(n_5225),
.B(n_5180),
.Y(n_5688)
);

AND2x4_ASAP7_75t_L g5689 ( 
.A(n_5280),
.B(n_5168),
.Y(n_5689)
);

OAI21x1_ASAP7_75t_L g5690 ( 
.A1(n_5293),
.A2(n_5241),
.B(n_5114),
.Y(n_5690)
);

AND2x2_ASAP7_75t_L g5691 ( 
.A(n_5341),
.B(n_5204),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5424),
.Y(n_5692)
);

BUFx3_ASAP7_75t_L g5693 ( 
.A(n_5364),
.Y(n_5693)
);

INVx8_ASAP7_75t_L g5694 ( 
.A(n_5371),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5441),
.Y(n_5695)
);

AO21x2_ASAP7_75t_L g5696 ( 
.A1(n_5529),
.A2(n_5198),
.B(n_5233),
.Y(n_5696)
);

OA21x2_ASAP7_75t_L g5697 ( 
.A1(n_5402),
.A2(n_5143),
.B(n_5233),
.Y(n_5697)
);

OAI21x1_ASAP7_75t_L g5698 ( 
.A1(n_5380),
.A2(n_5091),
.B(n_5168),
.Y(n_5698)
);

AO21x2_ASAP7_75t_L g5699 ( 
.A1(n_5541),
.A2(n_5143),
.B(n_5091),
.Y(n_5699)
);

OAI21x1_ASAP7_75t_L g5700 ( 
.A1(n_5339),
.A2(n_5091),
.B(n_5168),
.Y(n_5700)
);

OAI21x1_ASAP7_75t_L g5701 ( 
.A1(n_5339),
.A2(n_5080),
.B(n_5155),
.Y(n_5701)
);

AOI22xp33_ASAP7_75t_L g5702 ( 
.A1(n_5484),
.A2(n_2313),
.B1(n_2328),
.B2(n_2307),
.Y(n_5702)
);

AOI22xp33_ASAP7_75t_L g5703 ( 
.A1(n_5484),
.A2(n_2328),
.B1(n_2329),
.B2(n_2313),
.Y(n_5703)
);

NAND3xp33_ASAP7_75t_L g5704 ( 
.A(n_5439),
.B(n_2329),
.C(n_2328),
.Y(n_5704)
);

INVx8_ASAP7_75t_L g5705 ( 
.A(n_5544),
.Y(n_5705)
);

AO21x1_ASAP7_75t_L g5706 ( 
.A1(n_5407),
.A2(n_5080),
.B(n_63),
.Y(n_5706)
);

OAI21x1_ASAP7_75t_L g5707 ( 
.A1(n_5367),
.A2(n_5080),
.B(n_5155),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5470),
.Y(n_5708)
);

INVx2_ASAP7_75t_L g5709 ( 
.A(n_5471),
.Y(n_5709)
);

AND2x4_ASAP7_75t_L g5710 ( 
.A(n_5280),
.B(n_5155),
.Y(n_5710)
);

BUFx2_ASAP7_75t_L g5711 ( 
.A(n_5458),
.Y(n_5711)
);

BUFx12f_ASAP7_75t_L g5712 ( 
.A(n_5332),
.Y(n_5712)
);

NAND2xp5_ASAP7_75t_L g5713 ( 
.A(n_5402),
.B(n_5216),
.Y(n_5713)
);

NAND2x1p5_ASAP7_75t_L g5714 ( 
.A(n_5492),
.B(n_2473),
.Y(n_5714)
);

OAI21x1_ASAP7_75t_L g5715 ( 
.A1(n_5300),
.A2(n_5239),
.B(n_5216),
.Y(n_5715)
);

OAI21x1_ASAP7_75t_L g5716 ( 
.A1(n_5418),
.A2(n_5239),
.B(n_2569),
.Y(n_5716)
);

INVx5_ASAP7_75t_L g5717 ( 
.A(n_5332),
.Y(n_5717)
);

HB1xp67_ASAP7_75t_L g5718 ( 
.A(n_5278),
.Y(n_5718)
);

NAND3xp33_ASAP7_75t_L g5719 ( 
.A(n_5390),
.B(n_2329),
.C(n_1362),
.Y(n_5719)
);

OAI21x1_ASAP7_75t_L g5720 ( 
.A1(n_5516),
.A2(n_2569),
.B(n_2540),
.Y(n_5720)
);

CKINVDCx20_ASAP7_75t_R g5721 ( 
.A(n_5328),
.Y(n_5721)
);

INVx5_ASAP7_75t_L g5722 ( 
.A(n_5332),
.Y(n_5722)
);

INVx1_ASAP7_75t_SL g5723 ( 
.A(n_5495),
.Y(n_5723)
);

BUFx3_ASAP7_75t_L g5724 ( 
.A(n_5391),
.Y(n_5724)
);

AOI221xp5_ASAP7_75t_L g5725 ( 
.A1(n_5365),
.A2(n_1447),
.B1(n_1470),
.B2(n_1362),
.C(n_1267),
.Y(n_5725)
);

OAI21x1_ASAP7_75t_L g5726 ( 
.A1(n_5386),
.A2(n_2569),
.B(n_2540),
.Y(n_5726)
);

INVx2_ASAP7_75t_L g5727 ( 
.A(n_5489),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5507),
.Y(n_5728)
);

AO21x2_ASAP7_75t_L g5729 ( 
.A1(n_5348),
.A2(n_3083),
.B(n_3079),
.Y(n_5729)
);

OAI21x1_ASAP7_75t_L g5730 ( 
.A1(n_5566),
.A2(n_2569),
.B(n_2540),
.Y(n_5730)
);

OAI21x1_ASAP7_75t_L g5731 ( 
.A1(n_5375),
.A2(n_5582),
.B(n_5410),
.Y(n_5731)
);

OAI21x1_ASAP7_75t_L g5732 ( 
.A1(n_5351),
.A2(n_2589),
.B(n_2575),
.Y(n_5732)
);

AOI21xp5_ASAP7_75t_L g5733 ( 
.A1(n_5559),
.A2(n_2486),
.B(n_2473),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5450),
.Y(n_5734)
);

OR2x6_ASAP7_75t_L g5735 ( 
.A(n_5395),
.B(n_3083),
.Y(n_5735)
);

OAI21x1_ASAP7_75t_SL g5736 ( 
.A1(n_5462),
.A2(n_5520),
.B(n_5294),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5514),
.Y(n_5737)
);

BUFx4f_ASAP7_75t_SL g5738 ( 
.A(n_5503),
.Y(n_5738)
);

OAI21x1_ASAP7_75t_L g5739 ( 
.A1(n_5526),
.A2(n_2589),
.B(n_2575),
.Y(n_5739)
);

OAI21xp5_ASAP7_75t_L g5740 ( 
.A1(n_5510),
.A2(n_66),
.B(n_67),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5381),
.Y(n_5741)
);

INVx3_ASAP7_75t_L g5742 ( 
.A(n_5528),
.Y(n_5742)
);

OAI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5312),
.A2(n_5567),
.B(n_5562),
.Y(n_5743)
);

CKINVDCx20_ASAP7_75t_R g5744 ( 
.A(n_5536),
.Y(n_5744)
);

OAI21x1_ASAP7_75t_L g5745 ( 
.A1(n_5576),
.A2(n_2589),
.B(n_2575),
.Y(n_5745)
);

O2A1O1Ixp33_ASAP7_75t_L g5746 ( 
.A1(n_5431),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_5746)
);

OAI21x1_ASAP7_75t_L g5747 ( 
.A1(n_5444),
.A2(n_2589),
.B(n_2575),
.Y(n_5747)
);

BUFx2_ASAP7_75t_R g5748 ( 
.A(n_5302),
.Y(n_5748)
);

INVxp67_ASAP7_75t_L g5749 ( 
.A(n_5519),
.Y(n_5749)
);

NAND2xp5_ASAP7_75t_L g5750 ( 
.A(n_5575),
.B(n_69),
.Y(n_5750)
);

OAI21x1_ASAP7_75t_L g5751 ( 
.A1(n_5296),
.A2(n_2601),
.B(n_2595),
.Y(n_5751)
);

OAI21x1_ASAP7_75t_L g5752 ( 
.A1(n_5368),
.A2(n_2601),
.B(n_2595),
.Y(n_5752)
);

INVx4_ASAP7_75t_L g5753 ( 
.A(n_5544),
.Y(n_5753)
);

OAI21x1_ASAP7_75t_L g5754 ( 
.A1(n_5436),
.A2(n_2601),
.B(n_2595),
.Y(n_5754)
);

AOI21xp5_ASAP7_75t_L g5755 ( 
.A1(n_5438),
.A2(n_5520),
.B(n_5342),
.Y(n_5755)
);

NOR2xp33_ASAP7_75t_L g5756 ( 
.A(n_5545),
.B(n_70),
.Y(n_5756)
);

AND2x4_ASAP7_75t_L g5757 ( 
.A(n_5515),
.B(n_71),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_5326),
.Y(n_5758)
);

AO21x2_ASAP7_75t_L g5759 ( 
.A1(n_5323),
.A2(n_3088),
.B(n_3087),
.Y(n_5759)
);

BUFx6f_ASAP7_75t_L g5760 ( 
.A(n_5531),
.Y(n_5760)
);

OAI21x1_ASAP7_75t_L g5761 ( 
.A1(n_5448),
.A2(n_2601),
.B(n_2595),
.Y(n_5761)
);

AOI21xp5_ASAP7_75t_L g5762 ( 
.A1(n_5329),
.A2(n_2486),
.B(n_2473),
.Y(n_5762)
);

AO21x2_ASAP7_75t_L g5763 ( 
.A1(n_5297),
.A2(n_2602),
.B(n_2599),
.Y(n_5763)
);

OAI21x1_ASAP7_75t_L g5764 ( 
.A1(n_5447),
.A2(n_2639),
.B(n_2610),
.Y(n_5764)
);

OAI21x1_ASAP7_75t_L g5765 ( 
.A1(n_5454),
.A2(n_2639),
.B(n_2610),
.Y(n_5765)
);

OAI21x1_ASAP7_75t_L g5766 ( 
.A1(n_5524),
.A2(n_2639),
.B(n_2610),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5311),
.Y(n_5767)
);

INVx8_ASAP7_75t_L g5768 ( 
.A(n_5324),
.Y(n_5768)
);

INVxp67_ASAP7_75t_L g5769 ( 
.A(n_5320),
.Y(n_5769)
);

BUFx12f_ASAP7_75t_L g5770 ( 
.A(n_5287),
.Y(n_5770)
);

AOI21x1_ASAP7_75t_L g5771 ( 
.A1(n_5301),
.A2(n_2681),
.B(n_2674),
.Y(n_5771)
);

INVx2_ASAP7_75t_SL g5772 ( 
.A(n_5333),
.Y(n_5772)
);

NAND2x1p5_ASAP7_75t_L g5773 ( 
.A(n_5497),
.B(n_2473),
.Y(n_5773)
);

AOI21x1_ASAP7_75t_L g5774 ( 
.A1(n_5401),
.A2(n_2681),
.B(n_2674),
.Y(n_5774)
);

OR2x2_ASAP7_75t_L g5775 ( 
.A(n_5479),
.B(n_5397),
.Y(n_5775)
);

INVx4_ASAP7_75t_L g5776 ( 
.A(n_5324),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5311),
.Y(n_5777)
);

NAND2x1p5_ASAP7_75t_L g5778 ( 
.A(n_5497),
.B(n_2486),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5311),
.Y(n_5779)
);

INVx8_ASAP7_75t_L g5780 ( 
.A(n_5440),
.Y(n_5780)
);

BUFx8_ASAP7_75t_SL g5781 ( 
.A(n_5307),
.Y(n_5781)
);

OAI21x1_ASAP7_75t_L g5782 ( 
.A1(n_5477),
.A2(n_2639),
.B(n_2610),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5396),
.Y(n_5783)
);

OAI21x1_ASAP7_75t_L g5784 ( 
.A1(n_5330),
.A2(n_2721),
.B(n_2711),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5535),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5535),
.Y(n_5786)
);

OA21x2_ASAP7_75t_L g5787 ( 
.A1(n_5474),
.A2(n_2664),
.B(n_2742),
.Y(n_5787)
);

AOI22x1_ASAP7_75t_L g5788 ( 
.A1(n_5565),
.A2(n_2756),
.B1(n_2757),
.B2(n_2683),
.Y(n_5788)
);

BUFx8_ASAP7_75t_L g5789 ( 
.A(n_5584),
.Y(n_5789)
);

NOR2xp33_ASAP7_75t_L g5790 ( 
.A(n_5552),
.B(n_71),
.Y(n_5790)
);

OAI21x1_ASAP7_75t_L g5791 ( 
.A1(n_5558),
.A2(n_2731),
.B(n_2723),
.Y(n_5791)
);

NAND3xp33_ASAP7_75t_L g5792 ( 
.A(n_5509),
.B(n_2329),
.C(n_1447),
.Y(n_5792)
);

INVx2_ASAP7_75t_L g5793 ( 
.A(n_5325),
.Y(n_5793)
);

NAND3xp33_ASAP7_75t_L g5794 ( 
.A(n_5378),
.B(n_2329),
.C(n_1470),
.Y(n_5794)
);

INVx1_ASAP7_75t_SL g5795 ( 
.A(n_5467),
.Y(n_5795)
);

INVx1_ASAP7_75t_SL g5796 ( 
.A(n_5440),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5325),
.Y(n_5797)
);

NAND2xp5_ASAP7_75t_L g5798 ( 
.A(n_5281),
.B(n_72),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5417),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5325),
.Y(n_5800)
);

AO21x2_ASAP7_75t_L g5801 ( 
.A1(n_5485),
.A2(n_5508),
.B(n_5501),
.Y(n_5801)
);

OAI21x1_ASAP7_75t_L g5802 ( 
.A1(n_5561),
.A2(n_2738),
.B(n_2723),
.Y(n_5802)
);

OAI21x1_ASAP7_75t_L g5803 ( 
.A1(n_5571),
.A2(n_2740),
.B(n_2738),
.Y(n_5803)
);

AOI22xp5_ASAP7_75t_L g5804 ( 
.A1(n_5376),
.A2(n_2496),
.B1(n_2497),
.B2(n_2486),
.Y(n_5804)
);

OAI21x1_ASAP7_75t_L g5805 ( 
.A1(n_5578),
.A2(n_2740),
.B(n_2743),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_5583),
.B(n_73),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5417),
.Y(n_5807)
);

OAI21x1_ASAP7_75t_L g5808 ( 
.A1(n_5581),
.A2(n_2748),
.B(n_2743),
.Y(n_5808)
);

CKINVDCx20_ASAP7_75t_R g5809 ( 
.A(n_5453),
.Y(n_5809)
);

INVx5_ASAP7_75t_L g5810 ( 
.A(n_5387),
.Y(n_5810)
);

INVxp67_ASAP7_75t_SL g5811 ( 
.A(n_5577),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5349),
.A2(n_2604),
.B(n_2663),
.Y(n_5812)
);

AO21x2_ASAP7_75t_L g5813 ( 
.A1(n_5369),
.A2(n_2756),
.B(n_2683),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5417),
.Y(n_5814)
);

OAI21x1_ASAP7_75t_L g5815 ( 
.A1(n_5313),
.A2(n_2682),
.B(n_2680),
.Y(n_5815)
);

BUFx2_ASAP7_75t_L g5816 ( 
.A(n_5528),
.Y(n_5816)
);

BUFx10_ASAP7_75t_L g5817 ( 
.A(n_5353),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5518),
.Y(n_5818)
);

HB1xp67_ASAP7_75t_L g5819 ( 
.A(n_5563),
.Y(n_5819)
);

OAI21x1_ASAP7_75t_L g5820 ( 
.A1(n_5412),
.A2(n_2682),
.B(n_2680),
.Y(n_5820)
);

HB1xp67_ASAP7_75t_L g5821 ( 
.A(n_5387),
.Y(n_5821)
);

OAI21x1_ASAP7_75t_SL g5822 ( 
.A1(n_5463),
.A2(n_74),
.B(n_75),
.Y(n_5822)
);

AO21x2_ASAP7_75t_L g5823 ( 
.A1(n_5511),
.A2(n_2759),
.B(n_2758),
.Y(n_5823)
);

OAI21x1_ASAP7_75t_L g5824 ( 
.A1(n_5419),
.A2(n_2682),
.B(n_2680),
.Y(n_5824)
);

NOR2xp33_ASAP7_75t_L g5825 ( 
.A(n_5475),
.B(n_75),
.Y(n_5825)
);

OAI21x1_ASAP7_75t_SL g5826 ( 
.A1(n_5476),
.A2(n_76),
.B(n_77),
.Y(n_5826)
);

OAI21x1_ASAP7_75t_L g5827 ( 
.A1(n_5426),
.A2(n_2692),
.B(n_2682),
.Y(n_5827)
);

NAND2x1p5_ASAP7_75t_L g5828 ( 
.A(n_5343),
.B(n_2486),
.Y(n_5828)
);

CKINVDCx5p33_ASAP7_75t_R g5829 ( 
.A(n_5392),
.Y(n_5829)
);

OA21x2_ASAP7_75t_L g5830 ( 
.A1(n_5429),
.A2(n_2760),
.B(n_2759),
.Y(n_5830)
);

INVx3_ASAP7_75t_L g5831 ( 
.A(n_5551),
.Y(n_5831)
);

CKINVDCx5p33_ASAP7_75t_R g5832 ( 
.A(n_5551),
.Y(n_5832)
);

AO21x2_ASAP7_75t_L g5833 ( 
.A1(n_5580),
.A2(n_2760),
.B(n_2702),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5570),
.Y(n_5834)
);

BUFx8_ASAP7_75t_L g5835 ( 
.A(n_5531),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5570),
.Y(n_5836)
);

OAI21x1_ASAP7_75t_L g5837 ( 
.A1(n_5432),
.A2(n_2722),
.B(n_2692),
.Y(n_5837)
);

OAI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_5442),
.A2(n_76),
.B(n_78),
.Y(n_5838)
);

BUFx3_ASAP7_75t_L g5839 ( 
.A(n_5531),
.Y(n_5839)
);

OAI21x1_ASAP7_75t_SL g5840 ( 
.A1(n_5579),
.A2(n_80),
.B(n_81),
.Y(n_5840)
);

OAI21x1_ASAP7_75t_L g5841 ( 
.A1(n_5478),
.A2(n_2722),
.B(n_2692),
.Y(n_5841)
);

OAI21x1_ASAP7_75t_L g5842 ( 
.A1(n_5483),
.A2(n_2722),
.B(n_2692),
.Y(n_5842)
);

CKINVDCx20_ASAP7_75t_R g5843 ( 
.A(n_5273),
.Y(n_5843)
);

AOI22xp5_ASAP7_75t_L g5844 ( 
.A1(n_5843),
.A2(n_5437),
.B1(n_5290),
.B2(n_5451),
.Y(n_5844)
);

OAI21xp5_ASAP7_75t_L g5845 ( 
.A1(n_5631),
.A2(n_5385),
.B(n_5480),
.Y(n_5845)
);

BUFx3_ASAP7_75t_L g5846 ( 
.A(n_5627),
.Y(n_5846)
);

OA21x2_ASAP7_75t_L g5847 ( 
.A1(n_5592),
.A2(n_5370),
.B(n_5430),
.Y(n_5847)
);

OAI21xp5_ASAP7_75t_L g5848 ( 
.A1(n_5631),
.A2(n_5496),
.B(n_5434),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5668),
.Y(n_5849)
);

OA21x2_ASAP7_75t_L g5850 ( 
.A1(n_5601),
.A2(n_5446),
.B(n_5408),
.Y(n_5850)
);

OAI21x1_ASAP7_75t_L g5851 ( 
.A1(n_5673),
.A2(n_5573),
.B(n_5506),
.Y(n_5851)
);

INVx2_ASAP7_75t_L g5852 ( 
.A(n_5697),
.Y(n_5852)
);

BUFx3_ASAP7_75t_L g5853 ( 
.A(n_5627),
.Y(n_5853)
);

OR2x6_ASAP7_75t_L g5854 ( 
.A(n_5694),
.B(n_5350),
.Y(n_5854)
);

OA21x2_ASAP7_75t_L g5855 ( 
.A1(n_5785),
.A2(n_5413),
.B(n_5404),
.Y(n_5855)
);

INVx2_ASAP7_75t_L g5856 ( 
.A(n_5697),
.Y(n_5856)
);

AOI21xp5_ASAP7_75t_L g5857 ( 
.A1(n_5666),
.A2(n_5403),
.B(n_5547),
.Y(n_5857)
);

NAND2x1p5_ASAP7_75t_L g5858 ( 
.A(n_5653),
.B(n_5540),
.Y(n_5858)
);

OR2x2_ASAP7_75t_L g5859 ( 
.A(n_5718),
.B(n_5465),
.Y(n_5859)
);

OAI21x1_ASAP7_75t_L g5860 ( 
.A1(n_5743),
.A2(n_5502),
.B(n_5491),
.Y(n_5860)
);

OAI21x1_ASAP7_75t_L g5861 ( 
.A1(n_5590),
.A2(n_5445),
.B(n_5466),
.Y(n_5861)
);

INVx5_ASAP7_75t_L g5862 ( 
.A(n_5600),
.Y(n_5862)
);

A2O1A1Ixp33_ASAP7_75t_L g5863 ( 
.A1(n_5619),
.A2(n_5362),
.B(n_5428),
.C(n_5346),
.Y(n_5863)
);

OA21x2_ASAP7_75t_L g5864 ( 
.A1(n_5786),
.A2(n_5586),
.B(n_5398),
.Y(n_5864)
);

BUFx6f_ASAP7_75t_L g5865 ( 
.A(n_5630),
.Y(n_5865)
);

AO21x2_ASAP7_75t_L g5866 ( 
.A1(n_5659),
.A2(n_5383),
.B(n_5372),
.Y(n_5866)
);

AO31x2_ASAP7_75t_L g5867 ( 
.A1(n_5706),
.A2(n_5285),
.A3(n_5487),
.B(n_5379),
.Y(n_5867)
);

OAI21x1_ASAP7_75t_L g5868 ( 
.A1(n_5591),
.A2(n_5537),
.B(n_5521),
.Y(n_5868)
);

AOI21xp5_ASAP7_75t_L g5869 ( 
.A1(n_5666),
.A2(n_5277),
.B(n_5533),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5604),
.B(n_5461),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_SL g5871 ( 
.A(n_5603),
.B(n_5461),
.Y(n_5871)
);

HB1xp67_ASAP7_75t_L g5872 ( 
.A(n_5606),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5668),
.Y(n_5873)
);

OAI21x1_ASAP7_75t_L g5874 ( 
.A1(n_5626),
.A2(n_5700),
.B(n_5597),
.Y(n_5874)
);

AOI22x1_ASAP7_75t_L g5875 ( 
.A1(n_5660),
.A2(n_5421),
.B1(n_5423),
.B2(n_5387),
.Y(n_5875)
);

OAI21xp5_ASAP7_75t_L g5876 ( 
.A1(n_5593),
.A2(n_5427),
.B(n_5359),
.Y(n_5876)
);

NAND2xp5_ASAP7_75t_L g5877 ( 
.A(n_5606),
.B(n_5461),
.Y(n_5877)
);

OAI21xp5_ASAP7_75t_L g5878 ( 
.A1(n_5593),
.A2(n_5389),
.B(n_5354),
.Y(n_5878)
);

AO21x2_ASAP7_75t_L g5879 ( 
.A1(n_5659),
.A2(n_5366),
.B(n_5347),
.Y(n_5879)
);

INVx2_ASAP7_75t_SL g5880 ( 
.A(n_5694),
.Y(n_5880)
);

OAI21x1_ASAP7_75t_L g5881 ( 
.A1(n_5626),
.A2(n_5539),
.B(n_5549),
.Y(n_5881)
);

OA21x2_ASAP7_75t_L g5882 ( 
.A1(n_5713),
.A2(n_5411),
.B(n_5409),
.Y(n_5882)
);

CKINVDCx20_ASAP7_75t_R g5883 ( 
.A(n_5744),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5811),
.B(n_5613),
.Y(n_5884)
);

OA21x2_ASAP7_75t_L g5885 ( 
.A1(n_5713),
.A2(n_5405),
.B(n_5456),
.Y(n_5885)
);

AOI22xp33_ASAP7_75t_L g5886 ( 
.A1(n_5704),
.A2(n_5360),
.B1(n_5550),
.B2(n_5553),
.Y(n_5886)
);

OAI21x1_ASAP7_75t_L g5887 ( 
.A1(n_5663),
.A2(n_5472),
.B(n_5486),
.Y(n_5887)
);

BUFx10_ASAP7_75t_L g5888 ( 
.A(n_5825),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5635),
.Y(n_5889)
);

OAI21x1_ASAP7_75t_L g5890 ( 
.A1(n_5701),
.A2(n_5707),
.B(n_5588),
.Y(n_5890)
);

OAI21x1_ASAP7_75t_L g5891 ( 
.A1(n_5637),
.A2(n_5504),
.B(n_5499),
.Y(n_5891)
);

BUFx2_ASAP7_75t_L g5892 ( 
.A(n_5744),
.Y(n_5892)
);

AOI22xp5_ASAP7_75t_L g5893 ( 
.A1(n_5843),
.A2(n_5331),
.B1(n_5555),
.B2(n_5568),
.Y(n_5893)
);

NAND2xp5_ASAP7_75t_L g5894 ( 
.A(n_5811),
.B(n_5500),
.Y(n_5894)
);

AO31x2_ASAP7_75t_L g5895 ( 
.A1(n_5619),
.A2(n_5422),
.A3(n_5482),
.B(n_5481),
.Y(n_5895)
);

NOR2x1_ASAP7_75t_SL g5896 ( 
.A(n_5647),
.B(n_5540),
.Y(n_5896)
);

AOI21xp5_ASAP7_75t_L g5897 ( 
.A1(n_5644),
.A2(n_5527),
.B(n_5517),
.Y(n_5897)
);

NOR2xp67_ASAP7_75t_L g5898 ( 
.A(n_5632),
.B(n_5540),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5639),
.Y(n_5899)
);

AO21x2_ASAP7_75t_L g5900 ( 
.A1(n_5818),
.A2(n_5522),
.B(n_5298),
.Y(n_5900)
);

AOI21x1_ASAP7_75t_L g5901 ( 
.A1(n_5671),
.A2(n_5295),
.B(n_5542),
.Y(n_5901)
);

AO21x2_ASAP7_75t_L g5902 ( 
.A1(n_5798),
.A2(n_5494),
.B(n_5554),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_5737),
.Y(n_5903)
);

OAI21x1_ASAP7_75t_L g5904 ( 
.A1(n_5637),
.A2(n_5525),
.B(n_5513),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5711),
.B(n_5421),
.Y(n_5905)
);

CKINVDCx5p33_ASAP7_75t_R g5906 ( 
.A(n_5748),
.Y(n_5906)
);

AO21x2_ASAP7_75t_L g5907 ( 
.A1(n_5798),
.A2(n_5473),
.B(n_5460),
.Y(n_5907)
);

AO22x2_ASAP7_75t_L g5908 ( 
.A1(n_5795),
.A2(n_5775),
.B1(n_5769),
.B2(n_5796),
.Y(n_5908)
);

BUFx6f_ASAP7_75t_L g5909 ( 
.A(n_5630),
.Y(n_5909)
);

OAI21x1_ASAP7_75t_L g5910 ( 
.A1(n_5648),
.A2(n_5570),
.B(n_5464),
.Y(n_5910)
);

NAND2x1p5_ASAP7_75t_L g5911 ( 
.A(n_5640),
.B(n_5546),
.Y(n_5911)
);

AO21x2_ASAP7_75t_L g5912 ( 
.A1(n_5750),
.A2(n_5801),
.B(n_5624),
.Y(n_5912)
);

OAI21x1_ASAP7_75t_L g5913 ( 
.A1(n_5662),
.A2(n_5464),
.B(n_5455),
.Y(n_5913)
);

OA21x2_ASAP7_75t_L g5914 ( 
.A1(n_5749),
.A2(n_5464),
.B(n_5455),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_L g5915 ( 
.A(n_5672),
.B(n_5393),
.Y(n_5915)
);

INVx2_ASAP7_75t_L g5916 ( 
.A(n_5709),
.Y(n_5916)
);

INVxp67_ASAP7_75t_SL g5917 ( 
.A(n_5769),
.Y(n_5917)
);

INVx3_ASAP7_75t_L g5918 ( 
.A(n_5632),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5727),
.Y(n_5919)
);

AOI21xp5_ASAP7_75t_L g5920 ( 
.A1(n_5644),
.A2(n_5425),
.B(n_5546),
.Y(n_5920)
);

AND2x4_ASAP7_75t_L g5921 ( 
.A(n_5682),
.B(n_5425),
.Y(n_5921)
);

OA21x2_ASAP7_75t_L g5922 ( 
.A1(n_5749),
.A2(n_5393),
.B(n_5557),
.Y(n_5922)
);

OAI21x1_ASAP7_75t_L g5923 ( 
.A1(n_5742),
.A2(n_5556),
.B(n_5546),
.Y(n_5923)
);

OAI21x1_ASAP7_75t_L g5924 ( 
.A1(n_5594),
.A2(n_5556),
.B(n_5449),
.Y(n_5924)
);

BUFx2_ASAP7_75t_R g5925 ( 
.A(n_5609),
.Y(n_5925)
);

NOR2x1_ASAP7_75t_SL g5926 ( 
.A(n_5647),
.B(n_5556),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5602),
.Y(n_5927)
);

OAI21x1_ASAP7_75t_L g5928 ( 
.A1(n_5621),
.A2(n_5449),
.B(n_5557),
.Y(n_5928)
);

INVx2_ASAP7_75t_SL g5929 ( 
.A(n_5694),
.Y(n_5929)
);

AOI22xp33_ASAP7_75t_L g5930 ( 
.A1(n_5704),
.A2(n_2258),
.B1(n_2259),
.B2(n_2243),
.Y(n_5930)
);

OAI21x1_ASAP7_75t_L g5931 ( 
.A1(n_5621),
.A2(n_5449),
.B(n_5557),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5692),
.B(n_5695),
.Y(n_5932)
);

OA21x2_ASAP7_75t_L g5933 ( 
.A1(n_5643),
.A2(n_2702),
.B(n_2699),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5734),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5646),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5611),
.Y(n_5936)
);

AO21x2_ASAP7_75t_L g5937 ( 
.A1(n_5750),
.A2(n_2707),
.B(n_2699),
.Y(n_5937)
);

OAI21x1_ASAP7_75t_L g5938 ( 
.A1(n_5831),
.A2(n_5698),
.B(n_5633),
.Y(n_5938)
);

AO21x2_ASAP7_75t_L g5939 ( 
.A1(n_5801),
.A2(n_2708),
.B(n_2707),
.Y(n_5939)
);

OAI21x1_ASAP7_75t_L g5940 ( 
.A1(n_5831),
.A2(n_2844),
.B(n_2837),
.Y(n_5940)
);

NOR2xp67_ASAP7_75t_L g5941 ( 
.A(n_5686),
.B(n_82),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5664),
.Y(n_5942)
);

INVx1_ASAP7_75t_SL g5943 ( 
.A(n_5620),
.Y(n_5943)
);

OA21x2_ASAP7_75t_L g5944 ( 
.A1(n_5643),
.A2(n_2709),
.B(n_2708),
.Y(n_5944)
);

INVx3_ASAP7_75t_L g5945 ( 
.A(n_5753),
.Y(n_5945)
);

INVx3_ASAP7_75t_L g5946 ( 
.A(n_5689),
.Y(n_5946)
);

NAND2x1p5_ASAP7_75t_L g5947 ( 
.A(n_5640),
.B(n_5810),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5615),
.Y(n_5948)
);

OAI21x1_ASAP7_75t_L g5949 ( 
.A1(n_5625),
.A2(n_2844),
.B(n_2837),
.Y(n_5949)
);

OAI21x1_ASAP7_75t_L g5950 ( 
.A1(n_5736),
.A2(n_5676),
.B(n_5731),
.Y(n_5950)
);

AOI21x1_ASAP7_75t_L g5951 ( 
.A1(n_5617),
.A2(n_2709),
.B(n_83),
.Y(n_5951)
);

AND2x2_ASAP7_75t_SL g5952 ( 
.A(n_5776),
.B(n_84),
.Y(n_5952)
);

AO31x2_ASAP7_75t_L g5953 ( 
.A1(n_5612),
.A2(n_5777),
.A3(n_5779),
.B(n_5767),
.Y(n_5953)
);

INVxp67_ASAP7_75t_L g5954 ( 
.A(n_5783),
.Y(n_5954)
);

AOI21xp5_ASAP7_75t_L g5955 ( 
.A1(n_5622),
.A2(n_2497),
.B(n_2496),
.Y(n_5955)
);

OAI21x1_ASAP7_75t_L g5956 ( 
.A1(n_5733),
.A2(n_2844),
.B(n_2837),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5651),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5675),
.Y(n_5958)
);

OAI21x1_ASAP7_75t_L g5959 ( 
.A1(n_5733),
.A2(n_2882),
.B(n_2727),
.Y(n_5959)
);

NAND2x1p5_ASAP7_75t_L g5960 ( 
.A(n_5810),
.B(n_1267),
.Y(n_5960)
);

INVx2_ASAP7_75t_SL g5961 ( 
.A(n_5629),
.Y(n_5961)
);

BUFx10_ASAP7_75t_L g5962 ( 
.A(n_5825),
.Y(n_5962)
);

OAI21x1_ASAP7_75t_L g5963 ( 
.A1(n_5793),
.A2(n_2882),
.B(n_2727),
.Y(n_5963)
);

INVx3_ASAP7_75t_L g5964 ( 
.A(n_5689),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5683),
.Y(n_5965)
);

OAI21x1_ASAP7_75t_L g5966 ( 
.A1(n_5797),
.A2(n_2882),
.B(n_2727),
.Y(n_5966)
);

OAI21xp5_ASAP7_75t_L g5967 ( 
.A1(n_5624),
.A2(n_84),
.B(n_85),
.Y(n_5967)
);

OAI21x1_ASAP7_75t_L g5968 ( 
.A1(n_5800),
.A2(n_2882),
.B(n_2722),
.Y(n_5968)
);

INVx3_ASAP7_75t_L g5969 ( 
.A(n_5693),
.Y(n_5969)
);

BUFx6f_ASAP7_75t_L g5970 ( 
.A(n_5629),
.Y(n_5970)
);

NOR2x1_ASAP7_75t_SL g5971 ( 
.A(n_5647),
.B(n_1470),
.Y(n_5971)
);

AO31x2_ASAP7_75t_L g5972 ( 
.A1(n_5612),
.A2(n_2067),
.A3(n_2175),
.B(n_2109),
.Y(n_5972)
);

AOI21xp5_ASAP7_75t_L g5973 ( 
.A1(n_5622),
.A2(n_2497),
.B(n_2496),
.Y(n_5973)
);

OA21x2_ASAP7_75t_L g5974 ( 
.A1(n_5686),
.A2(n_86),
.B(n_87),
.Y(n_5974)
);

OAI21x1_ASAP7_75t_L g5975 ( 
.A1(n_5679),
.A2(n_2733),
.B(n_2730),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5684),
.Y(n_5976)
);

INVx1_ASAP7_75t_SL g5977 ( 
.A(n_5620),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_5657),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5708),
.Y(n_5979)
);

OA21x2_ASAP7_75t_L g5980 ( 
.A1(n_5710),
.A2(n_86),
.B(n_88),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5728),
.Y(n_5981)
);

NAND2x1p5_ASAP7_75t_L g5982 ( 
.A(n_5810),
.B(n_1470),
.Y(n_5982)
);

OAI21x1_ASAP7_75t_SL g5983 ( 
.A1(n_5618),
.A2(n_89),
.B(n_91),
.Y(n_5983)
);

OAI21x1_ASAP7_75t_L g5984 ( 
.A1(n_5766),
.A2(n_2733),
.B(n_2730),
.Y(n_5984)
);

INVx2_ASAP7_75t_L g5985 ( 
.A(n_5795),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5741),
.Y(n_5986)
);

INVxp67_ASAP7_75t_SL g5987 ( 
.A(n_5614),
.Y(n_5987)
);

BUFx2_ASAP7_75t_L g5988 ( 
.A(n_5789),
.Y(n_5988)
);

OAI21x1_ASAP7_75t_SL g5989 ( 
.A1(n_5652),
.A2(n_91),
.B(n_93),
.Y(n_5989)
);

INVx1_ASAP7_75t_SL g5990 ( 
.A(n_5781),
.Y(n_5990)
);

OAI21x1_ASAP7_75t_L g5991 ( 
.A1(n_5716),
.A2(n_2733),
.B(n_2730),
.Y(n_5991)
);

CKINVDCx11_ASAP7_75t_R g5992 ( 
.A(n_5721),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5699),
.Y(n_5993)
);

OR2x2_ASAP7_75t_L g5994 ( 
.A(n_5723),
.B(n_94),
.Y(n_5994)
);

INVx2_ASAP7_75t_L g5995 ( 
.A(n_5636),
.Y(n_5995)
);

NAND2xp5_ASAP7_75t_L g5996 ( 
.A(n_5638),
.B(n_94),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5699),
.Y(n_5997)
);

AOI21xp5_ASAP7_75t_L g5998 ( 
.A1(n_5680),
.A2(n_2497),
.B(n_2496),
.Y(n_5998)
);

INVx5_ASAP7_75t_L g5999 ( 
.A(n_5712),
.Y(n_5999)
);

OAI21x1_ASAP7_75t_L g6000 ( 
.A1(n_5715),
.A2(n_2761),
.B(n_2733),
.Y(n_6000)
);

NAND3xp33_ASAP7_75t_L g6001 ( 
.A(n_5642),
.B(n_2232),
.C(n_2229),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5691),
.B(n_95),
.Y(n_6002)
);

OA21x2_ASAP7_75t_L g6003 ( 
.A1(n_5710),
.A2(n_96),
.B(n_97),
.Y(n_6003)
);

OR2x6_ASAP7_75t_L g6004 ( 
.A(n_5780),
.B(n_2496),
.Y(n_6004)
);

OAI21x1_ASAP7_75t_L g6005 ( 
.A1(n_5678),
.A2(n_2767),
.B(n_2761),
.Y(n_6005)
);

INVx2_ASAP7_75t_L g6006 ( 
.A(n_5636),
.Y(n_6006)
);

INVx8_ASAP7_75t_L g6007 ( 
.A(n_5717),
.Y(n_6007)
);

AND2x4_ASAP7_75t_L g6008 ( 
.A(n_5682),
.B(n_97),
.Y(n_6008)
);

INVx5_ASAP7_75t_L g6009 ( 
.A(n_5687),
.Y(n_6009)
);

AND2x4_ASAP7_75t_L g6010 ( 
.A(n_5682),
.B(n_98),
.Y(n_6010)
);

OAI21x1_ASAP7_75t_L g6011 ( 
.A1(n_5720),
.A2(n_2767),
.B(n_2761),
.Y(n_6011)
);

OAI21x1_ASAP7_75t_L g6012 ( 
.A1(n_5656),
.A2(n_2767),
.B(n_2761),
.Y(n_6012)
);

AND2x4_ASAP7_75t_L g6013 ( 
.A(n_5724),
.B(n_100),
.Y(n_6013)
);

OAI21x1_ASAP7_75t_L g6014 ( 
.A1(n_5739),
.A2(n_2769),
.B(n_2767),
.Y(n_6014)
);

AO31x2_ASAP7_75t_L g6015 ( 
.A1(n_5596),
.A2(n_5836),
.A3(n_5834),
.B(n_5799),
.Y(n_6015)
);

OAI21x1_ASAP7_75t_L g6016 ( 
.A1(n_5685),
.A2(n_2795),
.B(n_2769),
.Y(n_6016)
);

OAI21x1_ASAP7_75t_L g6017 ( 
.A1(n_5661),
.A2(n_5599),
.B(n_5674),
.Y(n_6017)
);

BUFx3_ASAP7_75t_L g6018 ( 
.A(n_5809),
.Y(n_6018)
);

NOR2x1_ASAP7_75t_R g6019 ( 
.A(n_5717),
.B(n_100),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5696),
.Y(n_6020)
);

AO21x2_ASAP7_75t_L g6021 ( 
.A1(n_5589),
.A2(n_2125),
.B(n_101),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5696),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5723),
.Y(n_6023)
);

AOI21x1_ASAP7_75t_L g6024 ( 
.A1(n_5821),
.A2(n_5816),
.B(n_5819),
.Y(n_6024)
);

INVx2_ASAP7_75t_L g6025 ( 
.A(n_5796),
.Y(n_6025)
);

HB1xp67_ASAP7_75t_L g6026 ( 
.A(n_5614),
.Y(n_6026)
);

AOI21xp33_ASAP7_75t_SL g6027 ( 
.A1(n_5638),
.A2(n_103),
.B(n_104),
.Y(n_6027)
);

OA21x2_ASAP7_75t_L g6028 ( 
.A1(n_5807),
.A2(n_104),
.B(n_105),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5735),
.Y(n_6029)
);

AO21x2_ASAP7_75t_L g6030 ( 
.A1(n_5589),
.A2(n_105),
.B(n_106),
.Y(n_6030)
);

AND2x4_ASAP7_75t_L g6031 ( 
.A(n_5724),
.B(n_106),
.Y(n_6031)
);

INVx4_ASAP7_75t_L g6032 ( 
.A(n_5717),
.Y(n_6032)
);

OR2x2_ASAP7_75t_L g6033 ( 
.A(n_5819),
.B(n_107),
.Y(n_6033)
);

BUFx3_ASAP7_75t_L g6034 ( 
.A(n_5809),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5607),
.B(n_107),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5759),
.Y(n_6036)
);

NOR2xp67_ASAP7_75t_L g6037 ( 
.A(n_5717),
.B(n_5722),
.Y(n_6037)
);

CKINVDCx11_ASAP7_75t_R g6038 ( 
.A(n_5721),
.Y(n_6038)
);

OA21x2_ASAP7_75t_L g6039 ( 
.A1(n_5814),
.A2(n_109),
.B(n_110),
.Y(n_6039)
);

OA21x2_ASAP7_75t_L g6040 ( 
.A1(n_5616),
.A2(n_109),
.B(n_112),
.Y(n_6040)
);

AOI21xp5_ASAP7_75t_L g6041 ( 
.A1(n_5680),
.A2(n_2497),
.B(n_2496),
.Y(n_6041)
);

AO21x2_ASAP7_75t_L g6042 ( 
.A1(n_5822),
.A2(n_113),
.B(n_114),
.Y(n_6042)
);

HB1xp67_ASAP7_75t_L g6043 ( 
.A(n_5669),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5607),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5772),
.B(n_113),
.Y(n_6045)
);

BUFx2_ASAP7_75t_L g6046 ( 
.A(n_5693),
.Y(n_6046)
);

AND2x2_ASAP7_75t_L g6047 ( 
.A(n_5610),
.B(n_115),
.Y(n_6047)
);

OAI21x1_ASAP7_75t_L g6048 ( 
.A1(n_5745),
.A2(n_5667),
.B(n_5688),
.Y(n_6048)
);

OAI21x1_ASAP7_75t_L g6049 ( 
.A1(n_5650),
.A2(n_2815),
.B(n_2128),
.Y(n_6049)
);

AO31x2_ASAP7_75t_L g6050 ( 
.A1(n_5596),
.A2(n_2067),
.A3(n_2175),
.B(n_2109),
.Y(n_6050)
);

OR2x6_ASAP7_75t_L g6051 ( 
.A(n_5780),
.B(n_2497),
.Y(n_6051)
);

OAI21xp5_ASAP7_75t_L g6052 ( 
.A1(n_5670),
.A2(n_116),
.B(n_117),
.Y(n_6052)
);

OAI21x1_ASAP7_75t_L g6053 ( 
.A1(n_5650),
.A2(n_2815),
.B(n_2128),
.Y(n_6053)
);

OAI21x1_ASAP7_75t_L g6054 ( 
.A1(n_5605),
.A2(n_2815),
.B(n_2128),
.Y(n_6054)
);

BUFx12f_ASAP7_75t_L g6055 ( 
.A(n_5817),
.Y(n_6055)
);

NOR2xp33_ASAP7_75t_L g6056 ( 
.A(n_5758),
.B(n_118),
.Y(n_6056)
);

OAI21x1_ASAP7_75t_L g6057 ( 
.A1(n_5605),
.A2(n_2171),
.B(n_2165),
.Y(n_6057)
);

AO31x2_ASAP7_75t_L g6058 ( 
.A1(n_5756),
.A2(n_2067),
.A3(n_2175),
.B(n_2109),
.Y(n_6058)
);

CKINVDCx20_ASAP7_75t_R g6059 ( 
.A(n_5781),
.Y(n_6059)
);

AO21x2_ASAP7_75t_L g6060 ( 
.A1(n_5826),
.A2(n_119),
.B(n_120),
.Y(n_6060)
);

OAI21x1_ASAP7_75t_L g6061 ( 
.A1(n_5762),
.A2(n_2171),
.B(n_2165),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_L g6062 ( 
.A(n_5669),
.B(n_121),
.Y(n_6062)
);

AND2x2_ASAP7_75t_L g6063 ( 
.A(n_5832),
.B(n_121),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_5757),
.B(n_122),
.Y(n_6064)
);

A2O1A1Ixp33_ASAP7_75t_L g6065 ( 
.A1(n_5857),
.A2(n_5756),
.B(n_5806),
.C(n_5790),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5946),
.B(n_5832),
.Y(n_6066)
);

OAI22xp5_ASAP7_75t_L g6067 ( 
.A1(n_5869),
.A2(n_5670),
.B1(n_5642),
.B2(n_5608),
.Y(n_6067)
);

AOI21x1_ASAP7_75t_SL g6068 ( 
.A1(n_5894),
.A2(n_5738),
.B(n_5722),
.Y(n_6068)
);

NOR2xp67_ASAP7_75t_L g6069 ( 
.A(n_5862),
.B(n_5722),
.Y(n_6069)
);

NAND2xp5_ASAP7_75t_L g6070 ( 
.A(n_5912),
.B(n_5790),
.Y(n_6070)
);

AOI21x1_ASAP7_75t_SL g6071 ( 
.A1(n_5870),
.A2(n_5738),
.B(n_5722),
.Y(n_6071)
);

OAI22xp5_ASAP7_75t_L g6072 ( 
.A1(n_5869),
.A2(n_5598),
.B1(n_5649),
.B2(n_5829),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_5912),
.B(n_5806),
.Y(n_6073)
);

NAND2xp5_ASAP7_75t_L g6074 ( 
.A(n_5917),
.B(n_5719),
.Y(n_6074)
);

A2O1A1Ixp33_ASAP7_75t_L g6075 ( 
.A1(n_6052),
.A2(n_5628),
.B(n_5677),
.C(n_5746),
.Y(n_6075)
);

OR2x2_ASAP7_75t_L g6076 ( 
.A(n_5859),
.B(n_6025),
.Y(n_6076)
);

OAI22xp5_ASAP7_75t_L g6077 ( 
.A1(n_5893),
.A2(n_6062),
.B1(n_5908),
.B2(n_6051),
.Y(n_6077)
);

CKINVDCx11_ASAP7_75t_R g6078 ( 
.A(n_5992),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5932),
.Y(n_6079)
);

OAI22xp5_ASAP7_75t_L g6080 ( 
.A1(n_5908),
.A2(n_5623),
.B1(n_5705),
.B2(n_5735),
.Y(n_6080)
);

OA21x2_ASAP7_75t_L g6081 ( 
.A1(n_5987),
.A2(n_5938),
.B(n_6043),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5954),
.B(n_5768),
.Y(n_6082)
);

HB1xp67_ASAP7_75t_L g6083 ( 
.A(n_5985),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5932),
.Y(n_6084)
);

AOI21x1_ASAP7_75t_SL g6085 ( 
.A1(n_5870),
.A2(n_5687),
.B(n_5817),
.Y(n_6085)
);

AOI21xp5_ASAP7_75t_SL g6086 ( 
.A1(n_6019),
.A2(n_5746),
.B(n_5623),
.Y(n_6086)
);

AOI21xp5_ASAP7_75t_SL g6087 ( 
.A1(n_5974),
.A2(n_5735),
.B(n_5828),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5974),
.Y(n_6088)
);

AOI21xp5_ASAP7_75t_L g6089 ( 
.A1(n_6052),
.A2(n_5755),
.B(n_5681),
.Y(n_6089)
);

AND2x2_ASAP7_75t_L g6090 ( 
.A(n_5964),
.B(n_5839),
.Y(n_6090)
);

NAND2xp5_ASAP7_75t_L g6091 ( 
.A(n_6023),
.B(n_5780),
.Y(n_6091)
);

AND2x4_ASAP7_75t_L g6092 ( 
.A(n_5969),
.B(n_5774),
.Y(n_6092)
);

O2A1O1Ixp33_ASAP7_75t_L g6093 ( 
.A1(n_6027),
.A2(n_5840),
.B(n_5838),
.C(n_5681),
.Y(n_6093)
);

AOI21xp5_ASAP7_75t_L g6094 ( 
.A1(n_5967),
.A2(n_5755),
.B(n_5649),
.Y(n_6094)
);

AND2x2_ASAP7_75t_L g6095 ( 
.A(n_6046),
.B(n_5839),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5935),
.Y(n_6096)
);

BUFx12f_ASAP7_75t_L g6097 ( 
.A(n_5992),
.Y(n_6097)
);

AOI21xp5_ASAP7_75t_L g6098 ( 
.A1(n_5967),
.A2(n_5838),
.B(n_5794),
.Y(n_6098)
);

NAND2xp5_ASAP7_75t_L g6099 ( 
.A(n_5902),
.B(n_5665),
.Y(n_6099)
);

A2O1A1Ixp33_ASAP7_75t_L g6100 ( 
.A1(n_5876),
.A2(n_5740),
.B(n_5792),
.C(n_5804),
.Y(n_6100)
);

OAI22xp5_ASAP7_75t_SL g6101 ( 
.A1(n_5943),
.A2(n_5770),
.B1(n_5810),
.B2(n_5828),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_5902),
.B(n_5729),
.Y(n_6102)
);

AOI21xp5_ASAP7_75t_SL g6103 ( 
.A1(n_5980),
.A2(n_5830),
.B(n_5813),
.Y(n_6103)
);

NAND2xp5_ASAP7_75t_L g6104 ( 
.A(n_6044),
.B(n_5634),
.Y(n_6104)
);

AND2x2_ASAP7_75t_L g6105 ( 
.A(n_5945),
.B(n_5905),
.Y(n_6105)
);

AOI21xp5_ASAP7_75t_SL g6106 ( 
.A1(n_5980),
.A2(n_5830),
.B(n_5813),
.Y(n_6106)
);

OR2x2_ASAP7_75t_L g6107 ( 
.A(n_5884),
.B(n_5634),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_5927),
.B(n_5771),
.Y(n_6108)
);

INVx2_ASAP7_75t_L g6109 ( 
.A(n_6003),
.Y(n_6109)
);

OAI22xp5_ASAP7_75t_L g6110 ( 
.A1(n_5908),
.A2(n_5595),
.B1(n_5788),
.B2(n_5760),
.Y(n_6110)
);

AND2x2_ASAP7_75t_L g6111 ( 
.A(n_5921),
.B(n_5760),
.Y(n_6111)
);

AOI21xp5_ASAP7_75t_L g6112 ( 
.A1(n_5998),
.A2(n_6041),
.B(n_5848),
.Y(n_6112)
);

INVxp67_ASAP7_75t_L g6113 ( 
.A(n_5925),
.Y(n_6113)
);

OAI22xp5_ASAP7_75t_L g6114 ( 
.A1(n_6004),
.A2(n_5702),
.B1(n_5703),
.B2(n_5714),
.Y(n_6114)
);

HB1xp67_ASAP7_75t_L g6115 ( 
.A(n_5889),
.Y(n_6115)
);

O2A1O1Ixp33_ASAP7_75t_L g6116 ( 
.A1(n_6027),
.A2(n_5794),
.B(n_5702),
.C(n_5703),
.Y(n_6116)
);

NAND2xp5_ASAP7_75t_L g6117 ( 
.A(n_5855),
.B(n_5823),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5942),
.Y(n_6118)
);

O2A1O1Ixp33_ASAP7_75t_L g6119 ( 
.A1(n_5876),
.A2(n_5848),
.B(n_5863),
.C(n_5878),
.Y(n_6119)
);

NAND2xp5_ASAP7_75t_L g6120 ( 
.A(n_5855),
.B(n_5823),
.Y(n_6120)
);

OA22x2_ASAP7_75t_L g6121 ( 
.A1(n_5844),
.A2(n_5690),
.B1(n_5754),
.B2(n_5752),
.Y(n_6121)
);

HB1xp67_ASAP7_75t_L g6122 ( 
.A(n_5899),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5958),
.Y(n_6123)
);

HB1xp67_ASAP7_75t_L g6124 ( 
.A(n_5849),
.Y(n_6124)
);

AOI21xp5_ASAP7_75t_SL g6125 ( 
.A1(n_6003),
.A2(n_5778),
.B(n_5773),
.Y(n_6125)
);

AOI21xp5_ASAP7_75t_L g6126 ( 
.A1(n_5998),
.A2(n_6041),
.B(n_5977),
.Y(n_6126)
);

AOI21xp5_ASAP7_75t_L g6127 ( 
.A1(n_5943),
.A2(n_5654),
.B(n_5725),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5965),
.Y(n_6128)
);

OA21x2_ASAP7_75t_L g6129 ( 
.A1(n_5987),
.A2(n_5730),
.B(n_5732),
.Y(n_6129)
);

BUFx2_ASAP7_75t_L g6130 ( 
.A(n_6055),
.Y(n_6130)
);

OA21x2_ASAP7_75t_L g6131 ( 
.A1(n_6043),
.A2(n_5815),
.B(n_5812),
.Y(n_6131)
);

HB1xp67_ASAP7_75t_L g6132 ( 
.A(n_5873),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5976),
.Y(n_6133)
);

INVx1_ASAP7_75t_SL g6134 ( 
.A(n_5977),
.Y(n_6134)
);

OA21x2_ASAP7_75t_L g6135 ( 
.A1(n_5874),
.A2(n_5782),
.B(n_5751),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_5934),
.B(n_5835),
.Y(n_6136)
);

O2A1O1Ixp5_ASAP7_75t_L g6137 ( 
.A1(n_5871),
.A2(n_5654),
.B(n_5658),
.C(n_5641),
.Y(n_6137)
);

OA22x2_ASAP7_75t_L g6138 ( 
.A1(n_5844),
.A2(n_5761),
.B1(n_5726),
.B2(n_5747),
.Y(n_6138)
);

INVx2_ASAP7_75t_L g6139 ( 
.A(n_5953),
.Y(n_6139)
);

NAND2xp5_ASAP7_75t_L g6140 ( 
.A(n_5907),
.B(n_5641),
.Y(n_6140)
);

BUFx6f_ASAP7_75t_L g6141 ( 
.A(n_5865),
.Y(n_6141)
);

OAI22xp5_ASAP7_75t_L g6142 ( 
.A1(n_6051),
.A2(n_5658),
.B1(n_5725),
.B2(n_5655),
.Y(n_6142)
);

A2O1A1Ixp33_ASAP7_75t_L g6143 ( 
.A1(n_5845),
.A2(n_5764),
.B(n_5765),
.C(n_5820),
.Y(n_6143)
);

A2O1A1Ixp33_ASAP7_75t_L g6144 ( 
.A1(n_5845),
.A2(n_5824),
.B(n_5837),
.C(n_5827),
.Y(n_6144)
);

BUFx6f_ASAP7_75t_L g6145 ( 
.A(n_5865),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5979),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_5907),
.B(n_5833),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_5947),
.B(n_5763),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5953),
.Y(n_6149)
);

AO21x2_ASAP7_75t_L g6150 ( 
.A1(n_6026),
.A2(n_5645),
.B(n_5763),
.Y(n_6150)
);

OA21x2_ASAP7_75t_L g6151 ( 
.A1(n_6020),
.A2(n_5842),
.B(n_5841),
.Y(n_6151)
);

AND2x2_ASAP7_75t_L g6152 ( 
.A(n_6009),
.B(n_5655),
.Y(n_6152)
);

AOI221xp5_ASAP7_75t_L g6153 ( 
.A1(n_6026),
.A2(n_5645),
.B1(n_2243),
.B2(n_2262),
.C(n_2259),
.Y(n_6153)
);

OAI22xp5_ASAP7_75t_L g6154 ( 
.A1(n_6051),
.A2(n_5952),
.B1(n_5886),
.B2(n_6008),
.Y(n_6154)
);

HB1xp67_ASAP7_75t_L g6155 ( 
.A(n_5986),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5981),
.Y(n_6156)
);

BUFx3_ASAP7_75t_L g6157 ( 
.A(n_5883),
.Y(n_6157)
);

AND2x2_ASAP7_75t_L g6158 ( 
.A(n_6009),
.B(n_5787),
.Y(n_6158)
);

OAI22xp5_ASAP7_75t_L g6159 ( 
.A1(n_5886),
.A2(n_127),
.B1(n_123),
.B2(n_124),
.Y(n_6159)
);

AND2x4_ASAP7_75t_L g6160 ( 
.A(n_5862),
.B(n_6037),
.Y(n_6160)
);

A2O1A1Ixp33_ASAP7_75t_L g6161 ( 
.A1(n_6056),
.A2(n_5784),
.B(n_5802),
.C(n_5791),
.Y(n_6161)
);

OA21x2_ASAP7_75t_L g6162 ( 
.A1(n_5993),
.A2(n_5803),
.B(n_5805),
.Y(n_6162)
);

BUFx2_ASAP7_75t_L g6163 ( 
.A(n_5883),
.Y(n_6163)
);

CKINVDCx20_ASAP7_75t_R g6164 ( 
.A(n_6038),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_5862),
.B(n_5808),
.Y(n_6165)
);

NOR2xp67_ASAP7_75t_L g6166 ( 
.A(n_5862),
.B(n_124),
.Y(n_6166)
);

INVx2_ASAP7_75t_L g6167 ( 
.A(n_5953),
.Y(n_6167)
);

AND2x2_ASAP7_75t_L g6168 ( 
.A(n_6009),
.B(n_5918),
.Y(n_6168)
);

OA21x2_ASAP7_75t_L g6169 ( 
.A1(n_5997),
.A2(n_128),
.B(n_130),
.Y(n_6169)
);

BUFx3_ASAP7_75t_L g6170 ( 
.A(n_5846),
.Y(n_6170)
);

HB1xp67_ASAP7_75t_L g6171 ( 
.A(n_6040),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5852),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5872),
.Y(n_6173)
);

NOR2xp67_ASAP7_75t_L g6174 ( 
.A(n_6032),
.B(n_131),
.Y(n_6174)
);

INVx3_ASAP7_75t_L g6175 ( 
.A(n_6032),
.Y(n_6175)
);

O2A1O1Ixp5_ASAP7_75t_L g6176 ( 
.A1(n_6024),
.A2(n_135),
.B(n_132),
.C(n_134),
.Y(n_6176)
);

OA21x2_ASAP7_75t_L g6177 ( 
.A1(n_6022),
.A2(n_132),
.B(n_134),
.Y(n_6177)
);

A2O1A1Ixp33_ASAP7_75t_L g6178 ( 
.A1(n_6056),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_6178)
);

AND2x4_ASAP7_75t_L g6179 ( 
.A(n_6037),
.B(n_139),
.Y(n_6179)
);

HB1xp67_ASAP7_75t_L g6180 ( 
.A(n_6040),
.Y(n_6180)
);

AOI21xp5_ASAP7_75t_L g6181 ( 
.A1(n_5996),
.A2(n_139),
.B(n_140),
.Y(n_6181)
);

AND2x2_ASAP7_75t_L g6182 ( 
.A(n_6009),
.B(n_140),
.Y(n_6182)
);

NAND2xp5_ASAP7_75t_L g6183 ( 
.A(n_5919),
.B(n_5996),
.Y(n_6183)
);

INVx5_ASAP7_75t_L g6184 ( 
.A(n_5865),
.Y(n_6184)
);

AOI21x1_ASAP7_75t_SL g6185 ( 
.A1(n_5877),
.A2(n_6064),
.B(n_6035),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5872),
.Y(n_6186)
);

AND2x2_ASAP7_75t_L g6187 ( 
.A(n_5880),
.B(n_142),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_6028),
.Y(n_6188)
);

O2A1O1Ixp33_ASAP7_75t_L g6189 ( 
.A1(n_5863),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_6189)
);

A2O1A1Ixp33_ASAP7_75t_L g6190 ( 
.A1(n_5878),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_5929),
.B(n_146),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_L g6192 ( 
.A(n_5937),
.B(n_147),
.Y(n_6192)
);

BUFx3_ASAP7_75t_L g6193 ( 
.A(n_5853),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_6028),
.Y(n_6194)
);

AND2x2_ASAP7_75t_L g6195 ( 
.A(n_5898),
.B(n_148),
.Y(n_6195)
);

INVx3_ASAP7_75t_L g6196 ( 
.A(n_5909),
.Y(n_6196)
);

O2A1O1Ixp33_ASAP7_75t_L g6197 ( 
.A1(n_6035),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_6197)
);

BUFx6f_ASAP7_75t_L g6198 ( 
.A(n_5909),
.Y(n_6198)
);

OR2x2_ASAP7_75t_L g6199 ( 
.A(n_5916),
.B(n_152),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_5898),
.B(n_153),
.Y(n_6200)
);

BUFx3_ASAP7_75t_L g6201 ( 
.A(n_6059),
.Y(n_6201)
);

AND2x4_ASAP7_75t_L g6202 ( 
.A(n_6008),
.B(n_154),
.Y(n_6202)
);

OAI22xp5_ASAP7_75t_L g6203 ( 
.A1(n_5994),
.A2(n_158),
.B1(n_155),
.B2(n_156),
.Y(n_6203)
);

CKINVDCx5p33_ASAP7_75t_R g6204 ( 
.A(n_5906),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_6039),
.Y(n_6205)
);

NOR2xp67_ASAP7_75t_L g6206 ( 
.A(n_5856),
.B(n_158),
.Y(n_6206)
);

OA21x2_ASAP7_75t_L g6207 ( 
.A1(n_5995),
.A2(n_159),
.B(n_160),
.Y(n_6207)
);

OA21x2_ASAP7_75t_L g6208 ( 
.A1(n_6006),
.A2(n_159),
.B(n_161),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_6039),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_6015),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_6015),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_6015),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_6033),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_5911),
.B(n_6002),
.Y(n_6214)
);

AND2x2_ASAP7_75t_L g6215 ( 
.A(n_5911),
.B(n_163),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_5988),
.B(n_165),
.Y(n_6216)
);

OAI22xp5_ASAP7_75t_L g6217 ( 
.A1(n_6010),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_6217)
);

OAI22xp5_ASAP7_75t_L g6218 ( 
.A1(n_6010),
.A2(n_170),
.B1(n_167),
.B2(n_168),
.Y(n_6218)
);

OA22x2_ASAP7_75t_L g6219 ( 
.A1(n_5854),
.A2(n_173),
.B1(n_168),
.B2(n_172),
.Y(n_6219)
);

OA21x2_ASAP7_75t_L g6220 ( 
.A1(n_5890),
.A2(n_174),
.B(n_176),
.Y(n_6220)
);

O2A1O1Ixp33_ASAP7_75t_L g6221 ( 
.A1(n_5989),
.A2(n_178),
.B(n_174),
.C(n_177),
.Y(n_6221)
);

O2A1O1Ixp5_ASAP7_75t_L g6222 ( 
.A1(n_5901),
.A2(n_182),
.B(n_179),
.C(n_180),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5903),
.Y(n_6223)
);

BUFx6f_ASAP7_75t_L g6224 ( 
.A(n_5909),
.Y(n_6224)
);

OAI22xp5_ASAP7_75t_L g6225 ( 
.A1(n_5897),
.A2(n_183),
.B1(n_179),
.B2(n_180),
.Y(n_6225)
);

AND2x2_ASAP7_75t_L g6226 ( 
.A(n_5990),
.B(n_183),
.Y(n_6226)
);

OAI22xp5_ASAP7_75t_L g6227 ( 
.A1(n_5897),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_6227)
);

AOI21xp5_ASAP7_75t_SL g6228 ( 
.A1(n_5971),
.A2(n_184),
.B(n_186),
.Y(n_6228)
);

OAI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_5920),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_6030),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_5866),
.B(n_188),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_5915),
.Y(n_6232)
);

AOI21xp5_ASAP7_75t_L g6233 ( 
.A1(n_5896),
.A2(n_5926),
.B(n_6007),
.Y(n_6233)
);

NAND2xp5_ASAP7_75t_L g6234 ( 
.A(n_5867),
.B(n_192),
.Y(n_6234)
);

INVx2_ASAP7_75t_L g6235 ( 
.A(n_5939),
.Y(n_6235)
);

AND2x2_ASAP7_75t_L g6236 ( 
.A(n_5990),
.B(n_5961),
.Y(n_6236)
);

AND2x2_ASAP7_75t_L g6237 ( 
.A(n_5892),
.B(n_193),
.Y(n_6237)
);

A2O1A1Ixp33_ASAP7_75t_L g6238 ( 
.A1(n_5941),
.A2(n_197),
.B(n_194),
.C(n_195),
.Y(n_6238)
);

NAND2xp5_ASAP7_75t_L g6239 ( 
.A(n_5867),
.B(n_198),
.Y(n_6239)
);

AND2x2_ASAP7_75t_L g6240 ( 
.A(n_6047),
.B(n_198),
.Y(n_6240)
);

OAI22xp5_ASAP7_75t_L g6241 ( 
.A1(n_5854),
.A2(n_203),
.B1(n_200),
.B2(n_202),
.Y(n_6241)
);

HB1xp67_ASAP7_75t_L g6242 ( 
.A(n_5951),
.Y(n_6242)
);

AND2x2_ASAP7_75t_L g6243 ( 
.A(n_6045),
.B(n_205),
.Y(n_6243)
);

CKINVDCx5p33_ASAP7_75t_R g6244 ( 
.A(n_6018),
.Y(n_6244)
);

AND2x2_ASAP7_75t_L g6245 ( 
.A(n_6034),
.B(n_207),
.Y(n_6245)
);

AOI21xp5_ASAP7_75t_SL g6246 ( 
.A1(n_6013),
.A2(n_209),
.B(n_211),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_5915),
.Y(n_6247)
);

OA22x2_ASAP7_75t_L g6248 ( 
.A1(n_5854),
.A2(n_6031),
.B1(n_6013),
.B2(n_5983),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_5867),
.B(n_212),
.Y(n_6249)
);

NAND2xp5_ASAP7_75t_L g6250 ( 
.A(n_6058),
.B(n_213),
.Y(n_6250)
);

AND2x2_ASAP7_75t_L g6251 ( 
.A(n_5999),
.B(n_213),
.Y(n_6251)
);

A2O1A1Ixp33_ASAP7_75t_L g6252 ( 
.A1(n_5941),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_6252)
);

AOI211xp5_ASAP7_75t_L g6253 ( 
.A1(n_5955),
.A2(n_218),
.B(n_215),
.C(n_217),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_6058),
.B(n_6031),
.Y(n_6254)
);

INVx2_ASAP7_75t_L g6255 ( 
.A(n_5939),
.Y(n_6255)
);

O2A1O1Ixp33_ASAP7_75t_L g6256 ( 
.A1(n_6042),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_6256)
);

OAI22xp5_ASAP7_75t_L g6257 ( 
.A1(n_5920),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_6257)
);

O2A1O1Ixp33_ASAP7_75t_L g6258 ( 
.A1(n_6042),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_6258)
);

OA21x2_ASAP7_75t_L g6259 ( 
.A1(n_5950),
.A2(n_6017),
.B(n_5923),
.Y(n_6259)
);

NOR2x1_ASAP7_75t_SL g6260 ( 
.A(n_5999),
.B(n_1518),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_5999),
.B(n_226),
.Y(n_6261)
);

INVx2_ASAP7_75t_SL g6262 ( 
.A(n_5999),
.Y(n_6262)
);

INVx2_ASAP7_75t_L g6263 ( 
.A(n_6029),
.Y(n_6263)
);

AOI21xp5_ASAP7_75t_SL g6264 ( 
.A1(n_6021),
.A2(n_229),
.B(n_230),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5847),
.Y(n_6265)
);

INVx2_ASAP7_75t_L g6266 ( 
.A(n_6163),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_6155),
.Y(n_6267)
);

INVx2_ASAP7_75t_L g6268 ( 
.A(n_6157),
.Y(n_6268)
);

AND2x2_ASAP7_75t_L g6269 ( 
.A(n_6111),
.B(n_5970),
.Y(n_6269)
);

BUFx2_ASAP7_75t_L g6270 ( 
.A(n_6097),
.Y(n_6270)
);

INVx2_ASAP7_75t_L g6271 ( 
.A(n_6134),
.Y(n_6271)
);

OAI21x1_ASAP7_75t_L g6272 ( 
.A1(n_6140),
.A2(n_5924),
.B(n_6054),
.Y(n_6272)
);

INVx2_ASAP7_75t_L g6273 ( 
.A(n_6177),
.Y(n_6273)
);

NAND2xp5_ASAP7_75t_L g6274 ( 
.A(n_6072),
.B(n_5888),
.Y(n_6274)
);

OR2x6_ASAP7_75t_L g6275 ( 
.A(n_6119),
.B(n_6007),
.Y(n_6275)
);

NAND2xp5_ASAP7_75t_L g6276 ( 
.A(n_6072),
.B(n_5888),
.Y(n_6276)
);

NAND2xp5_ASAP7_75t_L g6277 ( 
.A(n_6067),
.B(n_6171),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_6177),
.Y(n_6278)
);

OAI21x1_ASAP7_75t_L g6279 ( 
.A1(n_6080),
.A2(n_6048),
.B(n_5851),
.Y(n_6279)
);

NOR2xp33_ASAP7_75t_L g6280 ( 
.A(n_6113),
.B(n_5925),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6115),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_6122),
.Y(n_6282)
);

AO21x2_ASAP7_75t_L g6283 ( 
.A1(n_6070),
.A2(n_6021),
.B(n_6001),
.Y(n_6283)
);

AND2x2_ASAP7_75t_L g6284 ( 
.A(n_6066),
.B(n_6063),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6124),
.Y(n_6285)
);

NOR2xp33_ASAP7_75t_L g6286 ( 
.A(n_6078),
.B(n_5962),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6132),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6096),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6118),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_6169),
.Y(n_6290)
);

INVx2_ASAP7_75t_L g6291 ( 
.A(n_6169),
.Y(n_6291)
);

BUFx6f_ASAP7_75t_L g6292 ( 
.A(n_6170),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_6236),
.B(n_5962),
.Y(n_6293)
);

NAND2x1p5_ASAP7_75t_L g6294 ( 
.A(n_6166),
.B(n_5875),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_6207),
.Y(n_6295)
);

OAI21x1_ASAP7_75t_L g6296 ( 
.A1(n_6137),
.A2(n_5860),
.B(n_5881),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6123),
.Y(n_6297)
);

INVx2_ASAP7_75t_L g6298 ( 
.A(n_6207),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6128),
.Y(n_6299)
);

INVx4_ASAP7_75t_L g6300 ( 
.A(n_6184),
.Y(n_6300)
);

AO21x2_ASAP7_75t_L g6301 ( 
.A1(n_6073),
.A2(n_5973),
.B(n_5879),
.Y(n_6301)
);

INVx2_ASAP7_75t_L g6302 ( 
.A(n_6208),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_6208),
.Y(n_6303)
);

INVx2_ASAP7_75t_SL g6304 ( 
.A(n_6201),
.Y(n_6304)
);

HB1xp67_ASAP7_75t_L g6305 ( 
.A(n_6180),
.Y(n_6305)
);

BUFx6f_ASAP7_75t_L g6306 ( 
.A(n_6193),
.Y(n_6306)
);

AO21x2_ASAP7_75t_L g6307 ( 
.A1(n_6231),
.A2(n_6239),
.B(n_6234),
.Y(n_6307)
);

OR2x2_ASAP7_75t_L g6308 ( 
.A(n_6183),
.B(n_6076),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_6220),
.Y(n_6309)
);

HB1xp67_ASAP7_75t_L g6310 ( 
.A(n_6067),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_6220),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_6133),
.Y(n_6312)
);

INVx4_ASAP7_75t_L g6313 ( 
.A(n_6184),
.Y(n_6313)
);

INVx3_ASAP7_75t_L g6314 ( 
.A(n_6160),
.Y(n_6314)
);

AND2x4_ASAP7_75t_L g6315 ( 
.A(n_6184),
.B(n_6060),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_6146),
.Y(n_6316)
);

INVx2_ASAP7_75t_L g6317 ( 
.A(n_6150),
.Y(n_6317)
);

AOI21x1_ASAP7_75t_L g6318 ( 
.A1(n_6130),
.A2(n_5850),
.B(n_5847),
.Y(n_6318)
);

INVx2_ASAP7_75t_L g6319 ( 
.A(n_6150),
.Y(n_6319)
);

INVxp67_ASAP7_75t_L g6320 ( 
.A(n_6249),
.Y(n_6320)
);

INVx2_ASAP7_75t_L g6321 ( 
.A(n_6088),
.Y(n_6321)
);

OR2x2_ASAP7_75t_L g6322 ( 
.A(n_6083),
.B(n_5972),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_6156),
.Y(n_6323)
);

AOI222xp33_ASAP7_75t_L g6324 ( 
.A1(n_6075),
.A2(n_6065),
.B1(n_6077),
.B2(n_6100),
.C1(n_6159),
.C2(n_6099),
.Y(n_6324)
);

HB1xp67_ASAP7_75t_L g6325 ( 
.A(n_6242),
.Y(n_6325)
);

INVx3_ASAP7_75t_L g6326 ( 
.A(n_6160),
.Y(n_6326)
);

INVx2_ASAP7_75t_L g6327 ( 
.A(n_6109),
.Y(n_6327)
);

INVx2_ASAP7_75t_SL g6328 ( 
.A(n_6164),
.Y(n_6328)
);

OR2x2_ASAP7_75t_L g6329 ( 
.A(n_6213),
.B(n_6079),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6081),
.Y(n_6330)
);

BUFx12f_ASAP7_75t_L g6331 ( 
.A(n_6204),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_6179),
.Y(n_6332)
);

INVx4_ASAP7_75t_L g6333 ( 
.A(n_6141),
.Y(n_6333)
);

INVx2_ASAP7_75t_L g6334 ( 
.A(n_6092),
.Y(n_6334)
);

INVx3_ASAP7_75t_L g6335 ( 
.A(n_6141),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6230),
.Y(n_6336)
);

AND2x4_ASAP7_75t_L g6337 ( 
.A(n_6196),
.B(n_5891),
.Y(n_6337)
);

INVx3_ASAP7_75t_L g6338 ( 
.A(n_6141),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_6188),
.Y(n_6339)
);

AND2x2_ASAP7_75t_L g6340 ( 
.A(n_6095),
.B(n_6005),
.Y(n_6340)
);

HB1xp67_ASAP7_75t_L g6341 ( 
.A(n_6081),
.Y(n_6341)
);

AO21x2_ASAP7_75t_L g6342 ( 
.A1(n_6127),
.A2(n_5879),
.B(n_5900),
.Y(n_6342)
);

BUFx3_ASAP7_75t_L g6343 ( 
.A(n_6145),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_6194),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_6205),
.Y(n_6345)
);

AOI21x1_ASAP7_75t_L g6346 ( 
.A1(n_6265),
.A2(n_5861),
.B(n_5933),
.Y(n_6346)
);

AO21x2_ASAP7_75t_L g6347 ( 
.A1(n_6147),
.A2(n_5900),
.B(n_6036),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_6209),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_6173),
.Y(n_6349)
);

NAND2xp5_ASAP7_75t_L g6350 ( 
.A(n_6094),
.B(n_5972),
.Y(n_6350)
);

OAI21xp5_ASAP7_75t_L g6351 ( 
.A1(n_6176),
.A2(n_5930),
.B(n_5960),
.Y(n_6351)
);

AOI22xp33_ASAP7_75t_L g6352 ( 
.A1(n_6089),
.A2(n_5882),
.B1(n_5864),
.B2(n_5885),
.Y(n_6352)
);

HB1xp67_ASAP7_75t_L g6353 ( 
.A(n_6074),
.Y(n_6353)
);

NOR2x1_ASAP7_75t_SL g6354 ( 
.A(n_6154),
.B(n_5858),
.Y(n_6354)
);

NAND2xp5_ASAP7_75t_L g6355 ( 
.A(n_6084),
.B(n_5972),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_6105),
.B(n_5904),
.Y(n_6356)
);

OR2x2_ASAP7_75t_L g6357 ( 
.A(n_6186),
.B(n_6050),
.Y(n_6357)
);

INVx2_ASAP7_75t_L g6358 ( 
.A(n_6145),
.Y(n_6358)
);

INVxp67_ASAP7_75t_SL g6359 ( 
.A(n_6189),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_6192),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_6198),
.Y(n_6361)
);

INVx2_ASAP7_75t_L g6362 ( 
.A(n_6198),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_6199),
.Y(n_6363)
);

INVx3_ASAP7_75t_L g6364 ( 
.A(n_6224),
.Y(n_6364)
);

INVxp67_ASAP7_75t_L g6365 ( 
.A(n_6174),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6250),
.Y(n_6366)
);

NAND2x1p5_ASAP7_75t_L g6367 ( 
.A(n_6166),
.B(n_5933),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_6223),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_6224),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6210),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_6112),
.B(n_5930),
.Y(n_6371)
);

BUFx3_ASAP7_75t_L g6372 ( 
.A(n_6244),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6211),
.Y(n_6373)
);

INVx2_ASAP7_75t_L g6374 ( 
.A(n_6131),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_6212),
.Y(n_6375)
);

INVx3_ASAP7_75t_L g6376 ( 
.A(n_6196),
.Y(n_6376)
);

INVx2_ASAP7_75t_L g6377 ( 
.A(n_6131),
.Y(n_6377)
);

AND2x2_ASAP7_75t_L g6378 ( 
.A(n_6090),
.B(n_5940),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_6108),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_6139),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_6206),
.Y(n_6381)
);

BUFx12f_ASAP7_75t_L g6382 ( 
.A(n_6226),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6206),
.Y(n_6383)
);

NAND2xp5_ASAP7_75t_L g6384 ( 
.A(n_6232),
.B(n_6050),
.Y(n_6384)
);

INVx2_ASAP7_75t_L g6385 ( 
.A(n_6149),
.Y(n_6385)
);

HB1xp67_ASAP7_75t_L g6386 ( 
.A(n_6104),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6172),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_6167),
.Y(n_6388)
);

INVx4_ASAP7_75t_L g6389 ( 
.A(n_6251),
.Y(n_6389)
);

AND2x4_ASAP7_75t_L g6390 ( 
.A(n_6262),
.B(n_5887),
.Y(n_6390)
);

BUFx2_ASAP7_75t_L g6391 ( 
.A(n_6214),
.Y(n_6391)
);

BUFx6f_ASAP7_75t_L g6392 ( 
.A(n_6261),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6129),
.Y(n_6393)
);

HB1xp67_ASAP7_75t_L g6394 ( 
.A(n_6107),
.Y(n_6394)
);

OAI21x1_ASAP7_75t_SL g6395 ( 
.A1(n_6233),
.A2(n_5885),
.B(n_5944),
.Y(n_6395)
);

BUFx2_ASAP7_75t_L g6396 ( 
.A(n_6248),
.Y(n_6396)
);

OR2x2_ASAP7_75t_L g6397 ( 
.A(n_6082),
.B(n_5895),
.Y(n_6397)
);

BUFx2_ASAP7_75t_L g6398 ( 
.A(n_6168),
.Y(n_6398)
);

NAND2xp5_ASAP7_75t_L g6399 ( 
.A(n_6247),
.B(n_5882),
.Y(n_6399)
);

INVx2_ASAP7_75t_L g6400 ( 
.A(n_6129),
.Y(n_6400)
);

INVx2_ASAP7_75t_L g6401 ( 
.A(n_6235),
.Y(n_6401)
);

INVx2_ASAP7_75t_L g6402 ( 
.A(n_6255),
.Y(n_6402)
);

INVx3_ASAP7_75t_L g6403 ( 
.A(n_6175),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6093),
.Y(n_6404)
);

AOI22xp33_ASAP7_75t_L g6405 ( 
.A1(n_6219),
.A2(n_5864),
.B1(n_5944),
.B2(n_5914),
.Y(n_6405)
);

INVx2_ASAP7_75t_L g6406 ( 
.A(n_6151),
.Y(n_6406)
);

BUFx3_ASAP7_75t_L g6407 ( 
.A(n_6216),
.Y(n_6407)
);

HB1xp67_ASAP7_75t_L g6408 ( 
.A(n_6121),
.Y(n_6408)
);

INVx2_ASAP7_75t_L g6409 ( 
.A(n_6151),
.Y(n_6409)
);

OR2x2_ASAP7_75t_L g6410 ( 
.A(n_6126),
.B(n_5895),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_6091),
.Y(n_6411)
);

BUFx6f_ASAP7_75t_L g6412 ( 
.A(n_6182),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6162),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_L g6414 ( 
.A(n_6098),
.B(n_5895),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6162),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_6256),
.Y(n_6416)
);

AND2x4_ASAP7_75t_L g6417 ( 
.A(n_6069),
.B(n_5949),
.Y(n_6417)
);

HB1xp67_ASAP7_75t_L g6418 ( 
.A(n_6138),
.Y(n_6418)
);

INVx2_ASAP7_75t_SL g6419 ( 
.A(n_6202),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_6258),
.Y(n_6420)
);

INVxp67_ASAP7_75t_L g6421 ( 
.A(n_6195),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6254),
.Y(n_6422)
);

BUFx12f_ASAP7_75t_L g6423 ( 
.A(n_6245),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6237),
.Y(n_6424)
);

OAI21xp5_ASAP7_75t_L g6425 ( 
.A1(n_6222),
.A2(n_5982),
.B(n_5975),
.Y(n_6425)
);

NAND2xp5_ASAP7_75t_L g6426 ( 
.A(n_6181),
.B(n_5922),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_6263),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6203),
.Y(n_6428)
);

INVx3_ASAP7_75t_L g6429 ( 
.A(n_6175),
.Y(n_6429)
);

INVxp67_ASAP7_75t_SL g6430 ( 
.A(n_6197),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6136),
.Y(n_6431)
);

OA21x2_ASAP7_75t_L g6432 ( 
.A1(n_6102),
.A2(n_6057),
.B(n_5913),
.Y(n_6432)
);

INVx2_ASAP7_75t_L g6433 ( 
.A(n_6135),
.Y(n_6433)
);

INVx2_ASAP7_75t_L g6434 ( 
.A(n_6259),
.Y(n_6434)
);

HB1xp67_ASAP7_75t_L g6435 ( 
.A(n_6117),
.Y(n_6435)
);

INVx2_ASAP7_75t_SL g6436 ( 
.A(n_6202),
.Y(n_6436)
);

OR2x6_ASAP7_75t_L g6437 ( 
.A(n_6086),
.B(n_5982),
.Y(n_6437)
);

BUFx3_ASAP7_75t_L g6438 ( 
.A(n_6240),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6200),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6135),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_6215),
.Y(n_6441)
);

OAI21xp5_ASAP7_75t_L g6442 ( 
.A1(n_6190),
.A2(n_6061),
.B(n_5959),
.Y(n_6442)
);

INVx2_ASAP7_75t_L g6443 ( 
.A(n_6152),
.Y(n_6443)
);

INVx2_ASAP7_75t_L g6444 ( 
.A(n_6158),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6243),
.Y(n_6445)
);

OAI21x1_ASAP7_75t_L g6446 ( 
.A1(n_6071),
.A2(n_5868),
.B(n_5910),
.Y(n_6446)
);

HB1xp67_ASAP7_75t_L g6447 ( 
.A(n_6120),
.Y(n_6447)
);

OAI21x1_ASAP7_75t_L g6448 ( 
.A1(n_6085),
.A2(n_5931),
.B(n_5928),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6225),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6227),
.Y(n_6450)
);

OA21x2_ASAP7_75t_L g6451 ( 
.A1(n_6161),
.A2(n_6016),
.B(n_6012),
.Y(n_6451)
);

OAI22xp5_ASAP7_75t_SL g6452 ( 
.A1(n_6310),
.A2(n_6101),
.B1(n_6110),
.B2(n_6159),
.Y(n_6452)
);

OR2x2_ASAP7_75t_L g6453 ( 
.A(n_6277),
.B(n_6144),
.Y(n_6453)
);

INVx4_ASAP7_75t_L g6454 ( 
.A(n_6331),
.Y(n_6454)
);

OAI22xp5_ASAP7_75t_L g6455 ( 
.A1(n_6310),
.A2(n_6277),
.B1(n_6352),
.B2(n_6274),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_6304),
.B(n_6187),
.Y(n_6456)
);

OAI21x1_ASAP7_75t_L g6457 ( 
.A1(n_6296),
.A2(n_6185),
.B(n_6068),
.Y(n_6457)
);

AOI22xp5_ASAP7_75t_SL g6458 ( 
.A1(n_6359),
.A2(n_6430),
.B1(n_6276),
.B2(n_6274),
.Y(n_6458)
);

AND2x4_ASAP7_75t_L g6459 ( 
.A(n_6328),
.B(n_6191),
.Y(n_6459)
);

OR2x6_ASAP7_75t_L g6460 ( 
.A(n_6292),
.B(n_6246),
.Y(n_6460)
);

OAI22xp5_ASAP7_75t_L g6461 ( 
.A1(n_6352),
.A2(n_6101),
.B1(n_6125),
.B2(n_6106),
.Y(n_6461)
);

O2A1O1Ixp33_ASAP7_75t_SL g6462 ( 
.A1(n_6276),
.A2(n_6178),
.B(n_6241),
.C(n_6238),
.Y(n_6462)
);

INVx2_ASAP7_75t_L g6463 ( 
.A(n_6438),
.Y(n_6463)
);

AND2x2_ASAP7_75t_L g6464 ( 
.A(n_6280),
.B(n_6165),
.Y(n_6464)
);

AND2x4_ASAP7_75t_L g6465 ( 
.A(n_6438),
.B(n_6260),
.Y(n_6465)
);

NOR2xp33_ASAP7_75t_SL g6466 ( 
.A(n_6280),
.B(n_6252),
.Y(n_6466)
);

A2O1A1Ixp33_ASAP7_75t_L g6467 ( 
.A1(n_6359),
.A2(n_6221),
.B(n_6142),
.C(n_6116),
.Y(n_6467)
);

BUFx3_ASAP7_75t_L g6468 ( 
.A(n_6270),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_6321),
.Y(n_6469)
);

INVx1_ASAP7_75t_SL g6470 ( 
.A(n_6382),
.Y(n_6470)
);

AOI221xp5_ASAP7_75t_L g6471 ( 
.A1(n_6408),
.A2(n_6103),
.B1(n_6264),
.B2(n_6087),
.C(n_6257),
.Y(n_6471)
);

AND2x2_ASAP7_75t_L g6472 ( 
.A(n_6407),
.B(n_6165),
.Y(n_6472)
);

OAI22xp5_ASAP7_75t_L g6473 ( 
.A1(n_6410),
.A2(n_6253),
.B1(n_6143),
.B2(n_6229),
.Y(n_6473)
);

OA21x2_ASAP7_75t_L g6474 ( 
.A1(n_6330),
.A2(n_6153),
.B(n_6148),
.Y(n_6474)
);

OR2x2_ASAP7_75t_L g6475 ( 
.A(n_6271),
.B(n_6217),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_6327),
.Y(n_6476)
);

AOI221xp5_ASAP7_75t_L g6477 ( 
.A1(n_6408),
.A2(n_6217),
.B1(n_6218),
.B2(n_6114),
.C(n_6228),
.Y(n_6477)
);

OR2x2_ASAP7_75t_L g6478 ( 
.A(n_6266),
.B(n_5922),
.Y(n_6478)
);

O2A1O1Ixp33_ASAP7_75t_L g6479 ( 
.A1(n_6324),
.A2(n_5914),
.B(n_5948),
.C(n_5936),
.Y(n_6479)
);

AND2x4_ASAP7_75t_L g6480 ( 
.A(n_6292),
.B(n_6049),
.Y(n_6480)
);

CKINVDCx6p67_ASAP7_75t_R g6481 ( 
.A(n_6372),
.Y(n_6481)
);

OA21x2_ASAP7_75t_L g6482 ( 
.A1(n_6330),
.A2(n_6000),
.B(n_5966),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6284),
.B(n_5956),
.Y(n_6483)
);

NAND2xp5_ASAP7_75t_L g6484 ( 
.A(n_6424),
.B(n_5957),
.Y(n_6484)
);

AND2x2_ASAP7_75t_L g6485 ( 
.A(n_6269),
.B(n_6053),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_6305),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_L g6487 ( 
.A(n_6445),
.B(n_5978),
.Y(n_6487)
);

AOI22xp5_ASAP7_75t_L g6488 ( 
.A1(n_6324),
.A2(n_5968),
.B1(n_5963),
.B2(n_5991),
.Y(n_6488)
);

AND2x4_ASAP7_75t_L g6489 ( 
.A(n_6292),
.B(n_5984),
.Y(n_6489)
);

AOI21xp5_ASAP7_75t_L g6490 ( 
.A1(n_6414),
.A2(n_6011),
.B(n_6014),
.Y(n_6490)
);

OR2x2_ASAP7_75t_L g6491 ( 
.A(n_6428),
.B(n_230),
.Y(n_6491)
);

AND2x4_ASAP7_75t_L g6492 ( 
.A(n_6292),
.B(n_231),
.Y(n_6492)
);

OAI22xp5_ASAP7_75t_L g6493 ( 
.A1(n_6371),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_6493)
);

AND2x2_ASAP7_75t_L g6494 ( 
.A(n_6293),
.B(n_236),
.Y(n_6494)
);

OAI22xp5_ASAP7_75t_L g6495 ( 
.A1(n_6371),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_6495)
);

OA21x2_ASAP7_75t_L g6496 ( 
.A1(n_6341),
.A2(n_6291),
.B(n_6290),
.Y(n_6496)
);

AO32x2_ASAP7_75t_L g6497 ( 
.A1(n_6419),
.A2(n_6436),
.A3(n_6389),
.B1(n_6333),
.B2(n_6418),
.Y(n_6497)
);

INVx2_ASAP7_75t_L g6498 ( 
.A(n_6306),
.Y(n_6498)
);

OAI21x1_ASAP7_75t_SL g6499 ( 
.A1(n_6354),
.A2(n_243),
.B(n_245),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6305),
.Y(n_6500)
);

OAI21xp5_ASAP7_75t_L g6501 ( 
.A1(n_6426),
.A2(n_6365),
.B(n_6351),
.Y(n_6501)
);

OR2x2_ASAP7_75t_L g6502 ( 
.A(n_6308),
.B(n_243),
.Y(n_6502)
);

OAI22xp5_ASAP7_75t_SL g6503 ( 
.A1(n_6275),
.A2(n_6404),
.B1(n_6286),
.B2(n_6423),
.Y(n_6503)
);

AND2x4_ASAP7_75t_L g6504 ( 
.A(n_6306),
.B(n_245),
.Y(n_6504)
);

OR2x2_ASAP7_75t_L g6505 ( 
.A(n_6353),
.B(n_6329),
.Y(n_6505)
);

AND2x2_ASAP7_75t_L g6506 ( 
.A(n_6391),
.B(n_6286),
.Y(n_6506)
);

AND2x4_ASAP7_75t_L g6507 ( 
.A(n_6306),
.B(n_246),
.Y(n_6507)
);

OR2x2_ASAP7_75t_L g6508 ( 
.A(n_6353),
.B(n_247),
.Y(n_6508)
);

AOI21xp33_ASAP7_75t_L g6509 ( 
.A1(n_6426),
.A2(n_247),
.B(n_248),
.Y(n_6509)
);

OR2x6_ASAP7_75t_L g6510 ( 
.A(n_6306),
.B(n_1518),
.Y(n_6510)
);

HB1xp67_ASAP7_75t_L g6511 ( 
.A(n_6268),
.Y(n_6511)
);

OAI21x1_ASAP7_75t_SL g6512 ( 
.A1(n_6318),
.A2(n_249),
.B(n_250),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_6367),
.Y(n_6513)
);

AOI221xp5_ASAP7_75t_L g6514 ( 
.A1(n_6418),
.A2(n_2243),
.B1(n_2262),
.B2(n_2259),
.C(n_2258),
.Y(n_6514)
);

OAI21xp5_ASAP7_75t_L g6515 ( 
.A1(n_6365),
.A2(n_6351),
.B(n_6425),
.Y(n_6515)
);

AOI31xp33_ASAP7_75t_SL g6516 ( 
.A1(n_6421),
.A2(n_254),
.A3(n_251),
.B(n_252),
.Y(n_6516)
);

OAI21x1_ASAP7_75t_L g6517 ( 
.A1(n_6279),
.A2(n_2171),
.B(n_2165),
.Y(n_6517)
);

NOR2x1_ASAP7_75t_SL g6518 ( 
.A(n_6437),
.B(n_252),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_6367),
.Y(n_6519)
);

NAND2xp5_ASAP7_75t_L g6520 ( 
.A(n_6416),
.B(n_254),
.Y(n_6520)
);

OR2x2_ASAP7_75t_L g6521 ( 
.A(n_6360),
.B(n_255),
.Y(n_6521)
);

HB1xp67_ASAP7_75t_L g6522 ( 
.A(n_6325),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_6412),
.Y(n_6523)
);

AND2x4_ASAP7_75t_SL g6524 ( 
.A(n_6389),
.B(n_255),
.Y(n_6524)
);

A2O1A1Ixp33_ASAP7_75t_L g6525 ( 
.A1(n_6309),
.A2(n_260),
.B(n_256),
.C(n_259),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_6339),
.Y(n_6526)
);

INVx3_ASAP7_75t_L g6527 ( 
.A(n_6372),
.Y(n_6527)
);

AO32x1_ASAP7_75t_L g6528 ( 
.A1(n_6333),
.A2(n_262),
.A3(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6398),
.B(n_263),
.Y(n_6529)
);

OR2x6_ASAP7_75t_L g6530 ( 
.A(n_6275),
.B(n_1518),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6344),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6345),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6348),
.Y(n_6533)
);

NAND2x1p5_ASAP7_75t_L g6534 ( 
.A(n_6300),
.B(n_1518),
.Y(n_6534)
);

A2O1A1Ixp33_ASAP7_75t_L g6535 ( 
.A1(n_6309),
.A2(n_267),
.B(n_264),
.C(n_266),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_6412),
.Y(n_6536)
);

AND2x2_ASAP7_75t_L g6537 ( 
.A(n_6343),
.B(n_268),
.Y(n_6537)
);

O2A1O1Ixp33_ASAP7_75t_L g6538 ( 
.A1(n_6320),
.A2(n_272),
.B(n_269),
.C(n_271),
.Y(n_6538)
);

OR2x2_ASAP7_75t_L g6539 ( 
.A(n_6285),
.B(n_272),
.Y(n_6539)
);

BUFx6f_ASAP7_75t_L g6540 ( 
.A(n_6392),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_L g6541 ( 
.A(n_6420),
.B(n_273),
.Y(n_6541)
);

INVx2_ASAP7_75t_L g6542 ( 
.A(n_6412),
.Y(n_6542)
);

A2O1A1Ixp33_ASAP7_75t_L g6543 ( 
.A1(n_6311),
.A2(n_276),
.B(n_273),
.C(n_275),
.Y(n_6543)
);

AOI22xp5_ASAP7_75t_L g6544 ( 
.A1(n_6291),
.A2(n_2258),
.B1(n_2259),
.B2(n_2243),
.Y(n_6544)
);

NAND2xp5_ASAP7_75t_L g6545 ( 
.A(n_6449),
.B(n_6450),
.Y(n_6545)
);

OR2x2_ASAP7_75t_L g6546 ( 
.A(n_6287),
.B(n_6267),
.Y(n_6546)
);

HB1xp67_ASAP7_75t_L g6547 ( 
.A(n_6325),
.Y(n_6547)
);

AND2x6_ASAP7_75t_L g6548 ( 
.A(n_6392),
.B(n_275),
.Y(n_6548)
);

OAI21xp5_ASAP7_75t_L g6549 ( 
.A1(n_6425),
.A2(n_6311),
.B(n_6341),
.Y(n_6549)
);

AND2x4_ASAP7_75t_L g6550 ( 
.A(n_6441),
.B(n_276),
.Y(n_6550)
);

OA21x2_ASAP7_75t_L g6551 ( 
.A1(n_6434),
.A2(n_277),
.B(n_279),
.Y(n_6551)
);

OAI22xp5_ASAP7_75t_L g6552 ( 
.A1(n_6396),
.A2(n_6294),
.B1(n_6405),
.B2(n_6437),
.Y(n_6552)
);

AND2x6_ASAP7_75t_L g6553 ( 
.A(n_6392),
.B(n_282),
.Y(n_6553)
);

INVx1_ASAP7_75t_SL g6554 ( 
.A(n_6392),
.Y(n_6554)
);

AOI21xp5_ASAP7_75t_L g6555 ( 
.A1(n_6350),
.A2(n_283),
.B(n_284),
.Y(n_6555)
);

NAND2xp5_ASAP7_75t_L g6556 ( 
.A(n_6307),
.B(n_285),
.Y(n_6556)
);

BUFx3_ASAP7_75t_L g6557 ( 
.A(n_6332),
.Y(n_6557)
);

INVx2_ASAP7_75t_L g6558 ( 
.A(n_6315),
.Y(n_6558)
);

AO22x2_ASAP7_75t_L g6559 ( 
.A1(n_6295),
.A2(n_6302),
.B1(n_6303),
.B2(n_6298),
.Y(n_6559)
);

INVx3_ASAP7_75t_L g6560 ( 
.A(n_6313),
.Y(n_6560)
);

AND2x6_ASAP7_75t_L g6561 ( 
.A(n_6315),
.B(n_287),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6370),
.Y(n_6562)
);

AND2x2_ASAP7_75t_L g6563 ( 
.A(n_6358),
.B(n_288),
.Y(n_6563)
);

AOI21xp5_ASAP7_75t_L g6564 ( 
.A1(n_6350),
.A2(n_289),
.B(n_291),
.Y(n_6564)
);

AND2x2_ASAP7_75t_L g6565 ( 
.A(n_6361),
.B(n_289),
.Y(n_6565)
);

AND2x2_ASAP7_75t_L g6566 ( 
.A(n_6362),
.B(n_291),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_6307),
.B(n_292),
.Y(n_6567)
);

INVx1_ASAP7_75t_L g6568 ( 
.A(n_6373),
.Y(n_6568)
);

AO32x2_ASAP7_75t_L g6569 ( 
.A1(n_6313),
.A2(n_295),
.A3(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_6569)
);

AND2x4_ASAP7_75t_L g6570 ( 
.A(n_6439),
.B(n_298),
.Y(n_6570)
);

A2O1A1Ixp33_ASAP7_75t_L g6571 ( 
.A1(n_6366),
.A2(n_301),
.B(n_299),
.C(n_300),
.Y(n_6571)
);

INVx3_ASAP7_75t_L g6572 ( 
.A(n_6314),
.Y(n_6572)
);

NOR2xp33_ASAP7_75t_L g6573 ( 
.A(n_6314),
.B(n_300),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_6369),
.B(n_6431),
.Y(n_6574)
);

AO32x2_ASAP7_75t_L g6575 ( 
.A1(n_6363),
.A2(n_304),
.A3(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_6575)
);

BUFx3_ASAP7_75t_L g6576 ( 
.A(n_6326),
.Y(n_6576)
);

INVx2_ASAP7_75t_L g6577 ( 
.A(n_6295),
.Y(n_6577)
);

A2O1A1Ixp33_ASAP7_75t_L g6578 ( 
.A1(n_6405),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_6578)
);

NAND2xp5_ASAP7_75t_L g6579 ( 
.A(n_6422),
.B(n_308),
.Y(n_6579)
);

AO32x2_ASAP7_75t_L g6580 ( 
.A1(n_6411),
.A2(n_312),
.A3(n_310),
.B1(n_311),
.B2(n_313),
.Y(n_6580)
);

AND2x2_ASAP7_75t_L g6581 ( 
.A(n_6378),
.B(n_310),
.Y(n_6581)
);

O2A1O1Ixp33_ASAP7_75t_L g6582 ( 
.A1(n_6342),
.A2(n_316),
.B(n_311),
.C(n_315),
.Y(n_6582)
);

AO22x2_ASAP7_75t_L g6583 ( 
.A1(n_6302),
.A2(n_6303),
.B1(n_6273),
.B2(n_6278),
.Y(n_6583)
);

INVx2_ASAP7_75t_L g6584 ( 
.A(n_6335),
.Y(n_6584)
);

INVx2_ASAP7_75t_L g6585 ( 
.A(n_6335),
.Y(n_6585)
);

OR2x6_ASAP7_75t_L g6586 ( 
.A(n_6338),
.B(n_1518),
.Y(n_6586)
);

OAI21xp5_ASAP7_75t_L g6587 ( 
.A1(n_6442),
.A2(n_317),
.B(n_320),
.Y(n_6587)
);

INVx2_ASAP7_75t_L g6588 ( 
.A(n_6468),
.Y(n_6588)
);

OR2x2_ASAP7_75t_L g6589 ( 
.A(n_6505),
.B(n_6545),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6540),
.Y(n_6590)
);

OAI221xp5_ASAP7_75t_L g6591 ( 
.A1(n_6467),
.A2(n_6383),
.B1(n_6381),
.B2(n_6379),
.C(n_6399),
.Y(n_6591)
);

INVxp67_ASAP7_75t_L g6592 ( 
.A(n_6548),
.Y(n_6592)
);

OR2x2_ASAP7_75t_L g6593 ( 
.A(n_6508),
.B(n_6475),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6559),
.Y(n_6594)
);

AND2x4_ASAP7_75t_L g6595 ( 
.A(n_6576),
.B(n_6281),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_6540),
.Y(n_6596)
);

O2A1O1Ixp5_ASAP7_75t_L g6597 ( 
.A1(n_6455),
.A2(n_6400),
.B(n_6393),
.C(n_6433),
.Y(n_6597)
);

INVx2_ASAP7_75t_L g6598 ( 
.A(n_6527),
.Y(n_6598)
);

INVx2_ASAP7_75t_L g6599 ( 
.A(n_6456),
.Y(n_6599)
);

AOI22xp33_ASAP7_75t_L g6600 ( 
.A1(n_6477),
.A2(n_6342),
.B1(n_6400),
.B2(n_6393),
.Y(n_6600)
);

INVx1_ASAP7_75t_L g6601 ( 
.A(n_6559),
.Y(n_6601)
);

OR2x2_ASAP7_75t_L g6602 ( 
.A(n_6511),
.B(n_6282),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6583),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_6583),
.Y(n_6604)
);

INVx1_ASAP7_75t_L g6605 ( 
.A(n_6496),
.Y(n_6605)
);

AND2x4_ASAP7_75t_L g6606 ( 
.A(n_6459),
.B(n_6338),
.Y(n_6606)
);

BUFx3_ASAP7_75t_L g6607 ( 
.A(n_6481),
.Y(n_6607)
);

NAND2xp5_ASAP7_75t_L g6608 ( 
.A(n_6496),
.B(n_6288),
.Y(n_6608)
);

INVx2_ASAP7_75t_L g6609 ( 
.A(n_6518),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_L g6610 ( 
.A(n_6555),
.B(n_6564),
.Y(n_6610)
);

BUFx2_ASAP7_75t_L g6611 ( 
.A(n_6497),
.Y(n_6611)
);

AND2x4_ASAP7_75t_SL g6612 ( 
.A(n_6454),
.B(n_6364),
.Y(n_6612)
);

AND2x2_ASAP7_75t_L g6613 ( 
.A(n_6470),
.B(n_6364),
.Y(n_6613)
);

AOI22xp33_ASAP7_75t_L g6614 ( 
.A1(n_6466),
.A2(n_6409),
.B1(n_6406),
.B2(n_6413),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6577),
.Y(n_6615)
);

INVxp67_ASAP7_75t_SL g6616 ( 
.A(n_6458),
.Y(n_6616)
);

INVx3_ASAP7_75t_SL g6617 ( 
.A(n_6492),
.Y(n_6617)
);

AO21x2_ASAP7_75t_L g6618 ( 
.A1(n_6556),
.A2(n_6319),
.B(n_6317),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_6506),
.B(n_6340),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6522),
.Y(n_6620)
);

OAI221xp5_ASAP7_75t_L g6621 ( 
.A1(n_6501),
.A2(n_6379),
.B1(n_6399),
.B2(n_6394),
.C(n_6442),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6547),
.Y(n_6622)
);

AND2x2_ASAP7_75t_L g6623 ( 
.A(n_6464),
.B(n_6356),
.Y(n_6623)
);

AND2x2_ASAP7_75t_L g6624 ( 
.A(n_6472),
.B(n_6403),
.Y(n_6624)
);

INVxp67_ASAP7_75t_L g6625 ( 
.A(n_6548),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6463),
.B(n_6403),
.Y(n_6626)
);

AND2x4_ASAP7_75t_L g6627 ( 
.A(n_6498),
.B(n_6429),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6567),
.Y(n_6628)
);

INVx2_ASAP7_75t_L g6629 ( 
.A(n_6569),
.Y(n_6629)
);

AND2x2_ASAP7_75t_L g6630 ( 
.A(n_6529),
.B(n_6376),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6486),
.Y(n_6631)
);

AND2x2_ASAP7_75t_L g6632 ( 
.A(n_6574),
.B(n_6334),
.Y(n_6632)
);

OR2x2_ASAP7_75t_L g6633 ( 
.A(n_6546),
.B(n_6491),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6500),
.Y(n_6634)
);

NAND2x1_ASAP7_75t_L g6635 ( 
.A(n_6499),
.B(n_6443),
.Y(n_6635)
);

INVxp33_ASAP7_75t_L g6636 ( 
.A(n_6499),
.Y(n_6636)
);

AND2x2_ASAP7_75t_L g6637 ( 
.A(n_6494),
.B(n_6581),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6582),
.B(n_6289),
.Y(n_6638)
);

NAND2xp5_ASAP7_75t_L g6639 ( 
.A(n_6578),
.B(n_6297),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6575),
.Y(n_6640)
);

OR2x2_ASAP7_75t_L g6641 ( 
.A(n_6502),
.B(n_6349),
.Y(n_6641)
);

BUFx2_ASAP7_75t_L g6642 ( 
.A(n_6497),
.Y(n_6642)
);

NAND2xp5_ASAP7_75t_SL g6643 ( 
.A(n_6461),
.B(n_6337),
.Y(n_6643)
);

HB1xp67_ASAP7_75t_L g6644 ( 
.A(n_6549),
.Y(n_6644)
);

NAND2xp5_ASAP7_75t_L g6645 ( 
.A(n_6509),
.B(n_6561),
.Y(n_6645)
);

AO21x2_ASAP7_75t_L g6646 ( 
.A1(n_6515),
.A2(n_6319),
.B(n_6317),
.Y(n_6646)
);

OR2x2_ASAP7_75t_L g6647 ( 
.A(n_6554),
.B(n_6299),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_6569),
.Y(n_6648)
);

INVx3_ASAP7_75t_L g6649 ( 
.A(n_6572),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6561),
.B(n_6312),
.Y(n_6650)
);

INVx2_ASAP7_75t_SL g6651 ( 
.A(n_6524),
.Y(n_6651)
);

INVx2_ASAP7_75t_SL g6652 ( 
.A(n_6504),
.Y(n_6652)
);

INVx2_ASAP7_75t_L g6653 ( 
.A(n_6510),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6520),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6541),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_6469),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6561),
.B(n_6316),
.Y(n_6657)
);

INVx3_ASAP7_75t_L g6658 ( 
.A(n_6465),
.Y(n_6658)
);

HB1xp67_ASAP7_75t_L g6659 ( 
.A(n_6551),
.Y(n_6659)
);

BUFx6f_ASAP7_75t_SL g6660 ( 
.A(n_6507),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6476),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_L g6662 ( 
.A(n_6548),
.B(n_6323),
.Y(n_6662)
);

OAI22xp5_ASAP7_75t_SL g6663 ( 
.A1(n_6503),
.A2(n_6433),
.B1(n_6337),
.B2(n_6440),
.Y(n_6663)
);

HB1xp67_ASAP7_75t_L g6664 ( 
.A(n_6551),
.Y(n_6664)
);

CKINVDCx5p33_ASAP7_75t_R g6665 ( 
.A(n_6553),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_6510),
.Y(n_6666)
);

INVx3_ASAP7_75t_L g6667 ( 
.A(n_6560),
.Y(n_6667)
);

OR2x2_ASAP7_75t_L g6668 ( 
.A(n_6579),
.B(n_6368),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6460),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6580),
.Y(n_6670)
);

BUFx3_ASAP7_75t_L g6671 ( 
.A(n_6550),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6526),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6534),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6531),
.Y(n_6674)
);

INVx2_ASAP7_75t_L g6675 ( 
.A(n_6557),
.Y(n_6675)
);

INVx2_ASAP7_75t_L g6676 ( 
.A(n_6586),
.Y(n_6676)
);

AND2x4_ASAP7_75t_L g6677 ( 
.A(n_6523),
.B(n_6444),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6532),
.Y(n_6678)
);

INVx2_ASAP7_75t_SL g6679 ( 
.A(n_6537),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6533),
.Y(n_6680)
);

AND2x4_ASAP7_75t_L g6681 ( 
.A(n_6536),
.B(n_6336),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6562),
.Y(n_6682)
);

AND2x4_ASAP7_75t_L g6683 ( 
.A(n_6542),
.B(n_6417),
.Y(n_6683)
);

AOI221xp5_ASAP7_75t_L g6684 ( 
.A1(n_6479),
.A2(n_6386),
.B1(n_6394),
.B2(n_6447),
.C(n_6435),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6473),
.B(n_6375),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6584),
.B(n_6448),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6568),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_6539),
.Y(n_6688)
);

AOI21xp5_ASAP7_75t_SL g6689 ( 
.A1(n_6587),
.A2(n_6535),
.B(n_6525),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6487),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6484),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6521),
.Y(n_6692)
);

AND2x2_ASAP7_75t_L g6693 ( 
.A(n_6585),
.B(n_6417),
.Y(n_6693)
);

OA21x2_ASAP7_75t_L g6694 ( 
.A1(n_6597),
.A2(n_6471),
.B(n_6457),
.Y(n_6694)
);

NAND2xp5_ASAP7_75t_SL g6695 ( 
.A(n_6637),
.B(n_6452),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_L g6696 ( 
.A(n_6679),
.B(n_6573),
.Y(n_6696)
);

NAND3xp33_ASAP7_75t_L g6697 ( 
.A(n_6616),
.B(n_6597),
.C(n_6644),
.Y(n_6697)
);

NAND3xp33_ASAP7_75t_L g6698 ( 
.A(n_6616),
.B(n_6644),
.C(n_6642),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_6652),
.B(n_6453),
.Y(n_6699)
);

AOI221xp5_ASAP7_75t_L g6700 ( 
.A1(n_6614),
.A2(n_6591),
.B1(n_6621),
.B2(n_6684),
.C(n_6600),
.Y(n_6700)
);

NAND3xp33_ASAP7_75t_L g6701 ( 
.A(n_6611),
.B(n_6495),
.C(n_6493),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6607),
.B(n_6483),
.Y(n_6702)
);

AND2x2_ASAP7_75t_L g6703 ( 
.A(n_6623),
.B(n_6485),
.Y(n_6703)
);

AND2x2_ASAP7_75t_L g6704 ( 
.A(n_6619),
.B(n_6630),
.Y(n_6704)
);

AOI22xp33_ASAP7_75t_L g6705 ( 
.A1(n_6670),
.A2(n_6415),
.B1(n_6413),
.B2(n_6409),
.Y(n_6705)
);

NAND2xp5_ASAP7_75t_SL g6706 ( 
.A(n_6609),
.B(n_6606),
.Y(n_6706)
);

NAND2xp5_ASAP7_75t_L g6707 ( 
.A(n_6692),
.B(n_6462),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6613),
.B(n_6563),
.Y(n_6708)
);

NAND2xp5_ASAP7_75t_L g6709 ( 
.A(n_6688),
.B(n_6570),
.Y(n_6709)
);

AOI211xp5_ASAP7_75t_L g6710 ( 
.A1(n_6591),
.A2(n_6516),
.B(n_6552),
.C(n_6538),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6612),
.B(n_6565),
.Y(n_6711)
);

AOI22xp33_ASAP7_75t_L g6712 ( 
.A1(n_6629),
.A2(n_6415),
.B1(n_6406),
.B2(n_6377),
.Y(n_6712)
);

OAI22xp5_ASAP7_75t_L g6713 ( 
.A1(n_6600),
.A2(n_6543),
.B1(n_6558),
.B2(n_6397),
.Y(n_6713)
);

OAI221xp5_ASAP7_75t_L g6714 ( 
.A1(n_6614),
.A2(n_6621),
.B1(n_6684),
.B2(n_6610),
.C(n_6604),
.Y(n_6714)
);

AOI21xp33_ASAP7_75t_L g6715 ( 
.A1(n_6636),
.A2(n_6519),
.B(n_6513),
.Y(n_6715)
);

AND2x2_ASAP7_75t_L g6716 ( 
.A(n_6624),
.B(n_6566),
.Y(n_6716)
);

NAND2xp5_ASAP7_75t_L g6717 ( 
.A(n_6593),
.B(n_6571),
.Y(n_6717)
);

AND2x2_ASAP7_75t_SL g6718 ( 
.A(n_6589),
.B(n_6480),
.Y(n_6718)
);

NAND2xp5_ASAP7_75t_L g6719 ( 
.A(n_6648),
.B(n_6512),
.Y(n_6719)
);

NAND2xp5_ASAP7_75t_L g6720 ( 
.A(n_6610),
.B(n_6512),
.Y(n_6720)
);

OAI22xp5_ASAP7_75t_L g6721 ( 
.A1(n_6685),
.A2(n_6478),
.B1(n_6530),
.B2(n_6488),
.Y(n_6721)
);

AND2x2_ASAP7_75t_L g6722 ( 
.A(n_6588),
.B(n_6530),
.Y(n_6722)
);

OAI22xp5_ASAP7_75t_L g6723 ( 
.A1(n_6685),
.A2(n_6377),
.B1(n_6374),
.B2(n_6489),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6617),
.B(n_6435),
.Y(n_6724)
);

NOR3xp33_ASAP7_75t_SL g6725 ( 
.A(n_6663),
.B(n_6490),
.C(n_6514),
.Y(n_6725)
);

AOI221xp5_ASAP7_75t_L g6726 ( 
.A1(n_6603),
.A2(n_6447),
.B1(n_6301),
.B2(n_6355),
.C(n_6384),
.Y(n_6726)
);

NAND2xp33_ASAP7_75t_SL g6727 ( 
.A(n_6635),
.B(n_6390),
.Y(n_6727)
);

OAI221xp5_ASAP7_75t_L g6728 ( 
.A1(n_6594),
.A2(n_6387),
.B1(n_6474),
.B2(n_6384),
.C(n_6322),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6601),
.Y(n_6729)
);

NOR3xp33_ASAP7_75t_SL g6730 ( 
.A(n_6663),
.B(n_6355),
.C(n_6528),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_L g6731 ( 
.A(n_6633),
.B(n_6301),
.Y(n_6731)
);

AOI21xp5_ASAP7_75t_SL g6732 ( 
.A1(n_6660),
.A2(n_6651),
.B(n_6665),
.Y(n_6732)
);

OAI21xp33_ASAP7_75t_L g6733 ( 
.A1(n_6675),
.A2(n_6357),
.B(n_6517),
.Y(n_6733)
);

NAND3xp33_ASAP7_75t_L g6734 ( 
.A(n_6592),
.B(n_6544),
.C(n_6474),
.Y(n_6734)
);

AND2x2_ASAP7_75t_SL g6735 ( 
.A(n_6645),
.B(n_6595),
.Y(n_6735)
);

NAND3xp33_ASAP7_75t_L g6736 ( 
.A(n_6625),
.B(n_6385),
.C(n_6380),
.Y(n_6736)
);

AND2x2_ASAP7_75t_L g6737 ( 
.A(n_6599),
.B(n_6446),
.Y(n_6737)
);

NAND3xp33_ASAP7_75t_L g6738 ( 
.A(n_6605),
.B(n_6385),
.C(n_6380),
.Y(n_6738)
);

AOI22xp5_ASAP7_75t_SL g6739 ( 
.A1(n_6639),
.A2(n_6451),
.B1(n_6528),
.B2(n_6482),
.Y(n_6739)
);

AND2x2_ASAP7_75t_L g6740 ( 
.A(n_6626),
.B(n_6451),
.Y(n_6740)
);

OAI21xp5_ASAP7_75t_SL g6741 ( 
.A1(n_6639),
.A2(n_6346),
.B(n_6427),
.Y(n_6741)
);

NAND3xp33_ASAP7_75t_L g6742 ( 
.A(n_6608),
.B(n_6388),
.C(n_6482),
.Y(n_6742)
);

NAND3xp33_ASAP7_75t_L g6743 ( 
.A(n_6608),
.B(n_6388),
.C(n_6432),
.Y(n_6743)
);

NAND2xp5_ASAP7_75t_L g6744 ( 
.A(n_6654),
.B(n_6283),
.Y(n_6744)
);

AOI22xp33_ASAP7_75t_L g6745 ( 
.A1(n_6640),
.A2(n_6347),
.B1(n_6402),
.B2(n_6401),
.Y(n_6745)
);

AND2x2_ASAP7_75t_L g6746 ( 
.A(n_6632),
.B(n_6272),
.Y(n_6746)
);

OAI221xp5_ASAP7_75t_L g6747 ( 
.A1(n_6689),
.A2(n_6401),
.B1(n_6402),
.B2(n_6432),
.C(n_6395),
.Y(n_6747)
);

AOI22xp33_ASAP7_75t_L g6748 ( 
.A1(n_6659),
.A2(n_6347),
.B1(n_2272),
.B2(n_2293),
.Y(n_6748)
);

OA21x2_ASAP7_75t_L g6749 ( 
.A1(n_6664),
.A2(n_326),
.B(n_327),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6598),
.B(n_326),
.Y(n_6750)
);

NAND2xp5_ASAP7_75t_L g6751 ( 
.A(n_6655),
.B(n_328),
.Y(n_6751)
);

NAND4xp25_ASAP7_75t_L g6752 ( 
.A(n_6658),
.B(n_333),
.C(n_330),
.D(n_331),
.Y(n_6752)
);

NAND2xp5_ASAP7_75t_L g6753 ( 
.A(n_6628),
.B(n_331),
.Y(n_6753)
);

OAI22xp5_ASAP7_75t_L g6754 ( 
.A1(n_6638),
.A2(n_336),
.B1(n_333),
.B2(n_334),
.Y(n_6754)
);

NAND3xp33_ASAP7_75t_L g6755 ( 
.A(n_6620),
.B(n_6622),
.C(n_6615),
.Y(n_6755)
);

NAND2xp5_ASAP7_75t_L g6756 ( 
.A(n_6671),
.B(n_336),
.Y(n_6756)
);

AND2x2_ASAP7_75t_L g6757 ( 
.A(n_6649),
.B(n_337),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6693),
.B(n_337),
.Y(n_6758)
);

AOI211xp5_ASAP7_75t_L g6759 ( 
.A1(n_6643),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_6759)
);

AOI22xp33_ASAP7_75t_L g6760 ( 
.A1(n_6618),
.A2(n_2272),
.B1(n_2293),
.B2(n_2263),
.Y(n_6760)
);

AND2x2_ASAP7_75t_L g6761 ( 
.A(n_6590),
.B(n_343),
.Y(n_6761)
);

OAI22xp5_ASAP7_75t_L g6762 ( 
.A1(n_6602),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_6596),
.B(n_346),
.Y(n_6763)
);

NAND3xp33_ASAP7_75t_L g6764 ( 
.A(n_6631),
.B(n_347),
.C(n_348),
.Y(n_6764)
);

NAND4xp25_ASAP7_75t_L g6765 ( 
.A(n_6667),
.B(n_354),
.C(n_350),
.D(n_352),
.Y(n_6765)
);

NAND3xp33_ASAP7_75t_L g6766 ( 
.A(n_6634),
.B(n_354),
.C(n_355),
.Y(n_6766)
);

AND2x2_ASAP7_75t_L g6767 ( 
.A(n_6627),
.B(n_357),
.Y(n_6767)
);

OAI22xp5_ASAP7_75t_L g6768 ( 
.A1(n_6641),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_6768)
);

NAND3xp33_ASAP7_75t_L g6769 ( 
.A(n_6662),
.B(n_360),
.C(n_361),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6627),
.B(n_361),
.Y(n_6770)
);

OAI21xp5_ASAP7_75t_SL g6771 ( 
.A1(n_6662),
.A2(n_363),
.B(n_365),
.Y(n_6771)
);

AOI22xp33_ASAP7_75t_L g6772 ( 
.A1(n_6618),
.A2(n_2272),
.B1(n_2293),
.B2(n_2263),
.Y(n_6772)
);

NAND4xp25_ASAP7_75t_L g6773 ( 
.A(n_6647),
.B(n_367),
.C(n_365),
.D(n_366),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_L g6774 ( 
.A(n_6677),
.B(n_368),
.Y(n_6774)
);

OAI22xp5_ASAP7_75t_L g6775 ( 
.A1(n_6650),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_6775)
);

NAND3xp33_ASAP7_75t_L g6776 ( 
.A(n_6669),
.B(n_2239),
.C(n_2232),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6683),
.B(n_370),
.Y(n_6777)
);

NAND4xp25_ASAP7_75t_L g6778 ( 
.A(n_6686),
.B(n_376),
.C(n_371),
.D(n_373),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6683),
.B(n_6681),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6690),
.B(n_376),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6691),
.B(n_378),
.Y(n_6781)
);

NAND4xp25_ASAP7_75t_L g6782 ( 
.A(n_6672),
.B(n_381),
.C(n_379),
.D(n_380),
.Y(n_6782)
);

AND2x2_ASAP7_75t_SL g6783 ( 
.A(n_6668),
.B(n_380),
.Y(n_6783)
);

AOI22xp33_ASAP7_75t_L g6784 ( 
.A1(n_6646),
.A2(n_2293),
.B1(n_2239),
.B2(n_2232),
.Y(n_6784)
);

INVx1_ASAP7_75t_SL g6785 ( 
.A(n_6735),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6749),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_6749),
.Y(n_6787)
);

OR2x2_ASAP7_75t_L g6788 ( 
.A(n_6697),
.B(n_6657),
.Y(n_6788)
);

HB1xp67_ASAP7_75t_L g6789 ( 
.A(n_6697),
.Y(n_6789)
);

NAND2x1_ASAP7_75t_L g6790 ( 
.A(n_6732),
.B(n_6674),
.Y(n_6790)
);

AND2x4_ASAP7_75t_L g6791 ( 
.A(n_6779),
.B(n_6711),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6704),
.B(n_6678),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6780),
.Y(n_6793)
);

AND2x2_ASAP7_75t_SL g6794 ( 
.A(n_6700),
.B(n_6680),
.Y(n_6794)
);

OR2x2_ASAP7_75t_L g6795 ( 
.A(n_6698),
.B(n_6682),
.Y(n_6795)
);

INVx3_ASAP7_75t_L g6796 ( 
.A(n_6708),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_6781),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6729),
.Y(n_6798)
);

INVxp67_ASAP7_75t_L g6799 ( 
.A(n_6698),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6719),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_6694),
.Y(n_6801)
);

AND2x4_ASAP7_75t_L g6802 ( 
.A(n_6716),
.B(n_6687),
.Y(n_6802)
);

AND2x2_ASAP7_75t_L g6803 ( 
.A(n_6702),
.B(n_6673),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6694),
.Y(n_6804)
);

INVx1_ASAP7_75t_L g6805 ( 
.A(n_6738),
.Y(n_6805)
);

INVx2_ASAP7_75t_L g6806 ( 
.A(n_6783),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6758),
.Y(n_6807)
);

INVx3_ASAP7_75t_L g6808 ( 
.A(n_6777),
.Y(n_6808)
);

INVx2_ASAP7_75t_L g6809 ( 
.A(n_6767),
.Y(n_6809)
);

INVx2_ASAP7_75t_L g6810 ( 
.A(n_6770),
.Y(n_6810)
);

AND2x2_ASAP7_75t_L g6811 ( 
.A(n_6703),
.B(n_6656),
.Y(n_6811)
);

AND2x4_ASAP7_75t_L g6812 ( 
.A(n_6706),
.B(n_6661),
.Y(n_6812)
);

HB1xp67_ASAP7_75t_L g6813 ( 
.A(n_6714),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6738),
.Y(n_6814)
);

AND2x4_ASAP7_75t_L g6815 ( 
.A(n_6750),
.B(n_6676),
.Y(n_6815)
);

INVx2_ASAP7_75t_L g6816 ( 
.A(n_6757),
.Y(n_6816)
);

BUFx2_ASAP7_75t_SL g6817 ( 
.A(n_6761),
.Y(n_6817)
);

AND2x4_ASAP7_75t_L g6818 ( 
.A(n_6722),
.B(n_6653),
.Y(n_6818)
);

AND2x4_ASAP7_75t_SL g6819 ( 
.A(n_6763),
.B(n_6666),
.Y(n_6819)
);

HB1xp67_ASAP7_75t_L g6820 ( 
.A(n_6769),
.Y(n_6820)
);

INVx2_ASAP7_75t_L g6821 ( 
.A(n_6718),
.Y(n_6821)
);

NOR2xp33_ASAP7_75t_L g6822 ( 
.A(n_6695),
.B(n_382),
.Y(n_6822)
);

INVxp67_ASAP7_75t_SL g6823 ( 
.A(n_6769),
.Y(n_6823)
);

NAND2xp5_ASAP7_75t_L g6824 ( 
.A(n_6730),
.B(n_6710),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_6774),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6753),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_6756),
.Y(n_6827)
);

AND2x4_ASAP7_75t_L g6828 ( 
.A(n_6724),
.B(n_383),
.Y(n_6828)
);

INVx3_ASAP7_75t_L g6829 ( 
.A(n_6737),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_6710),
.B(n_386),
.Y(n_6830)
);

AND2x2_ASAP7_75t_L g6831 ( 
.A(n_6720),
.B(n_386),
.Y(n_6831)
);

INVx2_ASAP7_75t_L g6832 ( 
.A(n_6699),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_6751),
.Y(n_6833)
);

NAND2xp5_ASAP7_75t_L g6834 ( 
.A(n_6764),
.B(n_390),
.Y(n_6834)
);

NAND2xp5_ASAP7_75t_L g6835 ( 
.A(n_6764),
.B(n_391),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_6766),
.B(n_391),
.Y(n_6836)
);

NAND2xp5_ASAP7_75t_L g6837 ( 
.A(n_6766),
.B(n_393),
.Y(n_6837)
);

AND2x4_ASAP7_75t_L g6838 ( 
.A(n_6709),
.B(n_395),
.Y(n_6838)
);

OR2x2_ASAP7_75t_L g6839 ( 
.A(n_6701),
.B(n_395),
.Y(n_6839)
);

INVx2_ASAP7_75t_L g6840 ( 
.A(n_6707),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6739),
.B(n_396),
.Y(n_6841)
);

INVx3_ASAP7_75t_L g6842 ( 
.A(n_6740),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6715),
.B(n_398),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6736),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_6717),
.Y(n_6845)
);

AND2x4_ASAP7_75t_L g6846 ( 
.A(n_6755),
.B(n_6696),
.Y(n_6846)
);

BUFx2_ASAP7_75t_L g6847 ( 
.A(n_6727),
.Y(n_6847)
);

INVx2_ASAP7_75t_L g6848 ( 
.A(n_6746),
.Y(n_6848)
);

AND2x2_ASAP7_75t_L g6849 ( 
.A(n_6759),
.B(n_401),
.Y(n_6849)
);

INVx3_ASAP7_75t_L g6850 ( 
.A(n_6731),
.Y(n_6850)
);

INVxp67_ASAP7_75t_SL g6851 ( 
.A(n_6759),
.Y(n_6851)
);

AND2x4_ASAP7_75t_L g6852 ( 
.A(n_6705),
.B(n_404),
.Y(n_6852)
);

NAND2x1p5_ASAP7_75t_L g6853 ( 
.A(n_6744),
.B(n_405),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6768),
.Y(n_6854)
);

NAND2xp5_ASAP7_75t_L g6855 ( 
.A(n_6726),
.B(n_406),
.Y(n_6855)
);

NAND2xp5_ASAP7_75t_L g6856 ( 
.A(n_6745),
.B(n_406),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6762),
.Y(n_6857)
);

NOR2xp33_ASAP7_75t_L g6858 ( 
.A(n_6741),
.B(n_407),
.Y(n_6858)
);

BUFx2_ASAP7_75t_L g6859 ( 
.A(n_6773),
.Y(n_6859)
);

INVx1_ASAP7_75t_SL g6860 ( 
.A(n_6789),
.Y(n_6860)
);

OAI21xp5_ASAP7_75t_L g6861 ( 
.A1(n_6789),
.A2(n_6771),
.B(n_6754),
.Y(n_6861)
);

HB1xp67_ASAP7_75t_L g6862 ( 
.A(n_6801),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6786),
.Y(n_6863)
);

OA21x2_ASAP7_75t_L g6864 ( 
.A1(n_6801),
.A2(n_6743),
.B(n_6742),
.Y(n_6864)
);

NAND2x1p5_ASAP7_75t_SL g6865 ( 
.A(n_6804),
.B(n_6712),
.Y(n_6865)
);

NAND3xp33_ASAP7_75t_SL g6866 ( 
.A(n_6804),
.B(n_6747),
.C(n_6713),
.Y(n_6866)
);

INVx1_ASAP7_75t_L g6867 ( 
.A(n_6787),
.Y(n_6867)
);

AND2x4_ASAP7_75t_L g6868 ( 
.A(n_6791),
.B(n_6725),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_6799),
.B(n_6743),
.Y(n_6869)
);

INVxp67_ASAP7_75t_SL g6870 ( 
.A(n_6799),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6796),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6792),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6820),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6807),
.Y(n_6874)
);

OA21x2_ASAP7_75t_L g6875 ( 
.A1(n_6841),
.A2(n_6742),
.B(n_6734),
.Y(n_6875)
);

OAI21x1_ASAP7_75t_L g6876 ( 
.A1(n_6841),
.A2(n_6723),
.B(n_6721),
.Y(n_6876)
);

INVx1_ASAP7_75t_SL g6877 ( 
.A(n_6785),
.Y(n_6877)
);

INVx3_ASAP7_75t_L g6878 ( 
.A(n_6791),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6851),
.Y(n_6879)
);

INVxp67_ASAP7_75t_SL g6880 ( 
.A(n_6788),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6851),
.Y(n_6881)
);

NOR3xp33_ASAP7_75t_SL g6882 ( 
.A(n_6824),
.B(n_6775),
.C(n_6778),
.Y(n_6882)
);

OA21x2_ASAP7_75t_L g6883 ( 
.A1(n_6824),
.A2(n_6728),
.B(n_6733),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_6832),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_6832),
.Y(n_6885)
);

NAND3xp33_ASAP7_75t_L g6886 ( 
.A(n_6813),
.B(n_6782),
.C(n_6765),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6839),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6811),
.Y(n_6888)
);

OA21x2_ASAP7_75t_L g6889 ( 
.A1(n_6805),
.A2(n_6814),
.B(n_6830),
.Y(n_6889)
);

BUFx2_ASAP7_75t_L g6890 ( 
.A(n_6847),
.Y(n_6890)
);

INVx4_ASAP7_75t_SL g6891 ( 
.A(n_6828),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6808),
.Y(n_6892)
);

BUFx3_ASAP7_75t_L g6893 ( 
.A(n_6808),
.Y(n_6893)
);

INVx2_ASAP7_75t_L g6894 ( 
.A(n_6819),
.Y(n_6894)
);

OAI21x1_ASAP7_75t_L g6895 ( 
.A1(n_6790),
.A2(n_6748),
.B(n_6752),
.Y(n_6895)
);

OA21x2_ASAP7_75t_L g6896 ( 
.A1(n_6830),
.A2(n_6784),
.B(n_6772),
.Y(n_6896)
);

INVx4_ASAP7_75t_SL g6897 ( 
.A(n_6828),
.Y(n_6897)
);

BUFx3_ASAP7_75t_L g6898 ( 
.A(n_6802),
.Y(n_6898)
);

INVx1_ASAP7_75t_SL g6899 ( 
.A(n_6817),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6831),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_6834),
.Y(n_6901)
);

OA21x2_ASAP7_75t_L g6902 ( 
.A1(n_6858),
.A2(n_6760),
.B(n_6776),
.Y(n_6902)
);

INVx3_ASAP7_75t_L g6903 ( 
.A(n_6838),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6838),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6834),
.Y(n_6905)
);

BUFx2_ASAP7_75t_L g6906 ( 
.A(n_6812),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6835),
.Y(n_6907)
);

INVx2_ASAP7_75t_L g6908 ( 
.A(n_6806),
.Y(n_6908)
);

INVx1_ASAP7_75t_L g6909 ( 
.A(n_6835),
.Y(n_6909)
);

NOR3xp33_ASAP7_75t_SL g6910 ( 
.A(n_6800),
.B(n_6844),
.C(n_6798),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6836),
.Y(n_6911)
);

NOR2x1_ASAP7_75t_L g6912 ( 
.A(n_6795),
.B(n_410),
.Y(n_6912)
);

OA21x2_ASAP7_75t_L g6913 ( 
.A1(n_6858),
.A2(n_410),
.B(n_411),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6836),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6837),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6837),
.Y(n_6916)
);

INVx2_ASAP7_75t_L g6917 ( 
.A(n_6806),
.Y(n_6917)
);

AND2x2_ASAP7_75t_L g6918 ( 
.A(n_6803),
.B(n_413),
.Y(n_6918)
);

INVx1_ASAP7_75t_SL g6919 ( 
.A(n_6846),
.Y(n_6919)
);

INVx1_ASAP7_75t_L g6920 ( 
.A(n_6823),
.Y(n_6920)
);

NOR2xp67_ASAP7_75t_L g6921 ( 
.A(n_6878),
.B(n_6842),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6862),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6862),
.Y(n_6923)
);

INVx3_ASAP7_75t_L g6924 ( 
.A(n_6898),
.Y(n_6924)
);

OR2x2_ASAP7_75t_L g6925 ( 
.A(n_6919),
.B(n_6842),
.Y(n_6925)
);

INVx1_ASAP7_75t_L g6926 ( 
.A(n_6906),
.Y(n_6926)
);

NAND2xp5_ASAP7_75t_L g6927 ( 
.A(n_6864),
.B(n_6794),
.Y(n_6927)
);

AND2x2_ASAP7_75t_L g6928 ( 
.A(n_6899),
.B(n_6848),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6864),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6891),
.Y(n_6930)
);

NAND2xp5_ASAP7_75t_L g6931 ( 
.A(n_6860),
.B(n_6813),
.Y(n_6931)
);

NOR2xp33_ASAP7_75t_L g6932 ( 
.A(n_6860),
.B(n_6880),
.Y(n_6932)
);

AND2x2_ASAP7_75t_L g6933 ( 
.A(n_6890),
.B(n_6821),
.Y(n_6933)
);

OR2x6_ASAP7_75t_L g6934 ( 
.A(n_6920),
.B(n_6879),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_6880),
.B(n_6793),
.Y(n_6935)
);

INVx2_ASAP7_75t_L g6936 ( 
.A(n_6891),
.Y(n_6936)
);

INVx1_ASAP7_75t_SL g6937 ( 
.A(n_6889),
.Y(n_6937)
);

NAND2xp5_ASAP7_75t_L g6938 ( 
.A(n_6870),
.B(n_6797),
.Y(n_6938)
);

INVx2_ASAP7_75t_L g6939 ( 
.A(n_6891),
.Y(n_6939)
);

OR2x2_ASAP7_75t_L g6940 ( 
.A(n_6865),
.B(n_6829),
.Y(n_6940)
);

OR2x2_ASAP7_75t_L g6941 ( 
.A(n_6877),
.B(n_6829),
.Y(n_6941)
);

NOR2xp33_ASAP7_75t_L g6942 ( 
.A(n_6869),
.B(n_6809),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6897),
.Y(n_6943)
);

INVx1_ASAP7_75t_L g6944 ( 
.A(n_6897),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6897),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6903),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_6868),
.B(n_6859),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6893),
.Y(n_6948)
);

INVx2_ASAP7_75t_L g6949 ( 
.A(n_6913),
.Y(n_6949)
);

OR2x2_ASAP7_75t_L g6950 ( 
.A(n_6872),
.B(n_6810),
.Y(n_6950)
);

NOR2xp33_ASAP7_75t_L g6951 ( 
.A(n_6866),
.B(n_6810),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6888),
.B(n_6822),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_6894),
.B(n_6816),
.Y(n_6953)
);

OR2x2_ASAP7_75t_L g6954 ( 
.A(n_6892),
.B(n_6840),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6889),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6904),
.Y(n_6956)
);

HB1xp67_ASAP7_75t_L g6957 ( 
.A(n_6875),
.Y(n_6957)
);

BUFx3_ASAP7_75t_L g6958 ( 
.A(n_6918),
.Y(n_6958)
);

AND2x4_ASAP7_75t_L g6959 ( 
.A(n_6871),
.B(n_6827),
.Y(n_6959)
);

NAND2xp5_ASAP7_75t_L g6960 ( 
.A(n_6875),
.B(n_6843),
.Y(n_6960)
);

NOR3xp33_ASAP7_75t_L g6961 ( 
.A(n_6866),
.B(n_6855),
.C(n_6856),
.Y(n_6961)
);

INVx1_ASAP7_75t_L g6962 ( 
.A(n_6912),
.Y(n_6962)
);

BUFx3_ASAP7_75t_L g6963 ( 
.A(n_6874),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6910),
.B(n_6826),
.Y(n_6964)
);

INVx4_ASAP7_75t_L g6965 ( 
.A(n_6881),
.Y(n_6965)
);

INVx2_ASAP7_75t_L g6966 ( 
.A(n_6873),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6900),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6861),
.B(n_6833),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6957),
.B(n_6927),
.Y(n_6969)
);

INVx2_ASAP7_75t_L g6970 ( 
.A(n_6958),
.Y(n_6970)
);

NAND2xp5_ASAP7_75t_SL g6971 ( 
.A(n_6921),
.B(n_6886),
.Y(n_6971)
);

INVx3_ASAP7_75t_L g6972 ( 
.A(n_6924),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6955),
.Y(n_6973)
);

OAI22xp5_ASAP7_75t_L g6974 ( 
.A1(n_6937),
.A2(n_6883),
.B1(n_6882),
.B2(n_6863),
.Y(n_6974)
);

OR2x6_ASAP7_75t_L g6975 ( 
.A(n_6936),
.B(n_6908),
.Y(n_6975)
);

OR2x2_ASAP7_75t_L g6976 ( 
.A(n_6931),
.B(n_6867),
.Y(n_6976)
);

INVx1_ASAP7_75t_SL g6977 ( 
.A(n_6937),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6925),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_6949),
.Y(n_6979)
);

NOR2xp33_ASAP7_75t_SL g6980 ( 
.A(n_6932),
.B(n_6884),
.Y(n_6980)
);

NOR2xp33_ASAP7_75t_L g6981 ( 
.A(n_6962),
.B(n_6917),
.Y(n_6981)
);

AND2x2_ASAP7_75t_L g6982 ( 
.A(n_6933),
.B(n_6928),
.Y(n_6982)
);

OR2x6_ASAP7_75t_L g6983 ( 
.A(n_6939),
.B(n_6885),
.Y(n_6983)
);

AND2x2_ASAP7_75t_L g6984 ( 
.A(n_6952),
.B(n_6876),
.Y(n_6984)
);

INVx3_ASAP7_75t_L g6985 ( 
.A(n_6963),
.Y(n_6985)
);

NOR2xp33_ASAP7_75t_SL g6986 ( 
.A(n_6932),
.B(n_6849),
.Y(n_6986)
);

INVx2_ASAP7_75t_L g6987 ( 
.A(n_6963),
.Y(n_6987)
);

OAI22xp5_ASAP7_75t_L g6988 ( 
.A1(n_6929),
.A2(n_6855),
.B1(n_6852),
.B2(n_6850),
.Y(n_6988)
);

HB1xp67_ASAP7_75t_L g6989 ( 
.A(n_6941),
.Y(n_6989)
);

NAND2xp5_ASAP7_75t_L g6990 ( 
.A(n_6951),
.B(n_6887),
.Y(n_6990)
);

OR2x2_ASAP7_75t_L g6991 ( 
.A(n_6940),
.B(n_6850),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_6951),
.B(n_6901),
.Y(n_6992)
);

NAND2xp5_ASAP7_75t_L g6993 ( 
.A(n_6922),
.B(n_6905),
.Y(n_6993)
);

HB1xp67_ASAP7_75t_L g6994 ( 
.A(n_6930),
.Y(n_6994)
);

NAND2xp5_ASAP7_75t_L g6995 ( 
.A(n_6942),
.B(n_6907),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6960),
.Y(n_6996)
);

OR2x2_ASAP7_75t_L g6997 ( 
.A(n_6954),
.B(n_6857),
.Y(n_6997)
);

CKINVDCx16_ASAP7_75t_R g6998 ( 
.A(n_6947),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6923),
.B(n_6909),
.Y(n_6999)
);

AND2x2_ASAP7_75t_L g7000 ( 
.A(n_6953),
.B(n_6895),
.Y(n_7000)
);

INVx2_ASAP7_75t_L g7001 ( 
.A(n_6943),
.Y(n_7001)
);

INVx2_ASAP7_75t_L g7002 ( 
.A(n_6944),
.Y(n_7002)
);

INVx2_ASAP7_75t_L g7003 ( 
.A(n_6945),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6935),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6982),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_L g7006 ( 
.A(n_6998),
.B(n_6926),
.Y(n_7006)
);

HB1xp67_ASAP7_75t_L g7007 ( 
.A(n_6975),
.Y(n_7007)
);

NAND2x1_ASAP7_75t_L g7008 ( 
.A(n_6985),
.B(n_6934),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6989),
.Y(n_7009)
);

NAND2xp5_ASAP7_75t_L g7010 ( 
.A(n_6984),
.B(n_6965),
.Y(n_7010)
);

NAND2xp5_ASAP7_75t_L g7011 ( 
.A(n_6972),
.B(n_6968),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6969),
.Y(n_7012)
);

NOR2x1_ASAP7_75t_L g7013 ( 
.A(n_6969),
.B(n_6934),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6997),
.Y(n_7014)
);

CKINVDCx16_ASAP7_75t_R g7015 ( 
.A(n_6980),
.Y(n_7015)
);

NAND4xp75_ASAP7_75t_L g7016 ( 
.A(n_7000),
.B(n_6964),
.C(n_6935),
.D(n_6938),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6975),
.Y(n_7017)
);

OAI21xp5_ASAP7_75t_L g7018 ( 
.A1(n_6974),
.A2(n_6961),
.B(n_6946),
.Y(n_7018)
);

INVx2_ASAP7_75t_SL g7019 ( 
.A(n_6970),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6991),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6995),
.Y(n_7021)
);

OR2x2_ASAP7_75t_L g7022 ( 
.A(n_6987),
.B(n_6950),
.Y(n_7022)
);

OR2x2_ASAP7_75t_L g7023 ( 
.A(n_6990),
.B(n_6966),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6990),
.Y(n_7024)
);

AOI22xp5_ASAP7_75t_L g7025 ( 
.A1(n_6996),
.A2(n_6914),
.B1(n_6915),
.B2(n_6911),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6983),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_SL g7027 ( 
.A(n_6980),
.B(n_6966),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6983),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6983),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_7007),
.Y(n_7030)
);

INVxp67_ASAP7_75t_SL g7031 ( 
.A(n_7013),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_7015),
.B(n_6981),
.Y(n_7032)
);

NOR4xp25_ASAP7_75t_L g7033 ( 
.A(n_7027),
.B(n_6977),
.C(n_6971),
.D(n_6979),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_7023),
.Y(n_7034)
);

OAI21xp33_ASAP7_75t_L g7035 ( 
.A1(n_7006),
.A2(n_6986),
.B(n_6978),
.Y(n_7035)
);

AOI22xp5_ASAP7_75t_L g7036 ( 
.A1(n_7013),
.A2(n_6986),
.B1(n_6973),
.B2(n_6916),
.Y(n_7036)
);

AOI21xp5_ASAP7_75t_L g7037 ( 
.A1(n_7008),
.A2(n_6992),
.B(n_6993),
.Y(n_7037)
);

AOI21xp33_ASAP7_75t_L g7038 ( 
.A1(n_7017),
.A2(n_6976),
.B(n_6845),
.Y(n_7038)
);

INVxp67_ASAP7_75t_SL g7039 ( 
.A(n_7011),
.Y(n_7039)
);

OAI221xp5_ASAP7_75t_L g7040 ( 
.A1(n_7018),
.A2(n_6999),
.B1(n_6993),
.B2(n_7004),
.C(n_6853),
.Y(n_7040)
);

OAI21xp5_ASAP7_75t_L g7041 ( 
.A1(n_7016),
.A2(n_6994),
.B(n_6999),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_7022),
.Y(n_7042)
);

NAND2x1p5_ASAP7_75t_L g7043 ( 
.A(n_7014),
.B(n_6959),
.Y(n_7043)
);

AOI22x1_ASAP7_75t_L g7044 ( 
.A1(n_7005),
.A2(n_7001),
.B1(n_7003),
.B2(n_7002),
.Y(n_7044)
);

OAI22xp5_ASAP7_75t_L g7045 ( 
.A1(n_7009),
.A2(n_6967),
.B1(n_6948),
.B2(n_6956),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_7010),
.Y(n_7046)
);

INVx2_ASAP7_75t_L g7047 ( 
.A(n_7024),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_7012),
.B(n_6815),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_7043),
.Y(n_7049)
);

NOR2xp33_ASAP7_75t_L g7050 ( 
.A(n_7031),
.B(n_7026),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_7048),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_7034),
.Y(n_7052)
);

AOI21xp33_ASAP7_75t_L g7053 ( 
.A1(n_7030),
.A2(n_7029),
.B(n_7028),
.Y(n_7053)
);

AND2x2_ASAP7_75t_L g7054 ( 
.A(n_7042),
.B(n_7019),
.Y(n_7054)
);

AOI221xp5_ASAP7_75t_L g7055 ( 
.A1(n_7033),
.A2(n_7038),
.B1(n_6988),
.B2(n_7037),
.C(n_7036),
.Y(n_7055)
);

NAND2xp5_ASAP7_75t_L g7056 ( 
.A(n_7039),
.B(n_7021),
.Y(n_7056)
);

INVxp67_ASAP7_75t_SL g7057 ( 
.A(n_7032),
.Y(n_7057)
);

INVxp67_ASAP7_75t_SL g7058 ( 
.A(n_7041),
.Y(n_7058)
);

NOR2xp33_ASAP7_75t_SL g7059 ( 
.A(n_7035),
.B(n_7020),
.Y(n_7059)
);

AND2x4_ASAP7_75t_L g7060 ( 
.A(n_7047),
.B(n_6818),
.Y(n_7060)
);

OR2x2_ASAP7_75t_L g7061 ( 
.A(n_7045),
.B(n_6854),
.Y(n_7061)
);

AND2x4_ASAP7_75t_SL g7062 ( 
.A(n_7046),
.B(n_7025),
.Y(n_7062)
);

INVx2_ASAP7_75t_L g7063 ( 
.A(n_7060),
.Y(n_7063)
);

OAI22xp5_ASAP7_75t_L g7064 ( 
.A1(n_7058),
.A2(n_7040),
.B1(n_7044),
.B2(n_6825),
.Y(n_7064)
);

AND2x2_ASAP7_75t_L g7065 ( 
.A(n_7054),
.B(n_6902),
.Y(n_7065)
);

OAI21xp33_ASAP7_75t_SL g7066 ( 
.A1(n_7055),
.A2(n_6896),
.B(n_415),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_7062),
.Y(n_7067)
);

INVx1_ASAP7_75t_SL g7068 ( 
.A(n_7061),
.Y(n_7068)
);

OR2x2_ASAP7_75t_L g7069 ( 
.A(n_7049),
.B(n_7052),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_7057),
.Y(n_7070)
);

AOI22xp5_ASAP7_75t_L g7071 ( 
.A1(n_7050),
.A2(n_7051),
.B1(n_7056),
.B2(n_7059),
.Y(n_7071)
);

AOI221xp5_ASAP7_75t_L g7072 ( 
.A1(n_7053),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_7072)
);

AND2x4_ASAP7_75t_SL g7073 ( 
.A(n_7067),
.B(n_2819),
.Y(n_7073)
);

OAI221xp5_ASAP7_75t_L g7074 ( 
.A1(n_7071),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.C(n_430),
.Y(n_7074)
);

O2A1O1Ixp5_ASAP7_75t_L g7075 ( 
.A1(n_7070),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_7075)
);

AND2x2_ASAP7_75t_L g7076 ( 
.A(n_7065),
.B(n_431),
.Y(n_7076)
);

OAI221xp5_ASAP7_75t_L g7077 ( 
.A1(n_7066),
.A2(n_437),
.B1(n_439),
.B2(n_440),
.C(n_441),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_L g7078 ( 
.A(n_7068),
.B(n_445),
.Y(n_7078)
);

NOR2xp33_ASAP7_75t_L g7079 ( 
.A(n_7063),
.B(n_446),
.Y(n_7079)
);

AOI32xp33_ASAP7_75t_L g7080 ( 
.A1(n_7064),
.A2(n_447),
.A3(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_7072),
.B(n_455),
.Y(n_7081)
);

INVx3_ASAP7_75t_L g7082 ( 
.A(n_7069),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_7082),
.Y(n_7083)
);

OAI221xp5_ASAP7_75t_L g7084 ( 
.A1(n_7080),
.A2(n_464),
.B1(n_465),
.B2(n_466),
.C(n_467),
.Y(n_7084)
);

NOR3x1_ASAP7_75t_L g7085 ( 
.A(n_7074),
.B(n_7077),
.C(n_7081),
.Y(n_7085)
);

AOI21xp5_ASAP7_75t_L g7086 ( 
.A1(n_7078),
.A2(n_466),
.B(n_467),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_7075),
.Y(n_7087)
);

A2O1A1Ixp33_ASAP7_75t_L g7088 ( 
.A1(n_7079),
.A2(n_473),
.B(n_470),
.C(n_471),
.Y(n_7088)
);

OAI21xp33_ASAP7_75t_L g7089 ( 
.A1(n_7073),
.A2(n_474),
.B(n_476),
.Y(n_7089)
);

OAI21xp33_ASAP7_75t_L g7090 ( 
.A1(n_7082),
.A2(n_478),
.B(n_479),
.Y(n_7090)
);

AOI221xp5_ASAP7_75t_L g7091 ( 
.A1(n_7082),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.C(n_483),
.Y(n_7091)
);

AND2x2_ASAP7_75t_L g7092 ( 
.A(n_7082),
.B(n_480),
.Y(n_7092)
);

AOI211xp5_ASAP7_75t_SL g7093 ( 
.A1(n_7082),
.A2(n_484),
.B(n_485),
.C(n_486),
.Y(n_7093)
);

HB1xp67_ASAP7_75t_L g7094 ( 
.A(n_7082),
.Y(n_7094)
);

OAI21xp5_ASAP7_75t_L g7095 ( 
.A1(n_7076),
.A2(n_486),
.B(n_487),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_7094),
.B(n_487),
.Y(n_7096)
);

OAI211xp5_ASAP7_75t_L g7097 ( 
.A1(n_7083),
.A2(n_488),
.B(n_489),
.C(n_490),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_L g7098 ( 
.A(n_7087),
.B(n_490),
.Y(n_7098)
);

NOR3x1_ASAP7_75t_L g7099 ( 
.A(n_7095),
.B(n_496),
.C(n_497),
.Y(n_7099)
);

O2A1O1Ixp33_ASAP7_75t_SL g7100 ( 
.A1(n_7088),
.A2(n_498),
.B(n_499),
.C(n_500),
.Y(n_7100)
);

AOI21xp5_ASAP7_75t_L g7101 ( 
.A1(n_7090),
.A2(n_499),
.B(n_501),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_7092),
.Y(n_7102)
);

NAND3xp33_ASAP7_75t_L g7103 ( 
.A(n_7093),
.B(n_1593),
.C(n_1585),
.Y(n_7103)
);

NAND3xp33_ASAP7_75t_L g7104 ( 
.A(n_7086),
.B(n_2324),
.C(n_2314),
.Y(n_7104)
);

OAI22xp5_ASAP7_75t_L g7105 ( 
.A1(n_7084),
.A2(n_503),
.B1(n_504),
.B2(n_506),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_7089),
.B(n_507),
.Y(n_7106)
);

O2A1O1Ixp33_ASAP7_75t_SL g7107 ( 
.A1(n_7091),
.A2(n_512),
.B(n_513),
.C(n_514),
.Y(n_7107)
);

NAND2xp5_ASAP7_75t_L g7108 ( 
.A(n_7102),
.B(n_7096),
.Y(n_7108)
);

AND2x2_ASAP7_75t_L g7109 ( 
.A(n_7099),
.B(n_7085),
.Y(n_7109)
);

NOR2x1_ASAP7_75t_L g7110 ( 
.A(n_7097),
.B(n_516),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_7100),
.Y(n_7111)
);

INVxp67_ASAP7_75t_L g7112 ( 
.A(n_7106),
.Y(n_7112)
);

NAND2xp5_ASAP7_75t_L g7113 ( 
.A(n_7101),
.B(n_7107),
.Y(n_7113)
);

NAND2xp5_ASAP7_75t_L g7114 ( 
.A(n_7105),
.B(n_518),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_7104),
.Y(n_7115)
);

AOI21xp33_ASAP7_75t_L g7116 ( 
.A1(n_7103),
.A2(n_522),
.B(n_524),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_7096),
.Y(n_7117)
);

NAND3xp33_ASAP7_75t_SL g7118 ( 
.A(n_7098),
.B(n_524),
.C(n_525),
.Y(n_7118)
);

NOR3xp33_ASAP7_75t_L g7119 ( 
.A(n_7108),
.B(n_526),
.C(n_528),
.Y(n_7119)
);

NAND2xp5_ASAP7_75t_SL g7120 ( 
.A(n_7111),
.B(n_2522),
.Y(n_7120)
);

NOR2xp33_ASAP7_75t_L g7121 ( 
.A(n_7112),
.B(n_7118),
.Y(n_7121)
);

NAND4xp25_ASAP7_75t_L g7122 ( 
.A(n_7110),
.B(n_529),
.C(n_530),
.D(n_532),
.Y(n_7122)
);

NOR2x1_ASAP7_75t_L g7123 ( 
.A(n_7113),
.B(n_533),
.Y(n_7123)
);

NOR3xp33_ASAP7_75t_L g7124 ( 
.A(n_7115),
.B(n_7114),
.C(n_7116),
.Y(n_7124)
);

NAND2xp5_ASAP7_75t_L g7125 ( 
.A(n_7117),
.B(n_535),
.Y(n_7125)
);

AND2x4_ASAP7_75t_L g7126 ( 
.A(n_7109),
.B(n_539),
.Y(n_7126)
);

NOR3x1_ASAP7_75t_L g7127 ( 
.A(n_7118),
.B(n_542),
.C(n_543),
.Y(n_7127)
);

NAND4xp75_ASAP7_75t_L g7128 ( 
.A(n_7109),
.B(n_543),
.C(n_544),
.D(n_545),
.Y(n_7128)
);

NOR3xp33_ASAP7_75t_L g7129 ( 
.A(n_7108),
.B(n_545),
.C(n_546),
.Y(n_7129)
);

AND4x1_ASAP7_75t_L g7130 ( 
.A(n_7109),
.B(n_547),
.C(n_549),
.D(n_550),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_7123),
.Y(n_7131)
);

AOI21xp5_ASAP7_75t_L g7132 ( 
.A1(n_7125),
.A2(n_554),
.B(n_555),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_L g7133 ( 
.A(n_7121),
.B(n_558),
.Y(n_7133)
);

AOI21xp33_ASAP7_75t_SL g7134 ( 
.A1(n_7126),
.A2(n_558),
.B(n_559),
.Y(n_7134)
);

AND2x2_ASAP7_75t_L g7135 ( 
.A(n_7127),
.B(n_559),
.Y(n_7135)
);

NAND3xp33_ASAP7_75t_L g7136 ( 
.A(n_7124),
.B(n_2324),
.C(n_562),
.Y(n_7136)
);

OR2x2_ASAP7_75t_L g7137 ( 
.A(n_7122),
.B(n_561),
.Y(n_7137)
);

NAND2xp5_ASAP7_75t_L g7138 ( 
.A(n_7130),
.B(n_563),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_7119),
.B(n_564),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_7128),
.Y(n_7140)
);

INVx2_ASAP7_75t_SL g7141 ( 
.A(n_7120),
.Y(n_7141)
);

AND2x2_ASAP7_75t_L g7142 ( 
.A(n_7129),
.B(n_564),
.Y(n_7142)
);

AND2x2_ASAP7_75t_L g7143 ( 
.A(n_7131),
.B(n_567),
.Y(n_7143)
);

NAND4xp25_ASAP7_75t_SL g7144 ( 
.A(n_7138),
.B(n_568),
.C(n_569),
.D(n_570),
.Y(n_7144)
);

OA22x2_ASAP7_75t_L g7145 ( 
.A1(n_7135),
.A2(n_570),
.B1(n_572),
.B2(n_574),
.Y(n_7145)
);

NOR2xp67_ASAP7_75t_L g7146 ( 
.A(n_7134),
.B(n_7132),
.Y(n_7146)
);

NOR2x1p5_ASAP7_75t_L g7147 ( 
.A(n_7137),
.B(n_580),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_7133),
.Y(n_7148)
);

INVx2_ASAP7_75t_L g7149 ( 
.A(n_7142),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_7140),
.B(n_582),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_7146),
.Y(n_7151)
);

AOI22xp5_ASAP7_75t_L g7152 ( 
.A1(n_7144),
.A2(n_7139),
.B1(n_7141),
.B2(n_7136),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_7147),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_7145),
.Y(n_7154)
);

NOR2x1_ASAP7_75t_L g7155 ( 
.A(n_7151),
.B(n_7149),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_7153),
.Y(n_7156)
);

INVx2_ASAP7_75t_L g7157 ( 
.A(n_7154),
.Y(n_7157)
);

NAND2x1p5_ASAP7_75t_L g7158 ( 
.A(n_7152),
.B(n_7148),
.Y(n_7158)
);

OAI211xp5_ASAP7_75t_SL g7159 ( 
.A1(n_7156),
.A2(n_7150),
.B(n_7143),
.C(n_584),
.Y(n_7159)
);

NAND4xp75_ASAP7_75t_L g7160 ( 
.A(n_7158),
.B(n_584),
.C(n_585),
.D(n_586),
.Y(n_7160)
);

OR3x2_ASAP7_75t_L g7161 ( 
.A(n_7156),
.B(n_585),
.C(n_587),
.Y(n_7161)
);

NOR3xp33_ASAP7_75t_L g7162 ( 
.A(n_7155),
.B(n_588),
.C(n_589),
.Y(n_7162)
);

NOR2x1p5_ASAP7_75t_L g7163 ( 
.A(n_7157),
.B(n_590),
.Y(n_7163)
);

NOR2x1_ASAP7_75t_L g7164 ( 
.A(n_7157),
.B(n_590),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_L g7165 ( 
.A(n_7155),
.B(n_591),
.Y(n_7165)
);

NOR3xp33_ASAP7_75t_L g7166 ( 
.A(n_7155),
.B(n_592),
.C(n_594),
.Y(n_7166)
);

NAND3x1_ASAP7_75t_L g7167 ( 
.A(n_7164),
.B(n_592),
.C(n_594),
.Y(n_7167)
);

OAI22xp5_ASAP7_75t_L g7168 ( 
.A1(n_7161),
.A2(n_7163),
.B1(n_7165),
.B2(n_7160),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_7159),
.Y(n_7169)
);

XNOR2xp5_ASAP7_75t_L g7170 ( 
.A(n_7162),
.B(n_595),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_7166),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_7164),
.Y(n_7172)
);

NOR2x1p5_ASAP7_75t_L g7173 ( 
.A(n_7172),
.B(n_7169),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_7168),
.Y(n_7174)
);

OAI22x1_ASAP7_75t_L g7175 ( 
.A1(n_7173),
.A2(n_7171),
.B1(n_7170),
.B2(n_7167),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_7174),
.Y(n_7176)
);

OAI22xp5_ASAP7_75t_SL g7177 ( 
.A1(n_7175),
.A2(n_610),
.B1(n_612),
.B2(n_614),
.Y(n_7177)
);

INVx4_ASAP7_75t_L g7178 ( 
.A(n_7176),
.Y(n_7178)
);

INVx2_ASAP7_75t_SL g7179 ( 
.A(n_7176),
.Y(n_7179)
);

OAI22xp5_ASAP7_75t_SL g7180 ( 
.A1(n_7176),
.A2(n_624),
.B1(n_625),
.B2(n_626),
.Y(n_7180)
);

OAI22xp5_ASAP7_75t_SL g7181 ( 
.A1(n_7176),
.A2(n_627),
.B1(n_630),
.B2(n_631),
.Y(n_7181)
);

AND2x4_ASAP7_75t_L g7182 ( 
.A(n_7176),
.B(n_631),
.Y(n_7182)
);

OA22x2_ASAP7_75t_L g7183 ( 
.A1(n_7179),
.A2(n_632),
.B1(n_633),
.B2(n_634),
.Y(n_7183)
);

INVx2_ASAP7_75t_L g7184 ( 
.A(n_7178),
.Y(n_7184)
);

HB1xp67_ASAP7_75t_L g7185 ( 
.A(n_7182),
.Y(n_7185)
);

AOI22xp5_ASAP7_75t_L g7186 ( 
.A1(n_7184),
.A2(n_7177),
.B1(n_7180),
.B2(n_7181),
.Y(n_7186)
);

AOI22xp33_ASAP7_75t_L g7187 ( 
.A1(n_7185),
.A2(n_637),
.B1(n_642),
.B2(n_643),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_7183),
.Y(n_7188)
);

O2A1O1Ixp5_ASAP7_75t_L g7189 ( 
.A1(n_7184),
.A2(n_649),
.B(n_651),
.C(n_1428),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_7188),
.Y(n_7190)
);

OAI21xp5_ASAP7_75t_SL g7191 ( 
.A1(n_7186),
.A2(n_651),
.B(n_2113),
.Y(n_7191)
);

OAI21xp5_ASAP7_75t_L g7192 ( 
.A1(n_7189),
.A2(n_2085),
.B(n_2122),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_7190),
.Y(n_7193)
);

INVx2_ASAP7_75t_L g7194 ( 
.A(n_7193),
.Y(n_7194)
);

AOI22x1_ASAP7_75t_L g7195 ( 
.A1(n_7194),
.A2(n_7192),
.B1(n_7191),
.B2(n_7187),
.Y(n_7195)
);

NAND2xp5_ASAP7_75t_L g7196 ( 
.A(n_7195),
.B(n_2085),
.Y(n_7196)
);

OAI21xp5_ASAP7_75t_L g7197 ( 
.A1(n_7195),
.A2(n_2122),
.B(n_2133),
.Y(n_7197)
);

AOI22x1_ASAP7_75t_L g7198 ( 
.A1(n_7195),
.A2(n_2101),
.B1(n_2113),
.B2(n_2121),
.Y(n_7198)
);

INVx2_ASAP7_75t_L g7199 ( 
.A(n_7196),
.Y(n_7199)
);

INVxp67_ASAP7_75t_SL g7200 ( 
.A(n_7197),
.Y(n_7200)
);

AOI21xp5_ASAP7_75t_L g7201 ( 
.A1(n_7200),
.A2(n_7198),
.B(n_2133),
.Y(n_7201)
);

OR2x6_ASAP7_75t_L g7202 ( 
.A(n_7199),
.B(n_2101),
.Y(n_7202)
);

AOI221xp5_ASAP7_75t_L g7203 ( 
.A1(n_7201),
.A2(n_2133),
.B1(n_2113),
.B2(n_2121),
.C(n_2101),
.Y(n_7203)
);

AOI22xp33_ASAP7_75t_SL g7204 ( 
.A1(n_7202),
.A2(n_2113),
.B1(n_2121),
.B2(n_2134),
.Y(n_7204)
);

AOI21xp5_ASAP7_75t_L g7205 ( 
.A1(n_7203),
.A2(n_2134),
.B(n_2522),
.Y(n_7205)
);

AOI211xp5_ASAP7_75t_L g7206 ( 
.A1(n_7205),
.A2(n_7204),
.B(n_2134),
.C(n_2543),
.Y(n_7206)
);


endmodule