module fake_jpeg_30604_n_444 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_444);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_17),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_74),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_32),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_88),
.Y(n_132)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_31),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_33),
.B(n_15),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_1),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_27),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_37),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_37),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_135),
.Y(n_165)
);

BUFx16f_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_49),
.B(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_45),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_46),
.Y(n_137)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_80),
.B1(n_67),
.B2(n_85),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_154),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_48),
.B1(n_47),
.B2(n_52),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_151),
.B(n_167),
.Y(n_180)
);

HAxp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_49),
.CON(n_141),
.SN(n_141)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_145),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_91),
.A2(n_53),
.B1(n_64),
.B2(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_160),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_34),
.B(n_20),
.C(n_41),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_162),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_51),
.B(n_63),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_152),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_66),
.B1(n_28),
.B2(n_31),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_96),
.A2(n_28),
.B1(n_31),
.B2(n_19),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_43),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_60),
.C(n_75),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_124),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_94),
.A2(n_79),
.B1(n_68),
.B2(n_59),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_86),
.B1(n_55),
.B2(n_28),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_175),
.B1(n_152),
.B2(n_143),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_87),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_173),
.Y(n_177)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_198),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_187),
.B1(n_194),
.B2(n_171),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_151),
.A2(n_93),
.B1(n_131),
.B2(n_105),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_191),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_93),
.B1(n_131),
.B2(n_105),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_138),
.C(n_109),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_111),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_114),
.B(n_118),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_212),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_195),
.B(n_193),
.C(n_192),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_158),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_213),
.Y(n_250)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_11),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_140),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_223),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_178),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_140),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_140),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_185),
.B(n_192),
.Y(n_247)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_191),
.C(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_224),
.C(n_219),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_180),
.B1(n_200),
.B2(n_183),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_240),
.B1(n_134),
.B2(n_175),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_180),
.B1(n_203),
.B2(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_244),
.B1(n_219),
.B2(n_210),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_183),
.B1(n_182),
.B2(n_203),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_185),
.B1(n_177),
.B2(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_114),
.B(n_153),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_182),
.B1(n_170),
.B2(n_189),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_211),
.B(n_190),
.Y(n_260)
);

XOR2x1_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_195),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_185),
.B(n_181),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_208),
.B(n_207),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_253),
.A2(n_243),
.B1(n_245),
.B2(n_247),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_256),
.C(n_262),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_260),
.A2(n_280),
.B(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_226),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_273),
.C(n_251),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_218),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

AO22x1_ASAP7_75t_SL g267 ( 
.A1(n_232),
.A2(n_228),
.B1(n_209),
.B2(n_213),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_236),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_271),
.B(n_244),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_196),
.C(n_181),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_248),
.Y(n_287)
);

OR2x4_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_202),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_228),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_202),
.C(n_193),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_209),
.Y(n_274)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_155),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_55),
.A3(n_137),
.B1(n_24),
.B2(n_58),
.Y(n_277)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_241),
.B1(n_245),
.B2(n_229),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_24),
.C(n_13),
.D(n_14),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_300),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_221),
.B(n_213),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_270),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_291),
.A2(n_299),
.B1(n_306),
.B2(n_107),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_298),
.B1(n_302),
.B2(n_307),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_295),
.A2(n_277),
.B(n_250),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_229),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_24),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_148),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_265),
.A2(n_236),
.B1(n_238),
.B2(n_251),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_173),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_257),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_143),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_238),
.B1(n_250),
.B2(n_233),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_267),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_253),
.A2(n_267),
.B1(n_278),
.B2(n_271),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_258),
.A2(n_250),
.B1(n_233),
.B2(n_214),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_311),
.B(n_332),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_255),
.C(n_263),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_313),
.C(n_314),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_262),
.C(n_261),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_259),
.C(n_274),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_282),
.A2(n_276),
.B1(n_266),
.B2(n_280),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_288),
.B1(n_284),
.B2(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_320),
.B(n_324),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_233),
.B(n_221),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_331),
.C(n_293),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_143),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_334),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_309),
.A2(n_179),
.B1(n_153),
.B2(n_166),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_323),
.A2(n_291),
.B1(n_306),
.B2(n_308),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_330),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_299),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_328),
.B(n_329),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_163),
.C(n_130),
.Y(n_331)
);

XNOR2x2_ASAP7_75t_SL g332 ( 
.A(n_287),
.B(n_24),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_168),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_292),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_335),
.A2(n_342),
.B1(n_357),
.B2(n_331),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_323),
.A2(n_303),
.B1(n_283),
.B2(n_289),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_355),
.A3(n_325),
.B1(n_320),
.B2(n_319),
.C1(n_333),
.C2(n_169),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_353),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_310),
.A2(n_286),
.B1(n_304),
.B2(n_292),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_344),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_321),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_283),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_356),
.C(n_163),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_304),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_358),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_147),
.B1(n_144),
.B2(n_107),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_24),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_324),
.A2(n_101),
.B1(n_95),
.B2(n_94),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_41),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_367),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_362),
.A2(n_365),
.B1(n_373),
.B2(n_344),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_311),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_370),
.Y(n_389)
);

OA21x2_ASAP7_75t_SL g364 ( 
.A1(n_339),
.A2(n_322),
.B(n_332),
.Y(n_364)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_343),
.B(n_334),
.Y(n_366)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_338),
.A2(n_95),
.B1(n_35),
.B2(n_19),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_117),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_117),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_374),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_346),
.B(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_378),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_337),
.A2(n_156),
.B1(n_134),
.B2(n_116),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_125),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_116),
.B(n_120),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_375),
.A2(n_357),
.B(n_349),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_130),
.C(n_129),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_352),
.C(n_347),
.Y(n_383)
);

INVx11_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_368),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_35),
.B1(n_43),
.B2(n_20),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_347),
.CI(n_353),
.CON(n_380),
.SN(n_380)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_384),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_383),
.B(n_388),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_335),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_394),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_359),
.B(n_370),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_351),
.B(n_12),
.Y(n_390)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_371),
.C(n_365),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_382),
.B(n_368),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_398),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_392),
.A2(n_351),
.B1(n_361),
.B2(n_360),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_388),
.A2(n_360),
.B(n_374),
.Y(n_400)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_375),
.B(n_366),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_403),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_SL g404 ( 
.A(n_386),
.B(n_373),
.C(n_376),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_404),
.A2(n_380),
.B1(n_393),
.B2(n_387),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_383),
.A2(n_35),
.B1(n_34),
.B2(n_125),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_393),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_14),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_11),
.Y(n_411)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_418),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_396),
.B(n_381),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_411),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_402),
.A2(n_380),
.B1(n_381),
.B2(n_389),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_413),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_399),
.A2(n_389),
.B(n_81),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_13),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_417),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_402),
.A2(n_57),
.B(n_12),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_112),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_397),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_427),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_401),
.C(n_407),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_423),
.A2(n_428),
.B(n_409),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_416),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_403),
.C(n_404),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_38),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_425),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_38),
.A3(n_112),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_2),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_417),
.B(n_12),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_433),
.B(n_434),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_428),
.A2(n_1),
.B(n_2),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_424),
.A2(n_426),
.B(n_421),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_435),
.A2(n_436),
.B(n_438),
.Y(n_439)
);

AOI322xp5_ASAP7_75t_L g438 ( 
.A1(n_429),
.A2(n_38),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_2),
.C2(n_8),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_437),
.A2(n_4),
.B(n_5),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_440),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_441)
);

OAI322xp33_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_4),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_439),
.C2(n_301),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_9),
.C(n_10),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_443),
.B(n_9),
.Y(n_444)
);


endmodule