module fake_jpeg_23666_n_132 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_18),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_13),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_16),
.B(n_19),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_49),
.C(n_34),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_32),
.A3(n_34),
.B1(n_27),
.B2(n_37),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_27),
.B1(n_24),
.B2(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_13),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_32),
.C(n_33),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.C(n_44),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.C(n_66),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_48),
.B1(n_42),
.B2(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_11),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_37),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_89),
.C(n_85),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_34),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_63),
.C(n_57),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_90),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_79),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_34),
.C(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_67),
.B(n_72),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_102),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_72),
.C(n_67),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_69),
.A3(n_21),
.B1(n_11),
.B2(n_43),
.C1(n_15),
.C2(n_13),
.Y(n_102)
);

AOI321xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_83),
.A3(n_89),
.B1(n_81),
.B2(n_87),
.C(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_106),
.Y(n_112)
);

AOI21x1_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_101),
.B(n_94),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_110),
.B(n_12),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_12),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_12),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_118),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_15),
.B1(n_21),
.B2(n_2),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_97),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_111),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_7),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_109),
.C(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_108),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_6),
.A3(n_9),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_10),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.C(n_127),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_1),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_119),
.C(n_7),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_128),
.Y(n_132)
);


endmodule