module real_jpeg_7474_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_92),
.B1(n_141),
.B2(n_193),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_2),
.A2(n_92),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_2),
.A2(n_92),
.B1(n_424),
.B2(n_426),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_79),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_79),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_4),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_156),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_4),
.A2(n_119),
.B1(n_156),
.B2(n_212),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_4),
.A2(n_156),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_5),
.A2(n_93),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_5),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_5),
.A2(n_177),
.B1(n_202),
.B2(n_259),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_5),
.A2(n_202),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_5),
.A2(n_202),
.B1(n_362),
.B2(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_47),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_6),
.A2(n_47),
.B1(n_371),
.B2(n_408),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_7),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_7),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_7),
.B(n_77),
.C(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_7),
.B(n_142),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_7),
.B(n_265),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_7),
.B(n_86),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_7),
.B(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_9),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_9),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_10),
.A2(n_190),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_10),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_10),
.A2(n_274),
.B1(n_291),
.B2(n_294),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_10),
.A2(n_274),
.B1(n_360),
.B2(n_362),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_10),
.A2(n_212),
.B1(n_274),
.B2(n_447),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_38),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_12),
.Y(n_392)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_14),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_14),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_15),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_15),
.A2(n_111),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_15),
.A2(n_111),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_15),
.A2(n_111),
.B1(n_152),
.B2(n_162),
.Y(n_331)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_232),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_230),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_204),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_20),
.B(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_124),
.C(n_173),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_21),
.A2(n_22),
.B1(n_124),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_87),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_23),
.A2(n_24),
.B(n_89),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_88),
.B1(n_89),
.B2(n_123),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_24),
.A2(n_45),
.B1(n_123),
.B2(n_435),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_25),
.A2(n_37),
.B1(n_176),
.B2(n_181),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_25),
.A2(n_258),
.B(n_263),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_25),
.A2(n_244),
.B(n_263),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_25),
.A2(n_402),
.B1(n_403),
.B2(n_406),
.Y(n_401)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_26),
.B(n_266),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_26),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_26),
.A2(n_335),
.B1(n_370),
.B2(n_373),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_26),
.A2(n_407),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_39),
.Y(n_371)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_41),
.Y(n_177)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_42),
.Y(n_408)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_43),
.Y(n_337)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_44),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_45),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_56),
.B1(n_78),
.B2(n_86),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_46),
.A2(n_56),
.B1(n_86),
.B2(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_55),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_55),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_56),
.A2(n_78),
.B1(n_86),
.B2(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_56),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_56),
.B(n_246),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_60),
.Y(n_189)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g190 ( 
.A(n_66),
.Y(n_190)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_69),
.A2(n_273),
.B(n_276),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_72),
.Y(n_269)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g348 ( 
.A(n_82),
.B(n_138),
.Y(n_348)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_85),
.Y(n_252)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_86),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_109),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_93),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_97),
.B(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_97),
.Y(n_210)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_104),
.B2(n_107),
.Y(n_98)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_99),
.Y(n_394)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_103),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_103),
.Y(n_329)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_109),
.A2(n_210),
.B(n_446),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_115),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_115),
.A2(n_415),
.B(n_416),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_124),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_163),
.B(n_172),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_164),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_142),
.B1(n_150),
.B2(n_157),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_127),
.A2(n_324),
.B(n_330),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_127),
.B(n_366),
.Y(n_365)
);

AOI22x1_ASAP7_75t_L g449 ( 
.A1(n_127),
.A2(n_142),
.B1(n_366),
.B2(n_450),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_127),
.A2(n_330),
.B(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_151),
.B1(n_192),
.B2(n_197),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_128),
.A2(n_197),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_128),
.A2(n_197),
.B1(n_359),
.B2(n_419),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_137),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_142),
.Y(n_197)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g275 ( 
.A(n_144),
.Y(n_275)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_149),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_155),
.Y(n_364)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g361 ( 
.A(n_160),
.Y(n_361)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_171),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_205),
.CI(n_206),
.CON(n_204),
.SN(n_204)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_173),
.B(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_191),
.C(n_198),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_174),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_185),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_175),
.B(n_185),
.Y(n_460)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_176),
.Y(n_441)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_184),
.Y(n_307)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_184),
.Y(n_405)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_186),
.Y(n_439)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_190),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_191),
.B(n_198),
.Y(n_433)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_192),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_197),
.B(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_197),
.A2(n_359),
.B(n_365),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B(n_203),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_199),
.A2(n_200),
.B1(n_210),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_203),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_204),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_214),
.B2(n_229),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_210),
.B(n_244),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_SL g415 ( 
.A1(n_212),
.A2(n_244),
.B(n_397),
.Y(n_415)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_228),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_241),
.B(n_245),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_216),
.A2(n_217),
.B1(n_273),
.B2(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_216),
.A2(n_245),
.B(n_318),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_216),
.A2(n_217),
.B1(n_423),
.B2(n_439),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_217),
.A2(n_276),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI311xp33_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_429),
.A3(n_468),
.B1(n_486),
.C1(n_491),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_377),
.B(n_428),
.Y(n_234)
);

AO21x1_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_350),
.B(n_376),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_312),
.B(n_349),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_279),
.B(n_311),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_256),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_239),
.B(n_256),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_250),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_240),
.A2(n_250),
.B1(n_251),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_244),
.A2(n_325),
.B(n_327),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_244),
.B(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_249),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_270),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_271),
.C(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_258),
.Y(n_305)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_277),
.B2(n_278),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_302),
.B(n_310),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_288),
.B(n_301),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_300),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_296),
.B(n_299),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_298),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_334),
.B(n_339),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_308),
.Y(n_310)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_314),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_332),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_322),
.B2(n_323),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_322),
.C(n_332),
.Y(n_351)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_326),
.Y(n_396)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_341),
.A3(n_342),
.B1(n_345),
.B2(n_348),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_351),
.B(n_352),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_357),
.B2(n_375),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_356),
.C(n_375),
.Y(n_378)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_367),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_368),
.C(n_369),
.Y(n_409)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_378),
.B(n_379),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_412),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_380)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_400),
.B2(n_401),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_383),
.B(n_400),
.Y(n_464)
);

OAI32xp33_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_387),
.A3(n_390),
.B1(n_393),
.B2(n_397),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_409),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_410),
.C(n_412),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_414),
.B1(n_417),
.B2(n_427),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_413),
.B(n_418),
.C(n_422),
.Y(n_477)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_422),
.Y(n_417)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_454),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_430),
.A2(n_454),
.B(n_487),
.C(n_490),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_451),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_451),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.C(n_436),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g467 ( 
.A(n_432),
.B(n_434),
.CI(n_436),
.CON(n_467),
.SN(n_467)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_444),
.C(n_449),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_444),
.A2(n_445),
.B1(n_449),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_467),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_467),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.C(n_461),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_457),
.B1(n_460),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.C(n_465),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_462),
.A2(n_463),
.B1(n_465),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_465),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_467),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_481),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_478),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_478),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.C(n_477),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_484),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_475),
.A2(n_476),
.B1(n_477),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_483),
.Y(n_488)
);


endmodule