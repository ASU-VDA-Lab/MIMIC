module fake_jpeg_18190_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_36),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

OAI211xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_34),
.B(n_31),
.C(n_19),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_35),
.C(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_53),
.B1(n_58),
.B2(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_20),
.C(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_67),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_71),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_60),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_80),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_93),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_22),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_44),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_41),
.CI(n_44),
.CON(n_105),
.SN(n_105)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_50),
.B1(n_51),
.B2(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_121),
.B1(n_84),
.B2(n_74),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_64),
.C(n_47),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_107),
.C(n_105),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_67),
.B(n_49),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_64),
.B(n_75),
.Y(n_145)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_47),
.Y(n_131)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_75),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_63),
.B1(n_44),
.B2(n_41),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_120),
.B1(n_87),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_41),
.B1(n_65),
.B2(n_21),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_23),
.B1(n_17),
.B2(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_131),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_140),
.B1(n_98),
.B2(n_106),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_81),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_135),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_76),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_70),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_20),
.C(n_72),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_74),
.B1(n_68),
.B2(n_90),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_94),
.B(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_139),
.B(n_135),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_104),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_149),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_98),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_64),
.C(n_29),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_29),
.C(n_33),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_161),
.B1(n_179),
.B2(n_181),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_167),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_176),
.C(n_127),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_118),
.B(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_114),
.B1(n_97),
.B2(n_113),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_162),
.B1(n_177),
.B2(n_167),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_120),
.A3(n_114),
.B1(n_121),
.B2(n_115),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_172),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_119),
.B(n_110),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_165),
.B(n_122),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_115),
.B1(n_113),
.B2(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_119),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_150),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_99),
.B1(n_103),
.B2(n_29),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_170),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_0),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_29),
.A3(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_133),
.B1(n_143),
.B2(n_138),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_24),
.C(n_17),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_124),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_123),
.B1(n_140),
.B2(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_24),
.B1(n_73),
.B2(n_2),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_189),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_188),
.B(n_197),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_202),
.B1(n_151),
.B2(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_141),
.B(n_142),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_193),
.C(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_138),
.C(n_73),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_73),
.B(n_1),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_199),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_200),
.B(n_204),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_8),
.C(n_15),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_8),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_178),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_2),
.B(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_155),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_158),
.B1(n_153),
.B2(n_163),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_213),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_180),
.B(n_152),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_218),
.B(n_219),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_161),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_196),
.B1(n_206),
.B2(n_204),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_179),
.C(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_233),
.C(n_194),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_175),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_7),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_227),
.B1(n_184),
.B2(n_202),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_175),
.B1(n_174),
.B2(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_171),
.C(n_158),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_242),
.B1(n_250),
.B2(n_253),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_238),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_184),
.C(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_240),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_203),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_207),
.B1(n_196),
.B2(n_172),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_218),
.B1(n_225),
.B2(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_4),
.C(n_5),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_221),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_270),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_R g256 ( 
.A(n_252),
.B(n_221),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_224),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

BUFx12f_ASAP7_75t_SL g258 ( 
.A(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_234),
.B1(n_242),
.B2(n_236),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_233),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_216),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_237),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_223),
.B(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_237),
.C(n_211),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_267),
.C(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_284),
.B1(n_9),
.B2(n_10),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_244),
.B1(n_223),
.B2(n_238),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_222),
.B1(n_253),
.B2(n_254),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_275),
.B(n_283),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_263),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_293),
.C(n_294),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_256),
.B(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_267),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_262),
.B(n_264),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_273),
.B(n_280),
.Y(n_299)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_270),
.A3(n_255),
.B1(n_249),
.B2(n_209),
.C(n_12),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_7),
.C(n_9),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_283),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_305),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_284),
.B(n_12),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_298),
.B(n_300),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_11),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_11),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_309),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_308),
.B(n_297),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_294),
.B(n_288),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_312),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_311),
.C(n_305),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_313),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_314),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_15),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_16),
.B(n_309),
.Y(n_320)
);


endmodule