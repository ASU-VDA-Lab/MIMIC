module fake_jpeg_26213_n_250 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_20),
.B1(n_33),
.B2(n_28),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_20),
.B1(n_24),
.B2(n_12),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_33),
.B1(n_28),
.B2(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_29),
.B(n_25),
.C(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_76),
.B1(n_42),
.B2(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_77),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_27),
.B(n_35),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_33),
.B1(n_31),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_25),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_26),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_47),
.B1(n_58),
.B2(n_13),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_21),
.B1(n_15),
.B2(n_12),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_34),
.B1(n_60),
.B2(n_42),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_86),
.B1(n_75),
.B2(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_89),
.B1(n_93),
.B2(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_59),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_88),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_42),
.B1(n_19),
.B2(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_42),
.B1(n_49),
.B2(n_46),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_74),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_77),
.B1(n_70),
.B2(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_36),
.CON(n_107),
.SN(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_106),
.B1(n_115),
.B2(n_80),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_64),
.B(n_62),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_107),
.B(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_75),
.B1(n_62),
.B2(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_93),
.B1(n_91),
.B2(n_72),
.Y(n_131)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_113),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_19),
.B(n_21),
.C(n_17),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_83),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_121),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_123),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_82),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_14),
.CI(n_65),
.CON(n_141),
.SN(n_141)
);

BUFx12f_ASAP7_75t_SL g127 ( 
.A(n_110),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_135),
.B(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_45),
.B1(n_65),
.B2(n_38),
.Y(n_148)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_107),
.B1(n_64),
.B2(n_16),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_21),
.B1(n_105),
.B2(n_56),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_68),
.B1(n_66),
.B2(n_45),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_148),
.B1(n_151),
.B2(n_40),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_65),
.B(n_1),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_143),
.B(n_149),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_32),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_68),
.C(n_38),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_155),
.C(n_157),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_23),
.B(n_10),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_54),
.B1(n_38),
.B2(n_24),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_38),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_26),
.C(n_30),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_26),
.C(n_30),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_166),
.C(n_174),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_163),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_133),
.C(n_30),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_151),
.B1(n_137),
.B2(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_26),
.C(n_30),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_184),
.B1(n_187),
.B2(n_183),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_187),
.B1(n_173),
.B2(n_174),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_140),
.B(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_190),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_150),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_193),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_157),
.B1(n_158),
.B2(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_146),
.C(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_160),
.C(n_168),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_148),
.B(n_139),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_141),
.B1(n_40),
.B2(n_24),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_30),
.B1(n_32),
.B2(n_8),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_8),
.B(n_10),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_162),
.B1(n_170),
.B2(n_171),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_195),
.B1(n_206),
.B2(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_180),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_165),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_1),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_185),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_169),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_32),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_178),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_215),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_212),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_196),
.A2(n_193),
.B1(n_9),
.B2(n_10),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_201),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_23),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_225),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_36),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_197),
.B(n_205),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_1),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_22),
.C(n_36),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_36),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_213),
.C(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_232),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_221),
.B(n_4),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_22),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_36),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_234),
.B1(n_23),
.B2(n_5),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_241),
.B(n_236),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_5),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_2),
.B(n_4),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_22),
.C(n_6),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_6),
.B(n_7),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_247),
.A2(n_6),
.B(n_7),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_6),
.B(n_7),
.Y(n_249)
);

OAI22x1_ASAP7_75t_SL g250 ( 
.A1(n_249),
.A2(n_22),
.B1(n_232),
.B2(n_127),
.Y(n_250)
);


endmodule