module fake_aes_1912_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_5), .B(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_16), .B(n_0), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
OAI22xp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_12), .B1(n_17), .B2(n_14), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_12), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_13), .B1(n_15), .B2(n_3), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_13), .B1(n_2), .B2(n_7), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_24), .B(n_20), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_24), .B(n_21), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_21), .B1(n_18), .B2(n_13), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_27), .B(n_23), .Y(n_31) );
NAND2x1_ASAP7_75t_L g32 ( .A(n_30), .B(n_13), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_30), .B(n_29), .Y(n_34) );
NOR2xp33_ASAP7_75t_L g35 ( .A(n_33), .B(n_1), .Y(n_35) );
AOI221xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_22), .B1(n_2), .B2(n_7), .C(n_1), .Y(n_36) );
NOR3x1_ASAP7_75t_L g37 ( .A(n_32), .B(n_8), .C(n_9), .Y(n_37) );
OAI211xp5_ASAP7_75t_SL g38 ( .A1(n_35), .A2(n_10), .B(n_22), .C(n_36), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
AOI22xp5_ASAP7_75t_SL g41 ( .A1(n_40), .A2(n_22), .B1(n_39), .B2(n_12), .Y(n_41) );
endmodule