module fake_netlist_6_2772_n_2439 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2439);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2439;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_161),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_48),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_62),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_112),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_136),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_132),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_72),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_230),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_60),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_48),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_150),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_113),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_107),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_164),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_72),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_126),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_90),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_70),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_101),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_180),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_96),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_212),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_116),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_148),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_69),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_46),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_82),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_170),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_73),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_114),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_124),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_144),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_142),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_156),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_105),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_87),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_94),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_78),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_77),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_81),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_17),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_127),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_82),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_215),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_27),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_204),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_78),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_200),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_22),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_4),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_10),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_73),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_47),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_211),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_60),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_192),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_4),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_37),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_65),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_121),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_160),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_94),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_55),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_146),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_19),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_130),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_188),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_213),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_185),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_206),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_183),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_133),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_31),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_22),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_77),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_59),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_10),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_25),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_104),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_91),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_97),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_85),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_147),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_63),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_69),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_87),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_172),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_43),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_153),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_201),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_75),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_208),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_131),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_117),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_125),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_207),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_157),
.Y(n_379)
);

BUFx2_ASAP7_75t_SL g380 ( 
.A(n_220),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_53),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_56),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_49),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_23),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_44),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_30),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_97),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_137),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_186),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_166),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_179),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_225),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_120),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_139),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_65),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_50),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_81),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_59),
.Y(n_399)
);

BUFx2_ASAP7_75t_SL g400 ( 
.A(n_99),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_18),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_67),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_57),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_96),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_174),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_39),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_227),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_30),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_216),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_15),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_51),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_71),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_119),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_49),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_224),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_95),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_9),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_63),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_154),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_64),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_98),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_167),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_1),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_3),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_31),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_223),
.Y(n_426)
);

BUFx10_ASAP7_75t_L g427 ( 
.A(n_86),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_54),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_85),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_38),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_46),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_11),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_228),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_25),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_66),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_47),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_42),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_50),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_169),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_7),
.Y(n_440)
);

BUFx2_ASAP7_75t_SL g441 ( 
.A(n_58),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_163),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_33),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_67),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_75),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_13),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_1),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_52),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_68),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_110),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_38),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_165),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_103),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_40),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_18),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_20),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_118),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_425),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_246),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_246),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_234),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_246),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_243),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_246),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_246),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_259),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_246),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_246),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_246),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_236),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_246),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_261),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_427),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_323),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_0),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_331),
.B(n_0),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_331),
.B(n_2),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_290),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_301),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_323),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_271),
.B(n_2),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_242),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_343),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_254),
.B(n_5),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_251),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_345),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_323),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_323),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_252),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_323),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_235),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_260),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_347),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_247),
.B(n_6),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_373),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_269),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_388),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_254),
.B(n_6),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_322),
.B(n_9),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_275),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_235),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_302),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_237),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_237),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_238),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_286),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_238),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_247),
.B(n_11),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_258),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_389),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_393),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_258),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_264),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_264),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_418),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_288),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_233),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_272),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_439),
.B(n_12),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_272),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_239),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_294),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_273),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_305),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_309),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_273),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_282),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_317),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_282),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_291),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_291),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_439),
.B(n_12),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_240),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_296),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_321),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_427),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_296),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_303),
.B(n_13),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_324),
.Y(n_544)
);

INVxp33_ASAP7_75t_SL g545 ( 
.A(n_325),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_303),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_327),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_304),
.B(n_14),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_328),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_304),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_333),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_265),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_265),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_334),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_335),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_338),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_267),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_297),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_241),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_267),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_435),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_281),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_306),
.B(n_14),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_281),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_292),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_306),
.B(n_16),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_339),
.Y(n_569)
);

INVxp33_ASAP7_75t_SL g570 ( 
.A(n_341),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_244),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_329),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_292),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_308),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_308),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_348),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_315),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_350),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_352),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_315),
.B(n_16),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_245),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_458),
.B(n_255),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_506),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_521),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_475),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_525),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_538),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_563),
.B(n_476),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_561),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_459),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_571),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_581),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_289),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_461),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_489),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_471),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_471),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_484),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_476),
.B(n_435),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_484),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_490),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_487),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_512),
.B(n_248),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_506),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_482),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_532),
.Y(n_616)
);

INVx6_ASAP7_75t_L g617 ( 
.A(n_553),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_492),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_487),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_494),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_499),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_553),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_470),
.B(n_254),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_486),
.B(n_289),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_464),
.B(n_255),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_491),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_491),
.Y(n_632)
);

CKINVDCx8_ASAP7_75t_R g633 ( 
.A(n_474),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_495),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_495),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_463),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_256),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_500),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_462),
.Y(n_641)
);

OA21x2_ASAP7_75t_L g642 ( 
.A1(n_470),
.A2(n_337),
.B(n_318),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_465),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_466),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_537),
.B(n_257),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_553),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_468),
.B(n_262),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_502),
.B(n_344),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_500),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_467),
.B(n_250),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_469),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_472),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_472),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_504),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_493),
.B(n_263),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_560),
.B(n_268),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_473),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_554),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_572),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_505),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_483),
.A2(n_310),
.B1(n_319),
.B2(n_287),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_555),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_559),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_562),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_510),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_479),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_507),
.B(n_445),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_508),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_520),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_562),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_520),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_649),
.B(n_344),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_526),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_647),
.B(n_545),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_625),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_624),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_678),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_626),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_611),
.B(n_570),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_626),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_653),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_557),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_649),
.B(n_344),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_591),
.B(n_441),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_653),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_656),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_624),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_611),
.B(n_529),
.Y(n_695)
);

CKINVDCx14_ASAP7_75t_R g696 ( 
.A(n_658),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_656),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_591),
.B(n_441),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_R g699 ( 
.A(n_586),
.B(n_480),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_654),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_624),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_589),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_627),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_593),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_584),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_584),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_584),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_593),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_607),
.B(n_509),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_593),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_584),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_646),
.B(n_541),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_641),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_585),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_646),
.B(n_529),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_638),
.B(n_533),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_626),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_594),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_583),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_594),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_646),
.B(n_533),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_607),
.B(n_511),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_638),
.B(n_544),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_617),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_642),
.B(n_318),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_585),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_590),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_594),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_645),
.B(n_513),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_641),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_625),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_583),
.Y(n_736)
);

BUFx4f_ASAP7_75t_L g737 ( 
.A(n_642),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_585),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_516),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_585),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_585),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_644),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_649),
.A2(n_478),
.B1(n_477),
.B2(n_642),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_585),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_648),
.B(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_646),
.B(n_544),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_582),
.A2(n_503),
.B1(n_519),
.B2(n_497),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_630),
.A2(n_549),
.B1(n_552),
.B2(n_547),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_644),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_648),
.B(n_518),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_666),
.B(n_657),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_598),
.Y(n_753)
);

NAND2x1_ASAP7_75t_L g754 ( 
.A(n_625),
.B(n_302),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_652),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_652),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_598),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_598),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_617),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_617),
.Y(n_760)
);

CKINVDCx8_ASAP7_75t_R g761 ( 
.A(n_592),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_627),
.B(n_522),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_649),
.A2(n_543),
.B1(n_565),
.B2(n_548),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_652),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_657),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_674),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_588),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_617),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_665),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_666),
.B(n_481),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_614),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_626),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_626),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_627),
.B(n_524),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_588),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_614),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_617),
.B(n_527),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_674),
.B(n_660),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_600),
.B(n_547),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_610),
.A2(n_552),
.B1(n_556),
.B2(n_549),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_622),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_640),
.B(n_483),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_665),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_665),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_640),
.B(n_556),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_605),
.B(n_558),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_635),
.A2(n_266),
.B1(n_330),
.B2(n_249),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_626),
.B(n_530),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_643),
.B(n_531),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_534),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_655),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_662),
.B(n_535),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_642),
.A2(n_580),
.B1(n_568),
.B2(n_625),
.Y(n_795)
);

BUFx10_ASAP7_75t_L g796 ( 
.A(n_606),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_655),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_622),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_655),
.Y(n_799)
);

INVx4_ASAP7_75t_SL g800 ( 
.A(n_625),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_588),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_622),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_664),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_659),
.B(n_558),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_625),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_664),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_588),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_663),
.B(n_380),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_619),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_631),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_664),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_632),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_665),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_569),
.Y(n_816)
);

INVx8_ASAP7_75t_L g817 ( 
.A(n_625),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_650),
.B(n_569),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_662),
.B(n_536),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_665),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_588),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_643),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_588),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_672),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_675),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_676),
.B(n_576),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_675),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_651),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_643),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_651),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_625),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_643),
.B(n_539),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_595),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_612),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_587),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_675),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_675),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_675),
.B(n_576),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_587),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_675),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_735),
.B(n_329),
.Y(n_841)
);

O2A1O1Ixp5_ASAP7_75t_L g842 ( 
.A1(n_737),
.A2(n_546),
.B(n_550),
.C(n_542),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_695),
.B(n_633),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_726),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_720),
.B(n_633),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_726),
.B(n_578),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_765),
.B(n_643),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_710),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_691),
.B(n_380),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_835),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_727),
.B(n_733),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_739),
.B(n_643),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_710),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_693),
.B(n_596),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_746),
.B(n_578),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_835),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_779),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_751),
.B(n_579),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_703),
.B(n_579),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_712),
.B(n_667),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_599),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_822),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_686),
.B(n_688),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_839),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_599),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_839),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_779),
.B(n_337),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_697),
.B(n_314),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_795),
.A2(n_379),
.B1(n_378),
.B2(n_349),
.Y(n_870)
);

AND2x6_ASAP7_75t_SL g871 ( 
.A(n_780),
.B(n_271),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_743),
.A2(n_379),
.B1(n_378),
.B2(n_349),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_700),
.B(n_838),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_779),
.B(n_368),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_775),
.B(n_601),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_680),
.B(n_485),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_775),
.B(n_601),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_683),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_775),
.A2(n_488),
.B1(n_498),
.B2(n_496),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_691),
.B(n_400),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_681),
.B(n_501),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_793),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_712),
.B(n_340),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_712),
.B(n_667),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_793),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_689),
.B(n_514),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_705),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_762),
.B(n_602),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_767),
.B(n_667),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_689),
.B(n_515),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_705),
.Y(n_891)
);

BUFx4f_ASAP7_75t_L g892 ( 
.A(n_679),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_711),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_788),
.B(n_637),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_711),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_797),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_778),
.B(n_602),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_748),
.B(n_270),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_763),
.B(n_603),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_774),
.B(n_603),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_829),
.B(n_609),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_737),
.B(n_609),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_683),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_752),
.A2(n_442),
.B1(n_276),
.B2(n_279),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_749),
.B(n_274),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_752),
.B(n_283),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_713),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_713),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_679),
.A2(n_362),
.B1(n_377),
.B2(n_340),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_679),
.A2(n_690),
.B1(n_737),
.B2(n_729),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_699),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_728),
.B(n_615),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_816),
.B(n_661),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_679),
.A2(n_377),
.B1(n_391),
.B2(n_362),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_826),
.B(n_673),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_SL g916 ( 
.A(n_781),
.B(n_385),
.C(n_360),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_735),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_719),
.B(n_399),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_722),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_784),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_694),
.B(n_701),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_735),
.B(n_329),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_723),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_728),
.B(n_759),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_797),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_725),
.B(n_747),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_691),
.A2(n_293),
.B1(n_295),
.B2(n_284),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_714),
.A2(n_391),
.B(n_457),
.C(n_395),
.Y(n_928)
);

NOR2x1p5_ASAP7_75t_L g929 ( 
.A(n_771),
.B(n_445),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_722),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_R g931 ( 
.A(n_696),
.B(n_298),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_691),
.A2(n_300),
.B1(n_316),
.B2(n_299),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_698),
.A2(n_784),
.B1(n_809),
.B2(n_701),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_799),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_702),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_724),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_724),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_759),
.B(n_615),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_760),
.B(n_618),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_694),
.B(n_395),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_354),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_732),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_805),
.B(n_355),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_792),
.B(n_667),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_698),
.B(n_400),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_723),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_799),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_760),
.B(n_618),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_787),
.B(n_320),
.Y(n_949)
);

INVx8_ASAP7_75t_L g950 ( 
.A(n_735),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_769),
.B(n_620),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_787),
.B(n_336),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_732),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_804),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_736),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_769),
.B(n_620),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_679),
.B(n_621),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_736),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_753),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_804),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_716),
.B(n_342),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_698),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_679),
.B(n_621),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_690),
.B(n_790),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_690),
.A2(n_457),
.B1(n_302),
.B2(n_329),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_792),
.B(n_668),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_690),
.B(n_791),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_807),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_811),
.B(n_813),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_690),
.B(n_623),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_698),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_761),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_811),
.B(n_346),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_690),
.A2(n_729),
.B1(n_742),
.B2(n_734),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_807),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_832),
.B(n_623),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_822),
.B(n_628),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_818),
.B(n_356),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_809),
.A2(n_419),
.B1(n_426),
.B2(n_415),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_729),
.B(n_628),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_714),
.B(n_629),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_717),
.B(n_629),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_813),
.B(n_357),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_754),
.B(n_302),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_704),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_717),
.A2(n_577),
.B(n_636),
.C(n_253),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_764),
.B(n_744),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_753),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_682),
.B(n_358),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_757),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_784),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_764),
.B(n_636),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_682),
.B(n_366),
.Y(n_993)
);

OAI221xp5_ASAP7_75t_L g994 ( 
.A1(n_771),
.A2(n_253),
.B1(n_421),
.B2(n_429),
.C(n_332),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_757),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_750),
.A2(n_302),
.B1(n_329),
.B2(n_376),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_755),
.B(n_616),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_830),
.B(n_421),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_756),
.B(n_616),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_800),
.B(n_277),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_812),
.A2(n_329),
.B1(n_376),
.B2(n_429),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_794),
.B(n_616),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_794),
.B(n_616),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_682),
.B(n_668),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_682),
.B(n_670),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_812),
.A2(n_329),
.B1(n_376),
.B2(n_396),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_818),
.B(n_361),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_828),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_819),
.B(n_616),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_809),
.B(n_801),
.Y(n_1010)
);

AND2x2_ASAP7_75t_SL g1011 ( 
.A(n_801),
.B(n_396),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_809),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_819),
.B(n_616),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_704),
.B(n_669),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_704),
.B(n_669),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_921),
.Y(n_1016)
);

NAND2x1p5_ASAP7_75t_L g1017 ( 
.A(n_917),
.B(n_682),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_851),
.B(n_706),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_918),
.B(n_810),
.C(n_731),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_955),
.B(n_810),
.Y(n_1020)
);

BUFx12f_ASAP7_75t_L g1021 ( 
.A(n_935),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_923),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_856),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_846),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_857),
.B(n_921),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_873),
.B(n_706),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_864),
.B(n_696),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_863),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_985),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_856),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_944),
.B(n_706),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_966),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_878),
.Y(n_1034)
);

AND3x1_ASAP7_75t_SL g1035 ( 
.A(n_929),
.B(n_994),
.C(n_278),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_865),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_958),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_862),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_SL g1039 ( 
.A(n_870),
.B(n_702),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_944),
.B(n_708),
.Y(n_1040)
);

AND2x2_ASAP7_75t_SL g1041 ( 
.A(n_872),
.B(n_397),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_857),
.B(n_800),
.Y(n_1042)
);

AOI211xp5_ASAP7_75t_L g1043 ( 
.A1(n_941),
.A2(n_789),
.B(n_833),
.C(n_731),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_848),
.B(n_708),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_848),
.B(n_708),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_846),
.B(n_684),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_865),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_917),
.B(n_806),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_920),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_917),
.B(n_806),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_921),
.B(n_800),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_916),
.B(n_365),
.C(n_363),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_853),
.B(n_718),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_966),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_985),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_935),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_855),
.B(n_684),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_858),
.B(n_1011),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_878),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_899),
.A2(n_277),
.B1(n_280),
.B2(n_278),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_850),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_850),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_972),
.B(n_420),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_950),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_911),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_853),
.B(n_718),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_903),
.B(n_800),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_862),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_950),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_998),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_847),
.A2(n_817),
.B(n_806),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_903),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_911),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1011),
.B(n_684),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_882),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_889),
.B(n_718),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_844),
.B(n_783),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_867),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_882),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_730),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_860),
.B(n_730),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_972),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_867),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_962),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_931),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_917),
.B(n_806),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1010),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_860),
.B(n_670),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_998),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_844),
.B(n_943),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_884),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_884),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_978),
.B(n_783),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_885),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_962),
.B(n_671),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1007),
.B(n_783),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_892),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_854),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_971),
.B(n_817),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_890),
.B(n_383),
.C(n_382),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_985),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_896),
.Y(n_1103)
);

BUFx4f_ASAP7_75t_L g1104 ( 
.A(n_971),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_896),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_925),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_SL g1107 ( 
.A(n_876),
.B(n_761),
.Y(n_1107)
);

NAND2x1_ASAP7_75t_L g1108 ( 
.A(n_907),
.B(n_730),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_869),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_925),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_886),
.B(n_796),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1010),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_871),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_934),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_907),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_934),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_917),
.A2(n_817),
.B(n_806),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_892),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_849),
.B(n_880),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_879),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_950),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_950),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_947),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_849),
.B(n_817),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_852),
.B(n_745),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_926),
.B(n_745),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_910),
.B(n_831),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_894),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_888),
.B(n_745),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_974),
.A2(n_831),
.B1(n_754),
.B2(n_833),
.Y(n_1130)
);

AND3x1_ASAP7_75t_SL g1131 ( 
.A(n_929),
.B(n_285),
.C(n_280),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_SL g1132 ( 
.A(n_1010),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_947),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_954),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_892),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_913),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_906),
.A2(n_417),
.B(n_397),
.C(n_312),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_915),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_969),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1010),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_875),
.A2(n_840),
.B1(n_837),
.B2(n_836),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_954),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_868),
.B(n_834),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_960),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_964),
.B(n_831),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_868),
.B(n_834),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_960),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_868),
.B(n_877),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_991),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_883),
.B(n_834),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_991),
.B(n_671),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_907),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_883),
.B(n_821),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_940),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_967),
.B(n_831),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_SL g1157 ( 
.A(n_949),
.B(n_386),
.C(n_384),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_902),
.A2(n_332),
.B1(n_440),
.B2(n_326),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_968),
.Y(n_1159)
);

AOI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_881),
.A2(n_437),
.B1(n_845),
.B2(n_843),
.C1(n_1008),
.C2(n_898),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_975),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_1002),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_R g1163 ( 
.A(n_849),
.B(n_398),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_975),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1003),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_924),
.A2(n_831),
.B(n_687),
.Y(n_1166)
);

BUFx8_ASAP7_75t_SL g1167 ( 
.A(n_849),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1009),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_880),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_859),
.A2(n_827),
.B1(n_825),
.B2(n_770),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_883),
.B(n_821),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_940),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_887),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1013),
.B(n_821),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_880),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_952),
.B(n_796),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_887),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_940),
.Y(n_1178)
);

OR2x4_ASAP7_75t_L g1179 ( 
.A(n_866),
.B(n_285),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_957),
.B(n_785),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_891),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_897),
.B(n_786),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_891),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_893),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_880),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1012),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_904),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_SL g1188 ( 
.A(n_933),
.B(n_404),
.C(n_401),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_893),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_945),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_945),
.B(n_814),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_895),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_874),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_895),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1000),
.Y(n_1195)
);

AND3x2_ASAP7_75t_L g1196 ( 
.A(n_945),
.B(n_312),
.C(n_311),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_SL g1197 ( 
.A(n_905),
.B(n_408),
.C(n_406),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_908),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_909),
.A2(n_432),
.B1(n_351),
.B2(n_326),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_908),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_945),
.B(n_815),
.Y(n_1201)
);

BUFx4_ASAP7_75t_SL g1202 ( 
.A(n_973),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_983),
.B(n_796),
.Y(n_1203)
);

BUFx5_ASAP7_75t_L g1204 ( 
.A(n_1000),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1000),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_919),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_927),
.B(n_824),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1000),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_SL g1209 ( 
.A1(n_979),
.A2(n_423),
.B1(n_412),
.B2(n_414),
.Y(n_1209)
);

OR2x2_ASAP7_75t_SL g1210 ( 
.A(n_961),
.B(n_311),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_919),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1020),
.B(n_932),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1051),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1033),
.B(n_976),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1166),
.A2(n_842),
.B(n_987),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1058),
.A2(n_980),
.B1(n_861),
.B2(n_914),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1046),
.B(n_824),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1051),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1058),
.A2(n_963),
.B1(n_970),
.B2(n_824),
.Y(n_1219)
);

NAND2x1_ASAP7_75t_L g1220 ( 
.A(n_1064),
.B(n_930),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_L g1221 ( 
.A1(n_1126),
.A2(n_938),
.B(n_939),
.C(n_912),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_SL g1222 ( 
.A1(n_1135),
.A2(n_951),
.B(n_948),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1070),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1162),
.A2(n_922),
.B(n_841),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1022),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1044),
.A2(n_1015),
.B(n_1014),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1045),
.A2(n_977),
.B(n_997),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1075),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1065),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1089),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1127),
.A2(n_922),
.B(n_841),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_999),
.B(n_936),
.Y(n_1232)
);

OAI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_1057),
.A2(n_430),
.B(n_424),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1032),
.A2(n_901),
.B(n_900),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1033),
.A2(n_687),
.A3(n_773),
.B1(n_721),
.B2(n_685),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1079),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_1124),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1066),
.A2(n_936),
.B(n_930),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1145),
.A2(n_956),
.B(n_981),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1054),
.B(n_937),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1024),
.B(n_982),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1127),
.A2(n_1018),
.B(n_1148),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1145),
.A2(n_992),
.B(n_989),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1039),
.A2(n_965),
.B(n_937),
.C(n_942),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1054),
.B(n_942),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_959),
.B(n_953),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1125),
.A2(n_820),
.B(n_953),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1114),
.A2(n_928),
.A3(n_986),
.B(n_959),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1136),
.B(n_988),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1111),
.B(n_297),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1114),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1030),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1071),
.A2(n_1005),
.B(n_1004),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1136),
.B(n_988),
.Y(n_1254)
);

O2A1O1Ixp5_ASAP7_75t_L g1255 ( 
.A1(n_1156),
.A2(n_990),
.B(n_995),
.C(n_993),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1090),
.B(n_990),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1132),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1055),
.A2(n_995),
.B(n_984),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1055),
.A2(n_984),
.B(n_1004),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_687),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1055),
.A2(n_984),
.B(n_1006),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1051),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1037),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1040),
.A2(n_1000),
.B(n_1001),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1102),
.A2(n_766),
.B(n_758),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1120),
.A2(n_359),
.B1(n_455),
.B2(n_313),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1165),
.B(n_1000),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1168),
.B(n_1091),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1076),
.A2(n_996),
.B(n_766),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1116),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1038),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1042),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1102),
.A2(n_772),
.B(n_758),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1107),
.B(n_369),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1156),
.A2(n_721),
.B(n_685),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1016),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1102),
.A2(n_777),
.B(n_772),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1129),
.A2(n_721),
.B(n_685),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1182),
.A2(n_773),
.B(n_709),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1116),
.A2(n_1161),
.B(n_1159),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1173),
.A2(n_782),
.B(n_777),
.Y(n_1282)
);

NOR2xp67_ASAP7_75t_SL g1283 ( 
.A(n_1097),
.B(n_370),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1159),
.A2(n_803),
.A3(n_798),
.B(n_782),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1065),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1170),
.A2(n_803),
.B(n_798),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1178),
.A2(n_773),
.B1(n_433),
.B2(n_450),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1057),
.B(n_371),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1082),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1135),
.A2(n_823),
.B(n_709),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1092),
.B(n_1088),
.Y(n_1291)
);

AO22x2_ASAP7_75t_L g1292 ( 
.A1(n_1019),
.A2(n_411),
.B1(n_364),
.B2(n_359),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1173),
.A2(n_677),
.B(n_669),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1039),
.A2(n_351),
.B(n_313),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1088),
.B(n_677),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1034),
.B(n_564),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1178),
.A2(n_374),
.B1(n_452),
.B2(n_413),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1173),
.A2(n_677),
.B(n_566),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1207),
.A2(n_440),
.B(n_402),
.C(n_403),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1160),
.B(n_434),
.C(n_431),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1088),
.B(n_375),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1183),
.A2(n_564),
.B(n_566),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1161),
.A2(n_416),
.A3(n_353),
.B(n_364),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1016),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1094),
.Y(n_1305)
);

OA22x2_ASAP7_75t_L g1306 ( 
.A1(n_1193),
.A2(n_387),
.B1(n_381),
.B2(n_372),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1081),
.A2(n_823),
.B(n_808),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_SL g1308 ( 
.A1(n_1023),
.A2(n_387),
.B(n_381),
.C(n_455),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1021),
.B(n_255),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1027),
.B(n_297),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1027),
.B(n_390),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1138),
.B(n_436),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1056),
.B(n_567),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1080),
.A2(n_823),
.B(n_808),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1143),
.A2(n_823),
.B(n_808),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1183),
.A2(n_573),
.B(n_574),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1043),
.B(n_447),
.C(n_446),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1146),
.A2(n_823),
.B(n_808),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1028),
.A2(n_394),
.B1(n_453),
.B2(n_409),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1016),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1060),
.A2(n_448),
.B1(n_444),
.B2(n_353),
.C(n_432),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1034),
.B(n_567),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1128),
.B(n_438),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1207),
.A2(n_444),
.B(n_372),
.C(n_448),
.Y(n_1324)
);

NOR2x1_ASAP7_75t_SL g1325 ( 
.A(n_1124),
.B(n_707),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1172),
.B(n_392),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1082),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1098),
.Y(n_1328)
);

NAND2x1_ASAP7_75t_L g1329 ( 
.A(n_1064),
.B(n_707),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_808),
.B(n_802),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1031),
.A2(n_575),
.B(n_573),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1052),
.B(n_451),
.C(n_456),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1183),
.A2(n_575),
.B(n_574),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1041),
.B(n_405),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1103),
.A2(n_411),
.B(n_402),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1021),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1153),
.A2(n_802),
.B(n_776),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1171),
.A2(n_1041),
.B(n_1130),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1189),
.Y(n_1339)
);

BUFx5_ASAP7_75t_L g1340 ( 
.A(n_1180),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1061),
.A2(n_407),
.B(n_403),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1117),
.A2(n_802),
.B(n_776),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1105),
.A2(n_416),
.A3(n_417),
.B(n_329),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1106),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1064),
.B(n_707),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1189),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1025),
.B(n_443),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1128),
.B(n_449),
.Y(n_1348)
);

NOR4xp25_ASAP7_75t_L g1349 ( 
.A(n_1137),
.B(n_297),
.C(n_307),
.D(n_367),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1074),
.B(n_802),
.C(n_776),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1135),
.A2(n_123),
.B(n_102),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1189),
.A2(n_802),
.B(n_776),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1049),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1073),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1029),
.A2(n_776),
.B(n_768),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1110),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1061),
.A2(n_768),
.B(n_741),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1017),
.A2(n_1050),
.B(n_1048),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1085),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1016),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1186),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1025),
.B(n_707),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1115),
.A2(n_768),
.B(n_741),
.Y(n_1363)
);

AND2x6_ASAP7_75t_L g1364 ( 
.A(n_1097),
.B(n_707),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1123),
.A2(n_768),
.B(n_741),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1186),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1025),
.B(n_709),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1017),
.A2(n_768),
.B(n_741),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1048),
.A2(n_741),
.B(n_740),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1133),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1072),
.B(n_108),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_R g1372 ( 
.A(n_1073),
.B(n_115),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1097),
.B(n_709),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1077),
.B(n_307),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1115),
.A2(n_1152),
.B(n_1062),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1115),
.A2(n_1152),
.B(n_1062),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1042),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1134),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1142),
.A2(n_740),
.B1(n_738),
.B2(n_715),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1223),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1238),
.A2(n_1108),
.B(n_1194),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1246),
.A2(n_1198),
.B(n_1194),
.Y(n_1382)
);

OR2x2_ASAP7_75t_SL g1383 ( 
.A(n_1300),
.B(n_1149),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1212),
.A2(n_1187),
.B1(n_1074),
.B2(n_1209),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1223),
.Y(n_1385)
);

OAI211xp5_ASAP7_75t_L g1386 ( 
.A1(n_1233),
.A2(n_1060),
.B(n_1187),
.C(n_1109),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1221),
.A2(n_1147),
.B(n_1144),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1237),
.B(n_1069),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1252),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1242),
.B(n_1119),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1221),
.A2(n_1164),
.B(n_1155),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1242),
.A2(n_1047),
.B(n_1036),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1229),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1215),
.A2(n_1083),
.B(n_1078),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1272),
.B(n_1228),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1375),
.A2(n_1200),
.B(n_1198),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1271),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1376),
.A2(n_1232),
.B(n_1352),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1312),
.A2(n_1099),
.B1(n_1063),
.B2(n_1101),
.C(n_1163),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1222),
.A2(n_1141),
.B(n_1188),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1255),
.A2(n_1181),
.B(n_1177),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1281),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1237),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1231),
.B(n_1119),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1281),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1323),
.B(n_1085),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1284),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1257),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1258),
.A2(n_1200),
.B(n_1152),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1284),
.Y(n_1410)
);

AOI22x1_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1211),
.B1(n_1192),
.B2(n_1184),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1294),
.A2(n_1112),
.B1(n_1140),
.B2(n_1087),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_SL g1413 ( 
.A(n_1237),
.B(n_1097),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1241),
.A2(n_1035),
.B1(n_1176),
.B2(n_1139),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1284),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1255),
.A2(n_1206),
.B(n_1158),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1271),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1230),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1338),
.A2(n_1197),
.B(n_1157),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1241),
.B(n_1203),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1361),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1249),
.B(n_1158),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1284),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1262),
.B(n_1154),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1363),
.A2(n_1050),
.B(n_1086),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1224),
.A2(n_1208),
.B(n_1086),
.Y(n_1426)
);

NAND2x1_ASAP7_75t_L g1427 ( 
.A(n_1290),
.B(n_1069),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1231),
.A2(n_1095),
.B(n_1151),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1234),
.A2(n_1095),
.B(n_1151),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1299),
.A2(n_1190),
.B(n_1068),
.C(n_1175),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1359),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1285),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1309),
.A2(n_1163),
.B1(n_1348),
.B2(n_1323),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1293),
.A2(n_1199),
.B(n_1180),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1370),
.A2(n_1154),
.B1(n_1104),
.B2(n_1119),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1341),
.A2(n_1104),
.B(n_1095),
.C(n_1151),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1265),
.A2(n_1199),
.B(n_1180),
.Y(n_1437)
);

CKINVDCx6p67_ASAP7_75t_R g1438 ( 
.A(n_1336),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1236),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1354),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1274),
.A2(n_1180),
.B(n_1204),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1213),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1278),
.A2(n_1180),
.B(n_1204),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1317),
.A2(n_1185),
.B1(n_1132),
.B2(n_1119),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1298),
.A2(n_1204),
.B(n_1104),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1230),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1251),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1325),
.A2(n_1122),
.B(n_1069),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1253),
.A2(n_1208),
.B(n_1122),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1249),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1227),
.A2(n_1201),
.B(n_1191),
.Y(n_1451)
);

NAND2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1237),
.B(n_1121),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1213),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1312),
.A2(n_1348),
.B1(n_1324),
.B2(n_1250),
.C(n_1310),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1256),
.B(n_1210),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1213),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1282),
.A2(n_1204),
.B(n_1122),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1302),
.A2(n_1201),
.B(n_1191),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1286),
.A2(n_1191),
.B(n_1201),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1262),
.B(n_1067),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1213),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1268),
.B(n_1084),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1270),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1316),
.A2(n_1169),
.B(n_1042),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1286),
.A2(n_1067),
.B(n_1179),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1333),
.A2(n_1169),
.B(n_1179),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1225),
.B(n_1072),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1218),
.Y(n_1468)
);

CKINVDCx8_ASAP7_75t_R g1469 ( 
.A(n_1371),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1370),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1226),
.A2(n_1204),
.B(n_1121),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1305),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1253),
.A2(n_1208),
.B(n_1121),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1321),
.A2(n_1067),
.B(n_1131),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1254),
.A2(n_1118),
.B1(n_1059),
.B2(n_1084),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1339),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1346),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1342),
.A2(n_1204),
.B(n_1100),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1342),
.A2(n_1204),
.B(n_1100),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1254),
.B(n_1059),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1216),
.A2(n_1124),
.B(n_1100),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1214),
.B(n_1059),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_SL g1483 ( 
.A1(n_1351),
.A2(n_1132),
.B(n_1190),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1264),
.A2(n_1124),
.B(n_1118),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1334),
.B(n_1059),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1244),
.A2(n_1196),
.A3(n_1100),
.B(n_376),
.Y(n_1486)
);

CKINVDCx6p67_ASAP7_75t_R g1487 ( 
.A(n_1263),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1314),
.A2(n_1118),
.B(n_1205),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1257),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1218),
.B(n_1118),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1218),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1372),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1328),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1314),
.A2(n_1205),
.B(n_1195),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1219),
.A2(n_1205),
.B(n_1195),
.C(n_1202),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1296),
.A2(n_1167),
.B1(n_422),
.B2(n_1205),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1291),
.B(n_1195),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1239),
.A2(n_1195),
.B(n_329),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1344),
.Y(n_1499)
);

CKINVDCx6p67_ASAP7_75t_R g1500 ( 
.A(n_1327),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1311),
.B(n_1167),
.Y(n_1501)
);

AOI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1243),
.A2(n_740),
.B(n_738),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1292),
.A2(n_1266),
.B1(n_1349),
.B2(n_1332),
.C(n_1374),
.Y(n_1503)
);

CKINVDCx6p67_ASAP7_75t_R g1504 ( 
.A(n_1217),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1356),
.A2(n_1113),
.B1(n_740),
.B2(n_738),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1353),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1378),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1240),
.Y(n_1508)
);

AO21x1_ASAP7_75t_L g1509 ( 
.A1(n_1373),
.A2(n_376),
.B(n_422),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1245),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1248),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1218),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1267),
.A2(n_376),
.B(n_422),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_SL g1514 ( 
.A1(n_1373),
.A2(n_376),
.B(n_226),
.C(n_221),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1296),
.A2(n_1113),
.B1(n_307),
.B2(n_454),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1273),
.B(n_307),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1248),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1273),
.B(n_1377),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1288),
.B(n_1313),
.C(n_1347),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1307),
.A2(n_376),
.B(n_738),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1295),
.B(n_17),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1307),
.A2(n_376),
.B(n_715),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1248),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1276),
.A2(n_715),
.B(n_709),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_SL g1525 ( 
.A1(n_1358),
.A2(n_218),
.B(n_214),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1357),
.A2(n_715),
.B(n_210),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1322),
.B(n_367),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1350),
.A2(n_715),
.B(n_205),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1322),
.A2(n_454),
.B1(n_367),
.B2(n_613),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1301),
.B(n_367),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1275),
.A2(n_454),
.B(n_21),
.C(n_24),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1248),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1364),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1303),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1292),
.A2(n_454),
.B1(n_613),
.B2(n_612),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1331),
.A2(n_613),
.B(n_612),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1303),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1326),
.B(n_19),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1279),
.A2(n_203),
.B(n_196),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1377),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1360),
.B(n_162),
.Y(n_1541)
);

BUFx2_ASAP7_75t_R g1542 ( 
.A(n_1362),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1247),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1366),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1277),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1247),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1292),
.A2(n_613),
.B1(n_612),
.B2(n_26),
.Y(n_1547)
);

CKINVDCx16_ASAP7_75t_R g1548 ( 
.A(n_1372),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1365),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1276),
.A2(n_173),
.B(n_134),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1277),
.Y(n_1551)
);

AOI22x1_ASAP7_75t_L g1552 ( 
.A1(n_1280),
.A2(n_613),
.B1(n_612),
.B2(n_26),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1289),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1371),
.A2(n_613),
.B1(n_612),
.B2(n_27),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1319),
.A2(n_21),
.B1(n_24),
.B2(n_28),
.Y(n_1555)
);

BUFx2_ASAP7_75t_SL g1556 ( 
.A(n_1364),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1260),
.A2(n_195),
.B(n_194),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1358),
.A2(n_193),
.B(n_190),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1269),
.A2(n_182),
.B(n_178),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1303),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1277),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1277),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1306),
.B(n_176),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1493),
.Y(n_1564)
);

NAND2xp33_ASAP7_75t_R g1565 ( 
.A(n_1429),
.B(n_1335),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1384),
.A2(n_1266),
.B1(n_1360),
.B2(n_1304),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1454),
.B(n_1420),
.Y(n_1567)
);

CKINVDCx6p67_ASAP7_75t_R g1568 ( 
.A(n_1489),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1493),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1433),
.A2(n_1266),
.B1(n_1306),
.B2(n_1335),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1472),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1472),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1393),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1491),
.B(n_1304),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1395),
.B(n_1297),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1386),
.A2(n_1340),
.B1(n_1304),
.B2(n_1320),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1515),
.A2(n_1283),
.B1(n_1287),
.B2(n_1367),
.C(n_1260),
.Y(n_1577)
);

CKINVDCx6p67_ASAP7_75t_R g1578 ( 
.A(n_1489),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1555),
.A2(n_1340),
.B1(n_1320),
.B2(n_1304),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1395),
.B(n_1320),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1491),
.B(n_1320),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1499),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1499),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1469),
.A2(n_1379),
.B1(n_1345),
.B2(n_1220),
.Y(n_1584)
);

BUFx8_ASAP7_75t_L g1585 ( 
.A(n_1397),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1503),
.A2(n_1340),
.B1(n_1279),
.B2(n_1261),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1507),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_SL g1588 ( 
.A1(n_1436),
.A2(n_1330),
.B(n_1315),
.C(n_1318),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1470),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1507),
.Y(n_1590)
);

OR2x6_ASAP7_75t_SL g1591 ( 
.A(n_1492),
.B(n_1303),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1399),
.A2(n_1337),
.B1(n_1318),
.B2(n_1315),
.C(n_1329),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1422),
.A2(n_1340),
.B1(n_1364),
.B2(n_1365),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1469),
.A2(n_1345),
.B1(n_1355),
.B2(n_1369),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1393),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1531),
.A2(n_1369),
.B(n_1355),
.C(n_1308),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1470),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1491),
.B(n_1364),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1403),
.B(n_1259),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1508),
.B(n_1343),
.Y(n_1600)
);

CKINVDCx6p67_ASAP7_75t_R g1601 ( 
.A(n_1440),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1484),
.A2(n_1368),
.B(n_1235),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1439),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1547),
.A2(n_1340),
.B1(n_1364),
.B2(n_1368),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1419),
.A2(n_1340),
.B1(n_1343),
.B2(n_32),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1512),
.B(n_1343),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1404),
.B(n_1235),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1449),
.A2(n_1235),
.B(n_1343),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1439),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1461),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1559),
.A2(n_1235),
.B(n_29),
.C(n_32),
.Y(n_1611)
);

BUFx4f_ASAP7_75t_SL g1612 ( 
.A(n_1431),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1512),
.B(n_158),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1447),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1516),
.B(n_28),
.Y(n_1615)
);

CKINVDCx6p67_ASAP7_75t_R g1616 ( 
.A(n_1408),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1563),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1516),
.B(n_34),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1419),
.A2(n_1455),
.B1(n_1563),
.B2(n_1519),
.Y(n_1619)
);

AOI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1406),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.C1(n_40),
.C2(n_41),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1397),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1419),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1512),
.B(n_155),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1519),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1424),
.B(n_145),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1380),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1508),
.B(n_45),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1463),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1455),
.B(n_56),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1414),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1510),
.B(n_1480),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1447),
.Y(n_1632)
);

AOI21xp33_ASAP7_75t_L g1633 ( 
.A1(n_1530),
.A2(n_62),
.B(n_68),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1398),
.A2(n_143),
.B(n_141),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1513),
.A2(n_70),
.B(n_74),
.Y(n_1635)
);

CKINVDCx6p67_ASAP7_75t_R g1636 ( 
.A(n_1408),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1510),
.B(n_74),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_SL g1638 ( 
.A(n_1556),
.B(n_140),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1476),
.Y(n_1639)
);

INVx5_ASAP7_75t_L g1640 ( 
.A(n_1533),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1414),
.B(n_1548),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1424),
.B(n_1490),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1473),
.A2(n_138),
.B(n_128),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1421),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1476),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1477),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1398),
.A2(n_76),
.B(n_79),
.Y(n_1647)
);

OR2x6_ASAP7_75t_L g1648 ( 
.A(n_1404),
.B(n_76),
.Y(n_1648)
);

INVx5_ASAP7_75t_L g1649 ( 
.A(n_1533),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1450),
.B(n_79),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1462),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1424),
.B(n_80),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1462),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1540),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1538),
.A2(n_98),
.B1(n_83),
.B2(n_84),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1428),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1548),
.B(n_80),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1417),
.B(n_83),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1504),
.B(n_84),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1540),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1432),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1428),
.Y(n_1662)
);

AOI222xp33_ASAP7_75t_L g1663 ( 
.A1(n_1554),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.C1(n_91),
.C2(n_92),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1518),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1461),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1504),
.A2(n_95),
.B1(n_89),
.B2(n_92),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1521),
.A2(n_88),
.B1(n_93),
.B2(n_1450),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1403),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1426),
.A2(n_93),
.B(n_1429),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1430),
.A2(n_1527),
.B1(n_1529),
.B2(n_1412),
.C(n_1385),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1428),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1521),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1482),
.B(n_1467),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1424),
.B(n_1490),
.Y(n_1674)
);

O2A1O1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1495),
.A2(n_1418),
.B(n_1446),
.C(n_1505),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1417),
.B(n_1450),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1450),
.B(n_1485),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1432),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1383),
.A2(n_1444),
.B1(n_1496),
.B2(n_1492),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1501),
.A2(n_1487),
.B1(n_1435),
.B2(n_1485),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1534),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1460),
.B(n_1518),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1404),
.B(n_1403),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1481),
.A2(n_1502),
.B(n_1537),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1552),
.A2(n_1404),
.B1(n_1474),
.B2(n_1429),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1460),
.B(n_1542),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1537),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1487),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1560),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_SL g1690 ( 
.A1(n_1552),
.A2(n_1429),
.B1(n_1408),
.B2(n_1413),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1500),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1506),
.B(n_1389),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1404),
.A2(n_1390),
.B(n_1427),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1498),
.A2(n_1557),
.B(n_1475),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1389),
.B(n_1500),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1474),
.A2(n_1390),
.B1(n_1465),
.B2(n_1539),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1383),
.B(n_1497),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1405),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1421),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1544),
.B(n_1456),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1461),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1394),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1456),
.B(n_1553),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1497),
.B(n_1490),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1390),
.A2(n_1533),
.B1(n_1438),
.B2(n_1556),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1390),
.A2(n_1427),
.B(n_1392),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1438),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1456),
.B(n_1562),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1545),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1490),
.B(n_1442),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1545),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1403),
.B(n_1390),
.Y(n_1712)
);

NAND2x1_ASAP7_75t_L g1713 ( 
.A(n_1533),
.B(n_1448),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1560),
.Y(n_1714)
);

BUFx10_ASAP7_75t_L g1715 ( 
.A(n_1541),
.Y(n_1715)
);

CKINVDCx11_ASAP7_75t_R g1716 ( 
.A(n_1461),
.Y(n_1716)
);

INVx3_ASAP7_75t_SL g1717 ( 
.A(n_1461),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1468),
.Y(n_1718)
);

CKINVDCx6p67_ASAP7_75t_R g1719 ( 
.A(n_1561),
.Y(n_1719)
);

AND2x2_ASAP7_75t_SL g1720 ( 
.A(n_1541),
.B(n_1392),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1468),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1535),
.A2(n_1411),
.B1(n_1474),
.B2(n_1514),
.C(n_1466),
.Y(n_1722)
);

CKINVDCx6p67_ASAP7_75t_R g1723 ( 
.A(n_1561),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1388),
.B(n_1452),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1394),
.Y(n_1725)
);

OR2x6_ASAP7_75t_L g1726 ( 
.A(n_1388),
.B(n_1452),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1541),
.A2(n_1400),
.B1(n_1474),
.B2(n_1442),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_R g1728 ( 
.A(n_1458),
.B(n_1451),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1405),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1402),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1453),
.B(n_1541),
.Y(n_1731)
);

CKINVDCx6p67_ASAP7_75t_R g1732 ( 
.A(n_1561),
.Y(n_1732)
);

INVx5_ASAP7_75t_L g1733 ( 
.A(n_1468),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1402),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1459),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1465),
.Y(n_1736)
);

OR2x6_ASAP7_75t_L g1737 ( 
.A(n_1388),
.B(n_1452),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1545),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1468),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_SL g1740 ( 
.A1(n_1413),
.A2(n_1539),
.B1(n_1525),
.B2(n_1526),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1511),
.A2(n_1523),
.B(n_1517),
.C(n_1532),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1465),
.A2(n_1539),
.B1(n_1400),
.B2(n_1483),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1448),
.B(n_1525),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1459),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1468),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1453),
.B(n_1551),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1524),
.A2(n_1478),
.B(n_1479),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1394),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1551),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1466),
.B(n_1486),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1488),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1459),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1466),
.B(n_1486),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1466),
.B(n_1486),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1558),
.B2(n_1400),
.Y(n_1755)
);

AND2x6_ASAP7_75t_L g1756 ( 
.A(n_1511),
.B(n_1532),
.Y(n_1756)
);

AO21x2_ASAP7_75t_L g1757 ( 
.A1(n_1502),
.A2(n_1543),
.B(n_1546),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1509),
.A2(n_1526),
.B1(n_1528),
.B2(n_1558),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1682),
.B(n_1486),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1641),
.B(n_1486),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1630),
.A2(n_1509),
.B1(n_1517),
.B2(n_1523),
.C(n_1528),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1624),
.A2(n_1546),
.B1(n_1543),
.B2(n_1416),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1630),
.A2(n_1549),
.B1(n_1410),
.B2(n_1423),
.C(n_1415),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1651),
.B(n_1451),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1704),
.B(n_1498),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1635),
.A2(n_1392),
.B(n_1471),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1566),
.A2(n_1550),
.B1(n_1488),
.B2(n_1451),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1730),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1567),
.A2(n_1416),
.B1(n_1387),
.B2(n_1391),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1567),
.A2(n_1416),
.B1(n_1387),
.B2(n_1391),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1673),
.B(n_1387),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1620),
.A2(n_1416),
.B1(n_1387),
.B2(n_1391),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1679),
.A2(n_1458),
.B1(n_1451),
.B2(n_1550),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1589),
.Y(n_1774)
);

AOI222xp33_ASAP7_75t_L g1775 ( 
.A1(n_1655),
.A2(n_1423),
.B1(n_1415),
.B2(n_1410),
.C1(n_1407),
.C2(n_1437),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1663),
.A2(n_1391),
.B1(n_1394),
.B2(n_1401),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1680),
.A2(n_1464),
.B1(n_1458),
.B2(n_1407),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1573),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1585),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1670),
.A2(n_1458),
.B1(n_1464),
.B2(n_1494),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1617),
.A2(n_1401),
.B1(n_1464),
.B2(n_1434),
.Y(n_1781)
);

CKINVDCx6p67_ASAP7_75t_R g1782 ( 
.A(n_1601),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1617),
.A2(n_1401),
.B1(n_1464),
.B2(n_1434),
.Y(n_1783)
);

AO21x1_ASAP7_75t_L g1784 ( 
.A1(n_1650),
.A2(n_1549),
.B(n_1522),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1655),
.A2(n_1401),
.B1(n_1437),
.B2(n_1382),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1729),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1704),
.B(n_1522),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1667),
.A2(n_1494),
.B1(n_1445),
.B2(n_1443),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1683),
.B(n_1409),
.Y(n_1789)
);

AO21x2_ASAP7_75t_L g1790 ( 
.A1(n_1669),
.A2(n_1409),
.B(n_1443),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1633),
.A2(n_1520),
.B1(n_1396),
.B2(n_1381),
.C(n_1536),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1692),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1648),
.A2(n_1536),
.B1(n_1396),
.B2(n_1445),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1667),
.A2(n_1536),
.B1(n_1520),
.B2(n_1381),
.C(n_1425),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1724),
.B(n_1726),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1652),
.B(n_1425),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1619),
.A2(n_1536),
.B1(n_1441),
.B2(n_1457),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1622),
.A2(n_1441),
.B1(n_1457),
.B2(n_1666),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1612),
.Y(n_1799)
);

AND2x6_ASAP7_75t_SL g1800 ( 
.A(n_1657),
.B(n_1695),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1622),
.A2(n_1666),
.B1(n_1619),
.B2(n_1570),
.C(n_1611),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1648),
.A2(n_1604),
.B(n_1650),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1611),
.A2(n_1570),
.B1(n_1605),
.B2(n_1672),
.C(n_1629),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1648),
.A2(n_1605),
.B1(n_1604),
.B2(n_1575),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1669),
.A2(n_1626),
.B1(n_1653),
.B2(n_1637),
.C(n_1627),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1621),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1577),
.A2(n_1579),
.B1(n_1576),
.B2(n_1690),
.C(n_1643),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1612),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1697),
.B(n_1677),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1716),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1683),
.B(n_1712),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1618),
.B(n_1686),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1597),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1631),
.B(n_1580),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1659),
.A2(n_1691),
.B1(n_1625),
.B2(n_1576),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1579),
.A2(n_1658),
.B1(n_1664),
.B2(n_1626),
.Y(n_1817)
);

BUFx12f_ASAP7_75t_L g1818 ( 
.A(n_1661),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1595),
.A2(n_1585),
.B1(n_1625),
.B2(n_1722),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1654),
.B(n_1660),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1688),
.A2(n_1690),
.B1(n_1707),
.B2(n_1711),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1602),
.A2(n_1685),
.B(n_1643),
.C(n_1720),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1595),
.A2(n_1578),
.B1(n_1568),
.B2(n_1676),
.Y(n_1824)
);

OAI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1675),
.A2(n_1596),
.B(n_1685),
.C(n_1742),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1600),
.B(n_1571),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1642),
.B(n_1674),
.Y(n_1827)
);

OA21x2_ASAP7_75t_L g1828 ( 
.A1(n_1602),
.A2(n_1608),
.B(n_1696),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1564),
.A2(n_1569),
.B1(n_1703),
.B2(n_1572),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1582),
.A2(n_1590),
.B1(n_1587),
.B2(n_1583),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1603),
.B(n_1609),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1616),
.A2(n_1636),
.B1(n_1674),
.B2(n_1628),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1708),
.B(n_1738),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1675),
.A2(n_1586),
.B1(n_1592),
.B2(n_1588),
.C(n_1696),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1614),
.A2(n_1632),
.B1(n_1586),
.B2(n_1606),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1588),
.A2(n_1742),
.B1(n_1694),
.B2(n_1594),
.C(n_1656),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1639),
.B(n_1645),
.Y(n_1838)
);

AOI222xp33_ASAP7_75t_L g1839 ( 
.A1(n_1720),
.A2(n_1638),
.B1(n_1699),
.B2(n_1646),
.C1(n_1613),
.C2(n_1623),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1574),
.B(n_1581),
.Y(n_1840)
);

AOI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1594),
.A2(n_1565),
.B(n_1727),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1746),
.B(n_1709),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1591),
.A2(n_1565),
.B1(n_1640),
.B2(n_1649),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1574),
.B(n_1581),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1606),
.A2(n_1613),
.B1(n_1623),
.B2(n_1683),
.Y(n_1845)
);

AO21x2_ASAP7_75t_L g1846 ( 
.A1(n_1758),
.A2(n_1706),
.B(n_1693),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1721),
.B(n_1644),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1734),
.B(n_1749),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1705),
.A2(n_1736),
.B1(n_1706),
.B2(n_1693),
.C(n_1584),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1681),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1678),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1687),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1689),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1740),
.A2(n_1593),
.B1(n_1723),
.B2(n_1732),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1712),
.A2(n_1715),
.B1(n_1724),
.B2(n_1726),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1714),
.B(n_1712),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1740),
.A2(n_1593),
.B1(n_1719),
.B2(n_1755),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1656),
.A2(n_1671),
.B1(n_1662),
.B2(n_1754),
.C(n_1753),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1721),
.B(n_1749),
.Y(n_1859)
);

BUFx4f_ASAP7_75t_SL g1860 ( 
.A(n_1717),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1715),
.A2(n_1647),
.B1(n_1755),
.B2(n_1607),
.Y(n_1861)
);

INVx11_ASAP7_75t_L g1862 ( 
.A(n_1756),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1698),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1749),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1733),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1724),
.A2(n_1726),
.B1(n_1737),
.B2(n_1743),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1734),
.B(n_1717),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_SL g1868 ( 
.A1(n_1662),
.A2(n_1671),
.B(n_1752),
.C(n_1744),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1640),
.A2(n_1649),
.B1(n_1607),
.B2(n_1737),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1735),
.A2(n_1752),
.B(n_1744),
.C(n_1750),
.Y(n_1870)
);

OAI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1735),
.A2(n_1634),
.B(n_1741),
.C(n_1698),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1607),
.A2(n_1737),
.B1(n_1634),
.B2(n_1741),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1610),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1745),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1718),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1610),
.B(n_1739),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1756),
.Y(n_1877)
);

BUFx12f_ASAP7_75t_L g1878 ( 
.A(n_1610),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_L g1879 ( 
.A(n_1743),
.B(n_1728),
.C(n_1745),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1610),
.B(n_1739),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1684),
.A2(n_1725),
.B1(n_1748),
.B2(n_1702),
.C(n_1751),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1665),
.B(n_1739),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1598),
.B(n_1733),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1743),
.A2(n_1640),
.B1(n_1649),
.B2(n_1668),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1640),
.A2(n_1649),
.B1(n_1668),
.B2(n_1598),
.Y(n_1885)
);

OAI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1733),
.A2(n_1728),
.B1(n_1665),
.B2(n_1739),
.Y(n_1886)
);

AOI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1684),
.A2(n_1713),
.B(n_1599),
.Y(n_1887)
);

CKINVDCx8_ASAP7_75t_R g1888 ( 
.A(n_1665),
.Y(n_1888)
);

AOI21xp33_ASAP7_75t_L g1889 ( 
.A1(n_1599),
.A2(n_1757),
.B(n_1701),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1756),
.A2(n_1733),
.B1(n_1701),
.B2(n_1747),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1701),
.Y(n_1891)
);

OAI221xp5_ASAP7_75t_L g1892 ( 
.A1(n_1617),
.A2(n_1454),
.B1(n_881),
.B2(n_876),
.C(n_748),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1589),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1635),
.A2(n_1436),
.B(n_1611),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1630),
.A2(n_748),
.B1(n_1567),
.B2(n_1300),
.C(n_477),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1630),
.A2(n_748),
.B1(n_1567),
.B2(n_1300),
.C(n_477),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1621),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1635),
.A2(n_1611),
.B(n_1567),
.C(n_1559),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1635),
.A2(n_1436),
.B(n_1611),
.Y(n_1902)
);

NOR2xp67_ASAP7_75t_L g1903 ( 
.A(n_1595),
.B(n_1099),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1573),
.B(n_935),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_L g1905 ( 
.A(n_1573),
.B(n_911),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1566),
.A2(n_1384),
.B1(n_1136),
.B2(n_1469),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1635),
.A2(n_1224),
.B(n_1559),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1692),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1566),
.A2(n_1384),
.B1(n_1136),
.B2(n_1469),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1692),
.Y(n_1913)
);

AOI222xp33_ASAP7_75t_L g1914 ( 
.A1(n_1566),
.A2(n_1300),
.B1(n_916),
.B2(n_1433),
.C1(n_1567),
.C2(n_410),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1567),
.B(n_1673),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1635),
.A2(n_1224),
.B(n_1559),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_R g1919 ( 
.A(n_1573),
.B(n_1229),
.Y(n_1919)
);

BUFx4f_ASAP7_75t_SL g1920 ( 
.A(n_1601),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1635),
.A2(n_1611),
.B(n_1567),
.C(n_1559),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1624),
.A2(n_1630),
.B1(n_1433),
.B2(n_1635),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1567),
.A2(n_1454),
.B(n_1419),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1567),
.A2(n_1620),
.B1(n_1663),
.B2(n_1433),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1892),
.A2(n_1927),
.B1(n_1926),
.B2(n_1898),
.C(n_1912),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1862),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1828),
.B(n_1759),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1916),
.B(n_1771),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1786),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1786),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1863),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1795),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1812),
.B(n_1789),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1868),
.B(n_1879),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1812),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1828),
.B(n_1760),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1768),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1809),
.B(n_1764),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1828),
.B(n_1823),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1774),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1850),
.B(n_1852),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1789),
.B(n_1877),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1789),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1898),
.A2(n_1927),
.B1(n_1926),
.B2(n_1910),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1899),
.A2(n_1901),
.B1(n_1912),
.B2(n_1921),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1853),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1814),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_SL g1951 ( 
.A(n_1810),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1866),
.B(n_1856),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1823),
.B(n_1769),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1826),
.B(n_1815),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1810),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1769),
.B(n_1770),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1770),
.B(n_1846),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1893),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1899),
.A2(n_1901),
.B1(n_1915),
.B2(n_1917),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1846),
.B(n_1841),
.Y(n_1960)
);

NOR2x1p5_ASAP7_75t_L g1961 ( 
.A(n_1810),
.B(n_1782),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1777),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1831),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1838),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1806),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1855),
.B(n_1796),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1837),
.B(n_1781),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1830),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1830),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1790),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1781),
.B(n_1783),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1810),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1867),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1848),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1815),
.B(n_1835),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1802),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1870),
.B(n_1820),
.Y(n_1977)
);

AO31x2_ASAP7_75t_L g1978 ( 
.A1(n_1900),
.A2(n_1923),
.A3(n_1766),
.B(n_1918),
.Y(n_1978)
);

NAND2x1p5_ASAP7_75t_L g1979 ( 
.A(n_1907),
.B(n_1788),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1783),
.B(n_1787),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1784),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1765),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1897),
.B(n_1857),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1922),
.B(n_1835),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1869),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1797),
.A2(n_1785),
.B(n_1861),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1805),
.B(n_1858),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1780),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1849),
.B(n_1872),
.Y(n_1989)
);

OR2x6_ASAP7_75t_L g1990 ( 
.A(n_1894),
.B(n_1902),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1880),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1860),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1881),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1872),
.B(n_1836),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1908),
.A2(n_1917),
.B1(n_1915),
.B2(n_1910),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1869),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1860),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1925),
.B(n_1792),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1794),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1871),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1773),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1843),
.B(n_1825),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1882),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1909),
.B(n_1913),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1785),
.B(n_1836),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1829),
.B(n_1900),
.Y(n_2006)
);

NOR2x1_ASAP7_75t_L g2007 ( 
.A(n_1843),
.B(n_1886),
.Y(n_2007)
);

NAND2x1p5_ASAP7_75t_L g2008 ( 
.A(n_1865),
.B(n_1874),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1772),
.B(n_1861),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1886),
.Y(n_2010)
);

NAND2x1_ASAP7_75t_L g2011 ( 
.A(n_1884),
.B(n_1885),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1878),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_1793),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1923),
.B(n_1834),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1799),
.B(n_1808),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1772),
.B(n_1767),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1890),
.B(n_1775),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1876),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1793),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1889),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1887),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1776),
.B(n_1804),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1821),
.B(n_1842),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1762),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1761),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1884),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1833),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1992),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1945),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_SL g2030 ( 
.A1(n_1990),
.A2(n_1921),
.B1(n_1908),
.B2(n_1920),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1980),
.B(n_1819),
.Y(n_2031)
);

NAND3xp33_ASAP7_75t_L g2032 ( 
.A(n_1990),
.B(n_1896),
.C(n_1895),
.Y(n_2032)
);

AND2x6_ASAP7_75t_L g2033 ( 
.A(n_1936),
.B(n_2007),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1980),
.B(n_1819),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1970),
.A2(n_1854),
.B(n_1791),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1932),
.Y(n_2036)
);

AOI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_1928),
.A2(n_1924),
.B1(n_1801),
.B2(n_1906),
.C(n_1911),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1990),
.A2(n_1924),
.B(n_1914),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1949),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1991),
.Y(n_2040)
);

BUFx2_ASAP7_75t_L g2041 ( 
.A(n_2027),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1980),
.B(n_1859),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1945),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_L g2044 ( 
.A(n_1990),
.B(n_1803),
.C(n_1804),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1947),
.A2(n_1816),
.B1(n_1798),
.B2(n_1824),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1949),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1941),
.B(n_1817),
.Y(n_2047)
);

OAI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1990),
.A2(n_1807),
.B1(n_1822),
.B2(n_1920),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1949),
.Y(n_2049)
);

OAI211xp5_ASAP7_75t_L g2050 ( 
.A1(n_1948),
.A2(n_1798),
.B(n_1817),
.C(n_1839),
.Y(n_2050)
);

INVx2_ASAP7_75t_SL g2051 ( 
.A(n_1991),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1977),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1992),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1950),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1939),
.B(n_1844),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1990),
.A2(n_1845),
.B(n_1885),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_2014),
.B(n_1800),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1939),
.B(n_1811),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1928),
.A2(n_2014),
.B1(n_1976),
.B2(n_2022),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_1936),
.B(n_1864),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1939),
.B(n_1813),
.Y(n_2061)
);

AND2x4_ASAP7_75t_SL g2062 ( 
.A(n_1929),
.B(n_1865),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1987),
.A2(n_1845),
.B(n_1776),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_SL g2064 ( 
.A(n_1998),
.B(n_1987),
.C(n_2000),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2027),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1951),
.Y(n_2066)
);

NOR2x1_ASAP7_75t_L g2067 ( 
.A(n_1937),
.B(n_1903),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1959),
.A2(n_1832),
.B1(n_1824),
.B2(n_1875),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1950),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1950),
.Y(n_2070)
);

AO21x1_ASAP7_75t_SL g2071 ( 
.A1(n_2002),
.A2(n_1832),
.B(n_1763),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2025),
.A2(n_1847),
.B1(n_1779),
.B2(n_1905),
.C(n_1840),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1934),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1979),
.A2(n_1883),
.B(n_1904),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1998),
.B(n_1847),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1982),
.B(n_1827),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_1974),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1974),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1982),
.B(n_1873),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1941),
.B(n_1891),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1977),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_2004),
.Y(n_2082)
);

NOR4xp25_ASAP7_75t_SL g2083 ( 
.A(n_1976),
.B(n_1778),
.C(n_1851),
.D(n_1888),
.Y(n_2083)
);

AOI211xp5_ASAP7_75t_L g2084 ( 
.A1(n_1960),
.A2(n_1919),
.B(n_1874),
.C(n_1818),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1934),
.Y(n_2085)
);

OAI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_1995),
.A2(n_1919),
.B1(n_1979),
.B2(n_2006),
.C(n_2025),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1943),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_2019),
.B(n_2001),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1975),
.A2(n_2002),
.B1(n_2006),
.B2(n_1954),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1943),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1975),
.A2(n_1954),
.B1(n_2017),
.B2(n_1967),
.Y(n_2091)
);

AOI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_1989),
.A2(n_1993),
.B(n_2000),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1933),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1944),
.Y(n_2094)
);

OAI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_1979),
.A2(n_2001),
.B1(n_1993),
.B2(n_2011),
.C(n_2004),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2022),
.A2(n_1967),
.B1(n_1994),
.B2(n_2016),
.Y(n_2096)
);

OAI33xp33_ASAP7_75t_L g2097 ( 
.A1(n_1965),
.A2(n_1931),
.A3(n_1969),
.B1(n_1968),
.B2(n_1983),
.B3(n_2020),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1931),
.B(n_1973),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1933),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2003),
.B(n_1930),
.Y(n_2100)
);

OAI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_1979),
.A2(n_2011),
.B1(n_1937),
.B2(n_1962),
.C(n_2013),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1936),
.B(n_1945),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1940),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1958),
.Y(n_2104)
);

NAND4xp25_ASAP7_75t_L g2105 ( 
.A(n_1967),
.B(n_1965),
.C(n_1989),
.D(n_1983),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1940),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2039),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2036),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2052),
.B(n_1973),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2046),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_2041),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2100),
.B(n_2061),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2081),
.B(n_2020),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_2029),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2036),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2061),
.B(n_1930),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2088),
.B(n_2019),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2049),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2058),
.B(n_1953),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2082),
.B(n_1960),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2054),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2058),
.B(n_1953),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_2029),
.Y(n_2123)
);

OR2x2_ASAP7_75t_L g2124 ( 
.A(n_2077),
.B(n_2013),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2078),
.B(n_1960),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2055),
.B(n_1953),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2098),
.B(n_2073),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2055),
.B(n_1942),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2069),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2085),
.B(n_1962),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2042),
.B(n_1942),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2042),
.B(n_1942),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2087),
.B(n_1988),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_2084),
.B(n_1935),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2029),
.B(n_2043),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_2065),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2090),
.B(n_2024),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2070),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_SL g2139 ( 
.A(n_2032),
.B(n_2007),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2043),
.B(n_1936),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2040),
.B(n_1988),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2043),
.B(n_1945),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_2080),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2040),
.B(n_1988),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2102),
.B(n_1966),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2102),
.B(n_1966),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2102),
.B(n_1966),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2051),
.B(n_1978),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2060),
.B(n_1946),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2096),
.B(n_2024),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2051),
.B(n_1952),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2060),
.B(n_1946),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2104),
.B(n_1963),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2094),
.B(n_1978),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2080),
.B(n_1978),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2075),
.B(n_1963),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2093),
.B(n_1978),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2099),
.B(n_1978),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2076),
.B(n_1952),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_2089),
.B(n_1984),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2075),
.B(n_1964),
.Y(n_2161)
);

INVxp67_ASAP7_75t_SL g2162 ( 
.A(n_2099),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2076),
.B(n_2031),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2031),
.B(n_1957),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2103),
.B(n_1978),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2131),
.B(n_2060),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2139),
.B(n_2057),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2125),
.B(n_1978),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2108),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2107),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_SL g2171 ( 
.A(n_2139),
.B(n_2101),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2125),
.B(n_2047),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2107),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2110),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2109),
.B(n_2091),
.Y(n_2175)
);

NAND2x1p5_ASAP7_75t_L g2176 ( 
.A(n_2134),
.B(n_1935),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2131),
.B(n_2033),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2110),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2109),
.B(n_2095),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_2145),
.B(n_2146),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2132),
.B(n_2033),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2132),
.B(n_2033),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2128),
.B(n_2033),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2128),
.B(n_2033),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2155),
.B(n_2047),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2108),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2111),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2111),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2155),
.B(n_2035),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_L g2190 ( 
.A(n_2150),
.B(n_2038),
.C(n_2067),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2118),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_2145),
.B(n_1935),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2160),
.B(n_2092),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2160),
.B(n_2057),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2150),
.B(n_2086),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2156),
.B(n_2034),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2156),
.B(n_2034),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2164),
.B(n_2126),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2108),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2115),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2161),
.B(n_2063),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2118),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2161),
.B(n_2105),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_2136),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2121),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2146),
.B(n_1946),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2126),
.B(n_1984),
.Y(n_2207)
);

NOR2x1p5_ASAP7_75t_SL g2208 ( 
.A(n_2157),
.B(n_1970),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2115),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2115),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2120),
.B(n_2035),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2119),
.B(n_2018),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2121),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2147),
.B(n_1946),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2129),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2164),
.B(n_2033),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2129),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2138),
.Y(n_2218)
);

NAND2x1p5_ASAP7_75t_L g2219 ( 
.A(n_2136),
.B(n_1938),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2120),
.B(n_2106),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2119),
.B(n_2079),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2127),
.B(n_1955),
.Y(n_2222)
);

OAI31xp33_ASAP7_75t_L g2223 ( 
.A1(n_2171),
.A2(n_2048),
.A3(n_2050),
.B(n_2044),
.Y(n_2223)
);

NOR2x1_ASAP7_75t_L g2224 ( 
.A(n_2167),
.B(n_1961),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2216),
.B(n_2122),
.Y(n_2225)
);

AO21x1_ASAP7_75t_L g2226 ( 
.A1(n_2190),
.A2(n_2113),
.B(n_2045),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2169),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2216),
.B(n_2122),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2195),
.A2(n_2064),
.B1(n_2059),
.B2(n_2037),
.Y(n_2229)
);

NOR4xp25_ASAP7_75t_SL g2230 ( 
.A(n_2176),
.B(n_2066),
.C(n_2097),
.D(n_2072),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2170),
.Y(n_2231)
);

NAND5xp2_ASAP7_75t_SL g2232 ( 
.A(n_2177),
.B(n_2066),
.C(n_2074),
.D(n_2068),
.E(n_2017),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2170),
.Y(n_2233)
);

NAND2xp33_ASAP7_75t_R g2234 ( 
.A(n_2194),
.B(n_2083),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2173),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2201),
.B(n_2113),
.Y(n_2236)
);

OAI211xp5_ASAP7_75t_L g2237 ( 
.A1(n_2193),
.A2(n_2179),
.B(n_2203),
.C(n_2175),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2173),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2169),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2177),
.B(n_2147),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2174),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2186),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2172),
.B(n_2124),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2186),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2196),
.B(n_2163),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2176),
.A2(n_2016),
.B(n_1986),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2181),
.B(n_2142),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2199),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2174),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2197),
.B(n_2163),
.Y(n_2250)
);

OAI22x1_ASAP7_75t_L g2251 ( 
.A1(n_2176),
.A2(n_1961),
.B1(n_2143),
.B2(n_2114),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2172),
.B(n_2124),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2187),
.B(n_2143),
.Y(n_2253)
);

NAND2xp33_ASAP7_75t_R g2254 ( 
.A(n_2181),
.B(n_2015),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2199),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2178),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2182),
.B(n_2142),
.Y(n_2257)
);

NAND2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2182),
.B(n_1951),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2188),
.A2(n_2030),
.B(n_2056),
.Y(n_2259)
);

OR2x6_ASAP7_75t_L g2260 ( 
.A(n_2219),
.B(n_2028),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2204),
.B(n_2192),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2178),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2183),
.B(n_2135),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2191),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2180),
.B(n_2149),
.Y(n_2265)
);

OAI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_2168),
.A2(n_2016),
.B(n_2017),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2183),
.B(n_2135),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2184),
.B(n_2135),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2207),
.B(n_2127),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_2198),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2184),
.B(n_2149),
.Y(n_2271)
);

NOR3xp33_ASAP7_75t_SL g2272 ( 
.A(n_2222),
.B(n_2137),
.C(n_2026),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2221),
.B(n_2159),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2200),
.Y(n_2274)
);

NAND3xp33_ASAP7_75t_L g2275 ( 
.A(n_2211),
.B(n_2022),
.C(n_2021),
.Y(n_2275)
);

INVx4_ASAP7_75t_L g2276 ( 
.A(n_2219),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2191),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2185),
.B(n_2130),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2226),
.A2(n_2009),
.B1(n_1971),
.B2(n_2192),
.Y(n_2279)
);

AOI322xp5_ASAP7_75t_L g2280 ( 
.A1(n_2266),
.A2(n_2198),
.A3(n_2009),
.B1(n_1971),
.B2(n_1994),
.C1(n_2221),
.C2(n_2005),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2231),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2226),
.A2(n_2211),
.B(n_2137),
.Y(n_2282)
);

AOI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2229),
.A2(n_2237),
.B1(n_2232),
.B2(n_2223),
.C(n_2275),
.Y(n_2283)
);

OAI32xp33_ASAP7_75t_L g2284 ( 
.A1(n_2234),
.A2(n_2168),
.A3(n_2189),
.B1(n_2219),
.B2(n_2185),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2224),
.B(n_2192),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2224),
.B(n_2236),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2259),
.A2(n_2009),
.B1(n_2189),
.B2(n_1971),
.Y(n_2287)
);

AOI31xp33_ASAP7_75t_L g2288 ( 
.A1(n_2254),
.A2(n_1951),
.A3(n_2180),
.B(n_2008),
.Y(n_2288)
);

AND2x4_ASAP7_75t_SL g2289 ( 
.A(n_2260),
.B(n_1929),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2231),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2243),
.B(n_2212),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2233),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2233),
.Y(n_2293)
);

OAI221xp5_ASAP7_75t_L g2294 ( 
.A1(n_2246),
.A2(n_1972),
.B1(n_1955),
.B2(n_1999),
.C(n_2028),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2261),
.A2(n_2206),
.B1(n_2214),
.B2(n_2180),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2235),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_L g2297 ( 
.A(n_2230),
.B(n_2021),
.C(n_2026),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2269),
.B(n_2202),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2243),
.B(n_2220),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2252),
.B(n_2220),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2265),
.Y(n_2301)
);

OAI21xp33_ASAP7_75t_SL g2302 ( 
.A1(n_2276),
.A2(n_2166),
.B(n_2112),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2252),
.B(n_2154),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2235),
.Y(n_2304)
);

OAI21xp33_ASAP7_75t_SL g2305 ( 
.A1(n_2276),
.A2(n_2166),
.B(n_2112),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2238),
.Y(n_2306)
);

OAI21xp33_ASAP7_75t_L g2307 ( 
.A1(n_2272),
.A2(n_2154),
.B(n_1957),
.Y(n_2307)
);

OAI21xp33_ASAP7_75t_L g2308 ( 
.A1(n_2251),
.A2(n_2148),
.B(n_2208),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2238),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2232),
.A2(n_1986),
.B(n_2005),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2253),
.Y(n_2311)
);

OAI21xp33_ASAP7_75t_SL g2312 ( 
.A1(n_2276),
.A2(n_2114),
.B(n_2218),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2241),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2258),
.A2(n_2214),
.B1(n_2206),
.B2(n_2005),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2265),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2240),
.B(n_2206),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2251),
.A2(n_1938),
.B1(n_1999),
.B2(n_1986),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2245),
.B(n_2202),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2250),
.B(n_2205),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2241),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_2311),
.Y(n_2321)
);

OAI221xp5_ASAP7_75t_L g2322 ( 
.A1(n_2283),
.A2(n_2260),
.B1(n_2270),
.B2(n_2278),
.C(n_2256),
.Y(n_2322)
);

INVxp67_ASAP7_75t_SL g2323 ( 
.A(n_2286),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2301),
.B(n_2315),
.Y(n_2324)
);

OR2x6_ASAP7_75t_L g2325 ( 
.A(n_2285),
.B(n_2260),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2279),
.B(n_2280),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2287),
.B(n_2288),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2281),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2287),
.A2(n_2260),
.B(n_2277),
.Y(n_2329)
);

OAI221xp5_ASAP7_75t_SL g2330 ( 
.A1(n_2297),
.A2(n_2278),
.B1(n_2148),
.B2(n_2228),
.C(n_2225),
.Y(n_2330)
);

OAI211xp5_ASAP7_75t_SL g2331 ( 
.A1(n_2317),
.A2(n_2294),
.B(n_2282),
.C(n_2310),
.Y(n_2331)
);

AOI211xp5_ASAP7_75t_L g2332 ( 
.A1(n_2284),
.A2(n_1992),
.B(n_1997),
.C(n_1972),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2290),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2292),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2293),
.Y(n_2335)
);

OAI321xp33_ASAP7_75t_L g2336 ( 
.A1(n_2310),
.A2(n_2277),
.A3(n_2264),
.B1(n_2262),
.B2(n_2256),
.C(n_2249),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2294),
.A2(n_2249),
.B(n_2264),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2295),
.B(n_2240),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2307),
.A2(n_2262),
.B(n_2265),
.Y(n_2339)
);

NAND2x1p5_ASAP7_75t_L g2340 ( 
.A(n_2314),
.B(n_1997),
.Y(n_2340)
);

OAI32xp33_ASAP7_75t_L g2341 ( 
.A1(n_2302),
.A2(n_2225),
.A3(n_2228),
.B1(n_2268),
.B2(n_2267),
.Y(n_2341)
);

NOR2x1_ASAP7_75t_L g2342 ( 
.A(n_2296),
.B(n_1997),
.Y(n_2342)
);

AND2x2_ASAP7_75t_SL g2343 ( 
.A(n_2289),
.B(n_1929),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2298),
.B(n_2273),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2305),
.B(n_2271),
.Y(n_2345)
);

OAI21xp33_ASAP7_75t_L g2346 ( 
.A1(n_2318),
.A2(n_2263),
.B(n_2267),
.Y(n_2346)
);

OAI22xp33_ASAP7_75t_SL g2347 ( 
.A1(n_2299),
.A2(n_2114),
.B1(n_2123),
.B2(n_2274),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2316),
.B(n_2271),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2304),
.Y(n_2349)
);

AOI322xp5_ASAP7_75t_L g2350 ( 
.A1(n_2308),
.A2(n_2268),
.A3(n_2263),
.B1(n_2257),
.B2(n_2247),
.C1(n_2116),
.C2(n_1956),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2318),
.A2(n_2247),
.B1(n_2257),
.B2(n_1951),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2328),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2333),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2322),
.A2(n_2312),
.B(n_2298),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2323),
.B(n_2319),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2321),
.B(n_2324),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2334),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2348),
.B(n_2325),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2335),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2342),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2325),
.B(n_2319),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2344),
.B(n_2300),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2325),
.Y(n_2363)
);

NAND2x1p5_ASAP7_75t_SL g2364 ( 
.A(n_2345),
.B(n_2227),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2349),
.Y(n_2365)
);

XNOR2xp5_ASAP7_75t_L g2366 ( 
.A(n_2351),
.B(n_1955),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2324),
.B(n_2320),
.Y(n_2367)
);

AOI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2331),
.A2(n_2313),
.B1(n_2309),
.B2(n_2306),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2346),
.Y(n_2369)
);

XNOR2x1_ASAP7_75t_L g2370 ( 
.A(n_2326),
.B(n_1972),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2338),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2332),
.A2(n_2291),
.B1(n_2303),
.B2(n_2053),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2339),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2336),
.B(n_2053),
.Y(n_2374)
);

OR2x2_ASAP7_75t_L g2375 ( 
.A(n_2330),
.B(n_2227),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_R g2376 ( 
.A(n_2343),
.B(n_2012),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2356),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2358),
.Y(n_2378)
);

NOR3xp33_ASAP7_75t_L g2379 ( 
.A(n_2363),
.B(n_2327),
.C(n_2332),
.Y(n_2379)
);

NOR3xp33_ASAP7_75t_SL g2380 ( 
.A(n_2371),
.B(n_2341),
.C(n_2329),
.Y(n_2380)
);

NAND3xp33_ASAP7_75t_L g2381 ( 
.A(n_2368),
.B(n_2350),
.C(n_2337),
.Y(n_2381)
);

NOR2x1_ASAP7_75t_L g2382 ( 
.A(n_2360),
.B(n_2239),
.Y(n_2382)
);

OAI211xp5_ASAP7_75t_SL g2383 ( 
.A1(n_2373),
.A2(n_2340),
.B(n_2347),
.C(n_2255),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2376),
.B(n_2363),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2367),
.Y(n_2385)
);

AOI211xp5_ASAP7_75t_L g2386 ( 
.A1(n_2354),
.A2(n_2340),
.B(n_2012),
.C(n_2274),
.Y(n_2386)
);

O2A1O1Ixp33_ASAP7_75t_L g2387 ( 
.A1(n_2374),
.A2(n_2255),
.B(n_2248),
.C(n_2244),
.Y(n_2387)
);

INVx1_ASAP7_75t_SL g2388 ( 
.A(n_2358),
.Y(n_2388)
);

AOI221x1_ASAP7_75t_L g2389 ( 
.A1(n_2364),
.A2(n_2248),
.B1(n_2244),
.B2(n_2242),
.C(n_2239),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2370),
.B(n_2242),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2370),
.B(n_2369),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2381),
.A2(n_2374),
.B1(n_2375),
.B2(n_2372),
.Y(n_2392)
);

OAI211xp5_ASAP7_75t_SL g2393 ( 
.A1(n_2380),
.A2(n_2355),
.B(n_2353),
.C(n_2365),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2391),
.A2(n_2361),
.B(n_2366),
.Y(n_2394)
);

NOR2x1_ASAP7_75t_L g2395 ( 
.A(n_2378),
.B(n_2352),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2379),
.A2(n_2361),
.B1(n_2362),
.B2(n_2357),
.Y(n_2396)
);

AOI221x1_ASAP7_75t_L g2397 ( 
.A1(n_2377),
.A2(n_2364),
.B1(n_2359),
.B2(n_2376),
.C(n_2218),
.Y(n_2397)
);

AOI221x1_ASAP7_75t_L g2398 ( 
.A1(n_2385),
.A2(n_2217),
.B1(n_2215),
.B2(n_2205),
.C(n_2213),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2388),
.B(n_2215),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2382),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2384),
.B(n_2012),
.Y(n_2401)
);

AOI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2383),
.A2(n_2386),
.B1(n_2390),
.B2(n_2387),
.C(n_2389),
.Y(n_2402)
);

OAI221xp5_ASAP7_75t_L g2403 ( 
.A1(n_2383),
.A2(n_2130),
.B1(n_2123),
.B2(n_2217),
.C(n_1999),
.Y(n_2403)
);

BUFx12f_ASAP7_75t_L g2404 ( 
.A(n_2401),
.Y(n_2404)
);

OAI332xp33_ASAP7_75t_L g2405 ( 
.A1(n_2400),
.A2(n_2117),
.A3(n_2010),
.B1(n_2158),
.B2(n_2157),
.B3(n_2165),
.C1(n_1996),
.C2(n_1985),
.Y(n_2405)
);

INVx3_ASAP7_75t_L g2406 ( 
.A(n_2399),
.Y(n_2406)
);

AOI22xp33_ASAP7_75t_R g2407 ( 
.A1(n_2393),
.A2(n_1981),
.B1(n_2071),
.B2(n_1968),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2396),
.B(n_2214),
.Y(n_2408)
);

AOI21xp33_ASAP7_75t_SL g2409 ( 
.A1(n_2392),
.A2(n_2117),
.B(n_2008),
.Y(n_2409)
);

OAI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2395),
.A2(n_2210),
.B(n_2209),
.Y(n_2410)
);

BUFx12f_ASAP7_75t_L g2411 ( 
.A(n_2404),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2409),
.B(n_2402),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2406),
.Y(n_2413)
);

AO22x2_ASAP7_75t_L g2414 ( 
.A1(n_2406),
.A2(n_2397),
.B1(n_2394),
.B2(n_2398),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2408),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_SL g2416 ( 
.A(n_2410),
.B(n_2403),
.C(n_2153),
.Y(n_2416)
);

NOR4xp25_ASAP7_75t_L g2417 ( 
.A(n_2407),
.B(n_2210),
.C(n_2209),
.D(n_2200),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2405),
.B(n_2123),
.Y(n_2418)
);

OAI211xp5_ASAP7_75t_SL g2419 ( 
.A1(n_2412),
.A2(n_2405),
.B(n_2153),
.C(n_2123),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2413),
.B(n_2133),
.C(n_2158),
.Y(n_2420)
);

NAND3xp33_ASAP7_75t_SL g2421 ( 
.A(n_2413),
.B(n_2008),
.C(n_1929),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2414),
.B(n_2138),
.Y(n_2422)
);

AOI21xp33_ASAP7_75t_SL g2423 ( 
.A1(n_2414),
.A2(n_2008),
.B(n_2133),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2415),
.Y(n_2424)
);

CKINVDCx12_ASAP7_75t_R g2425 ( 
.A(n_2424),
.Y(n_2425)
);

O2A1O1Ixp5_ASAP7_75t_L g2426 ( 
.A1(n_2422),
.A2(n_2418),
.B(n_2411),
.C(n_2417),
.Y(n_2426)
);

NOR3xp33_ASAP7_75t_L g2427 ( 
.A(n_2423),
.B(n_2418),
.C(n_2416),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2421),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_2428),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2429),
.Y(n_2430)
);

AOI22xp5_ASAP7_75t_SL g2431 ( 
.A1(n_2430),
.A2(n_2425),
.B1(n_2426),
.B2(n_2427),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2430),
.B(n_2420),
.Y(n_2432)
);

NAND3xp33_ASAP7_75t_L g2433 ( 
.A(n_2431),
.B(n_2432),
.C(n_2419),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2431),
.Y(n_2434)
);

XNOR2xp5_ASAP7_75t_L g2435 ( 
.A(n_2433),
.B(n_2062),
.Y(n_2435)
);

AOI31xp33_ASAP7_75t_L g2436 ( 
.A1(n_2434),
.A2(n_2023),
.A3(n_2144),
.B(n_2141),
.Y(n_2436)
);

AOI322xp5_ASAP7_75t_L g2437 ( 
.A1(n_2435),
.A2(n_2140),
.A3(n_2151),
.B1(n_2152),
.B2(n_2149),
.C1(n_2162),
.C2(n_2116),
.Y(n_2437)
);

OAI221xp5_ASAP7_75t_R g2438 ( 
.A1(n_2437),
.A2(n_2436),
.B1(n_2208),
.B2(n_2162),
.C(n_2062),
.Y(n_2438)
);

AOI211xp5_ASAP7_75t_L g2439 ( 
.A1(n_2438),
.A2(n_2141),
.B(n_2144),
.C(n_2140),
.Y(n_2439)
);


endmodule