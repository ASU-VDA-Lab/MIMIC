module real_aes_8587_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g257 ( .A1(n_0), .A2(n_258), .B(n_259), .C(n_262), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_1), .B(n_246), .Y(n_263) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_90), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g459 ( .A(n_2), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_3), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_4), .A2(n_135), .B(n_138), .C(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_5), .A2(n_130), .B(n_576), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_6), .A2(n_130), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_7), .B(n_246), .Y(n_582) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_8), .A2(n_165), .B(n_202), .Y(n_201) );
AND2x6_ASAP7_75t_L g135 ( .A(n_9), .B(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_10), .A2(n_135), .B(n_138), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g520 ( .A(n_11), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_12), .B(n_40), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_13), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_13), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_14), .B(n_222), .Y(n_554) );
INVx1_ASAP7_75t_L g156 ( .A(n_15), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_16), .B(n_174), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_17), .A2(n_175), .B(n_538), .C(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_18), .B(n_246), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_19), .B(n_150), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_20), .A2(n_138), .B(n_141), .C(n_149), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_21), .A2(n_210), .B(n_261), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_22), .B(n_222), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_23), .A2(n_56), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_23), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_24), .B(n_222), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g567 ( .A(n_25), .Y(n_567) );
INVx1_ASAP7_75t_L g492 ( .A(n_26), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_27), .A2(n_138), .B(n_149), .C(n_205), .Y(n_204) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_28), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_29), .Y(n_550) );
INVx1_ASAP7_75t_L g508 ( .A(n_30), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_31), .A2(n_130), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_33), .A2(n_178), .B(n_187), .C(n_189), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_34), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_35), .A2(n_261), .B(n_579), .C(n_581), .Y(n_578) );
INVxp67_ASAP7_75t_L g509 ( .A(n_36), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_37), .B(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_38), .A2(n_138), .B(n_149), .C(n_491), .Y(n_490) );
CKINVDCx14_ASAP7_75t_R g577 ( .A(n_39), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_41), .A2(n_262), .B(n_518), .C(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_42), .B(n_129), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_43), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_44), .B(n_174), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_45), .B(n_130), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_46), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_47), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_48), .A2(n_178), .B(n_187), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_49), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g260 ( .A(n_50), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_51), .A2(n_447), .B1(n_448), .B2(n_451), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_51), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_52), .A2(n_465), .B1(n_466), .B2(n_475), .C1(n_755), .C2(n_759), .Y(n_464) );
INVx1_ASAP7_75t_L g232 ( .A(n_53), .Y(n_232) );
INVx1_ASAP7_75t_L g526 ( .A(n_54), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_55), .B(n_130), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_56), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_57), .Y(n_158) );
CKINVDCx14_ASAP7_75t_R g516 ( .A(n_58), .Y(n_516) );
INVx1_ASAP7_75t_L g136 ( .A(n_59), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_60), .B(n_130), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_61), .B(n_246), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_62), .A2(n_148), .B(n_171), .C(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g155 ( .A(n_63), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_64), .A2(n_103), .B1(n_471), .B2(n_472), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_64), .Y(n_472) );
INVx1_ASAP7_75t_SL g580 ( .A(n_65), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_67), .B(n_174), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_68), .B(n_246), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_69), .B(n_175), .Y(n_220) );
INVx1_ASAP7_75t_L g570 ( .A(n_70), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_71), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_72), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_73), .A2(n_138), .B(n_169), .C(n_178), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_74), .Y(n_241) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_76), .A2(n_130), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_77), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_78), .A2(n_130), .B(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_79), .A2(n_129), .B(n_504), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_80), .Y(n_489) );
INVx1_ASAP7_75t_L g536 ( .A(n_81), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_82), .B(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_83), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_84), .A2(n_130), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g539 ( .A(n_85), .Y(n_539) );
INVx2_ASAP7_75t_L g153 ( .A(n_86), .Y(n_153) );
INVx1_ASAP7_75t_L g553 ( .A(n_87), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_88), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_89), .B(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g456 ( .A(n_90), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g478 ( .A(n_90), .B(n_458), .Y(n_478) );
INVx2_ASAP7_75t_L g480 ( .A(n_90), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_91), .A2(n_470), .B1(n_473), .B2(n_474), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_91), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_92), .A2(n_138), .B(n_178), .C(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_93), .B(n_130), .Y(n_185) );
INVx1_ASAP7_75t_L g190 ( .A(n_94), .Y(n_190) );
INVxp67_ASAP7_75t_L g244 ( .A(n_95), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_96), .A2(n_105), .B1(n_114), .B2(n_765), .Y(n_104) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_97), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_97), .B(n_165), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g170 ( .A(n_99), .Y(n_170) );
INVx1_ASAP7_75t_L g216 ( .A(n_100), .Y(n_216) );
INVx2_ASAP7_75t_L g529 ( .A(n_101), .Y(n_529) );
AND2x2_ASAP7_75t_L g234 ( .A(n_102), .B(n_152), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_103), .Y(n_471) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_SL g766 ( .A(n_107), .Y(n_766) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g458 ( .A(n_108), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_117), .B(n_463), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g764 ( .A(n_116), .Y(n_764) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_453), .B(n_460), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_445), .B1(n_446), .B2(n_452), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_120), .A2(n_482), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g452 ( .A(n_121), .Y(n_452) );
AND3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_349), .C(n_406), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_294), .C(n_330), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_196), .B(n_248), .C(n_281), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g251 ( .A(n_126), .B(n_252), .Y(n_251) );
INVx5_ASAP7_75t_L g280 ( .A(n_126), .Y(n_280) );
AND2x2_ASAP7_75t_L g353 ( .A(n_126), .B(n_269), .Y(n_353) );
AND2x2_ASAP7_75t_L g391 ( .A(n_126), .B(n_297), .Y(n_391) );
AND2x2_ASAP7_75t_L g411 ( .A(n_126), .B(n_253), .Y(n_411) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_157), .Y(n_126) );
AOI21xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_137), .B(n_150), .Y(n_127) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_131), .B(n_135), .Y(n_217) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_134), .Y(n_144) );
INVx3_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_134), .Y(n_222) );
BUFx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx4_ASAP7_75t_SL g179 ( .A(n_135), .Y(n_179) );
INVx5_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
BUFx3_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_147), .Y(n_141) );
INVx2_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_146), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_146), .A2(n_192), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_146), .A2(n_553), .B(n_554), .C(n_555), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_146), .A2(n_555), .B(n_570), .C(n_571), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_147), .A2(n_174), .B(n_492), .C(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_148), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_151), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_152), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_152), .A2(n_229), .B(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_217), .B(n_489), .C(n_490), .Y(n_488) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_152), .A2(n_514), .B(n_521), .Y(n_513) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g166 ( .A(n_153), .B(n_154), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_159), .A2(n_549), .B(n_556), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_160), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_183), .Y(n_160) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_161), .Y(n_292) );
AND2x2_ASAP7_75t_L g306 ( .A(n_161), .B(n_252), .Y(n_306) );
INVx1_ASAP7_75t_L g329 ( .A(n_161), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_161), .B(n_280), .Y(n_368) );
OR2x2_ASAP7_75t_L g405 ( .A(n_161), .B(n_250), .Y(n_405) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_162), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_162), .B(n_253), .Y(n_348) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g269 ( .A(n_163), .B(n_253), .Y(n_269) );
BUFx2_ASAP7_75t_L g297 ( .A(n_163), .Y(n_297) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_181), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_164), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_164), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_164), .A2(n_215), .B(n_223), .Y(n_214) );
INVx3_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_164), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_164), .B(n_557), .Y(n_556) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_164), .A2(n_566), .B(n_572), .Y(n_565) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_165), .A2(n_203), .B(n_204), .Y(n_202) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_165), .Y(n_238) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_173), .C(n_176), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_172), .A2(n_174), .B1(n_508), .B2(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_172), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_172), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_174), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g258 ( .A(n_174), .Y(n_258) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_175), .B(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g581 ( .A(n_177), .Y(n_581) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_179), .A2(n_188), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_179), .A2(n_188), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_179), .A2(n_188), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_179), .A2(n_188), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_179), .A2(n_188), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_179), .A2(n_188), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_179), .A2(n_188), .B(n_577), .C(n_578), .Y(n_576) );
INVx5_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
BUFx2_ASAP7_75t_L g273 ( .A(n_183), .Y(n_273) );
AND2x2_ASAP7_75t_L g430 ( .A(n_183), .B(n_284), .Y(n_430) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_194), .Y(n_183) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g262 ( .A(n_193), .Y(n_262) );
INVx1_ASAP7_75t_L g540 ( .A(n_193), .Y(n_540) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_235), .Y(n_197) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_198), .A2(n_331), .B1(n_338), .B2(n_339), .C(n_342), .Y(n_330) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_212), .Y(n_198) );
AND2x2_ASAP7_75t_L g236 ( .A(n_199), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_199), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g265 ( .A(n_200), .B(n_213), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_200), .B(n_214), .Y(n_275) );
OR2x2_ASAP7_75t_L g286 ( .A(n_200), .B(n_237), .Y(n_286) );
AND2x2_ASAP7_75t_L g289 ( .A(n_200), .B(n_277), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_200), .B(n_226), .Y(n_305) );
OR2x2_ASAP7_75t_L g321 ( .A(n_200), .B(n_214), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_200), .B(n_237), .Y(n_383) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_201), .B(n_226), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_201), .B(n_214), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B(n_209), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g299 ( .A(n_212), .B(n_286), .Y(n_299) );
INVx2_ASAP7_75t_L g325 ( .A(n_212), .Y(n_325) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
AND2x2_ASAP7_75t_L g247 ( .A(n_213), .B(n_227), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_213), .B(n_237), .Y(n_304) );
OR2x2_ASAP7_75t_L g315 ( .A(n_213), .B(n_227), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_213), .B(n_277), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_213), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_407) );
INVx5_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_214), .B(n_237), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_217), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_217), .A2(n_567), .B(n_568), .Y(n_566) );
INVx4_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
INVx2_ASAP7_75t_L g518 ( .A(n_222), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g501 ( .A(n_225), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_226), .B(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_226), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g293 ( .A(n_226), .B(n_265), .Y(n_293) );
OR2x2_ASAP7_75t_L g337 ( .A(n_226), .B(n_237), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_226), .B(n_289), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_226), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_226), .B(n_403), .Y(n_402) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_227), .B(n_236), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_227), .A2(n_271), .B(n_274), .C(n_278), .Y(n_270) );
OR2x2_ASAP7_75t_L g308 ( .A(n_227), .B(n_304), .Y(n_308) );
OR2x2_ASAP7_75t_L g344 ( .A(n_227), .B(n_286), .Y(n_344) );
OAI311xp33_ASAP7_75t_L g350 ( .A1(n_227), .A2(n_289), .A3(n_351), .B1(n_354), .C1(n_361), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_227), .B(n_237), .Y(n_401) );
AND2x2_ASAP7_75t_L g409 ( .A(n_227), .B(n_264), .Y(n_409) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_227), .Y(n_427) );
AND2x2_ASAP7_75t_L g444 ( .A(n_227), .B(n_265), .Y(n_444) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_247), .Y(n_235) );
AND2x2_ASAP7_75t_L g272 ( .A(n_236), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g428 ( .A(n_236), .Y(n_428) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g277 ( .A(n_237), .Y(n_277) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
INVxp67_ASAP7_75t_L g359 ( .A(n_237), .Y(n_359) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_245), .Y(n_237) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_238), .A2(n_524), .B(n_530), .Y(n_523) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_238), .A2(n_534), .B(n_541), .Y(n_533) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_238), .A2(n_575), .B(n_582), .Y(n_574) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_246), .A2(n_254), .B(n_263), .Y(n_253) );
AND2x2_ASAP7_75t_L g437 ( .A(n_247), .B(n_285), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_264), .B1(n_266), .B2(n_267), .C(n_270), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_250), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g290 ( .A(n_250), .B(n_280), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_250), .B(n_252), .Y(n_298) );
OR2x2_ASAP7_75t_L g310 ( .A(n_250), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_250), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g352 ( .A(n_250), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_250), .Y(n_372) );
AND2x2_ASAP7_75t_L g424 ( .A(n_250), .B(n_348), .Y(n_424) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_250), .A2(n_301), .A3(n_400), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_251), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g396 ( .A(n_251), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_251), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g284 ( .A(n_252), .B(n_280), .Y(n_284) );
INVx1_ASAP7_75t_L g371 ( .A(n_252), .Y(n_371) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g421 ( .A(n_253), .B(n_280), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_261), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g555 ( .A(n_262), .Y(n_555) );
INVx1_ASAP7_75t_SL g431 ( .A(n_264), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_265), .B(n_336), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_266), .A2(n_378), .B1(n_416), .B2(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_269), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_269), .B(n_290), .Y(n_443) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g413 ( .A(n_272), .B(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_273), .A2(n_332), .B(n_334), .Y(n_331) );
OR2x2_ASAP7_75t_L g339 ( .A(n_273), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g360 ( .A(n_273), .B(n_348), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_273), .B(n_371), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_273), .B(n_411), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g387 ( .A1(n_274), .A2(n_388), .B1(n_393), .B2(n_396), .C(n_397), .Y(n_387) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g364 ( .A(n_275), .B(n_337), .Y(n_364) );
INVx1_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
INVx2_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_280), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g347 ( .A(n_280), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g435 ( .A(n_280), .B(n_405), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B1(n_287), .B2(n_290), .C1(n_291), .C2(n_293), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_284), .A2(n_334), .B1(n_362), .B2(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_284), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OAI21xp33_ASAP7_75t_SL g322 ( .A1(n_293), .A2(n_323), .B(n_326), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_299), .B(n_300), .C(n_322), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_298), .A2(n_301), .B1(n_306), .B2(n_307), .C(n_309), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_298), .B(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g392 ( .A(n_298), .Y(n_392) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
AND2x2_ASAP7_75t_L g394 ( .A(n_303), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g311 ( .A(n_306), .Y(n_311) );
AND2x2_ASAP7_75t_L g317 ( .A(n_306), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_316), .B2(n_319), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_313), .B(n_325), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_314), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g414 ( .A(n_318), .Y(n_414) );
AND2x2_ASAP7_75t_L g433 ( .A(n_318), .B(n_348), .Y(n_433) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_325), .B(n_382), .Y(n_441) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_328), .B(n_396), .Y(n_439) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
BUFx2_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
OAI21xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_345), .B(n_347), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_365), .C(n_387), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_369), .B(n_373), .C(n_376), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_366), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp67_ASAP7_75t_SL g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g395 ( .A(n_375), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B(n_384), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g400 ( .A(n_378), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_402), .B2(n_404), .Y(n_397) );
INVx2_ASAP7_75t_SL g418 ( .A(n_405), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_422), .C(n_434), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_418), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_429), .B2(n_431), .C(n_432), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_423), .A2(n_435), .B(n_436), .C(n_438), .Y(n_434) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_442), .B2(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_452), .A2(n_476), .B1(n_479), .B2(n_481), .Y(n_475) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_456), .Y(n_462) );
NOR2x2_ASAP7_75t_L g761 ( .A(n_457), .B(n_480), .Y(n_761) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g479 ( .A(n_458), .B(n_480), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_460), .B(n_464), .C(n_762), .Y(n_463) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g473 ( .A(n_470), .Y(n_473) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g756 ( .A(n_477), .Y(n_756) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g758 ( .A(n_479), .Y(n_758) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OR5x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_649), .C(n_713), .D(n_729), .E(n_744), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_583), .C(n_610), .D(n_633), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_531), .B(n_542), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g562 ( .A(n_487), .Y(n_562) );
AND2x4_ASAP7_75t_L g596 ( .A(n_487), .B(n_585), .Y(n_596) );
OR2x2_ASAP7_75t_L g606 ( .A(n_487), .B(n_564), .Y(n_606) );
OR2x2_ASAP7_75t_L g652 ( .A(n_487), .B(n_499), .Y(n_652) );
AND2x2_ASAP7_75t_L g666 ( .A(n_487), .B(n_563), .Y(n_666) );
AND2x2_ASAP7_75t_L g709 ( .A(n_487), .B(n_599), .Y(n_709) );
AND2x2_ASAP7_75t_L g716 ( .A(n_487), .B(n_574), .Y(n_716) );
AND2x2_ASAP7_75t_L g735 ( .A(n_487), .B(n_625), .Y(n_735) );
AND2x2_ASAP7_75t_L g753 ( .A(n_487), .B(n_595), .Y(n_753) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g718 ( .A(n_496), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_512), .Y(n_496) );
AND2x2_ASAP7_75t_L g628 ( .A(n_497), .B(n_563), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_497), .B(n_648), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g661 ( .A1(n_497), .A2(n_662), .A3(n_665), .B1(n_667), .B2(n_671), .Y(n_661) );
AND2x2_ASAP7_75t_L g731 ( .A(n_497), .B(n_625), .Y(n_731) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g595 ( .A(n_499), .B(n_564), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_499), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_499), .B(n_584), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_499), .B(n_716), .Y(n_715) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B(n_510), .Y(n_499) );
INVx1_ASAP7_75t_L g600 ( .A(n_500), .Y(n_600) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OA21x2_ASAP7_75t_L g599 ( .A1(n_503), .A2(n_511), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g602 ( .A(n_512), .B(n_546), .Y(n_602) );
AND2x2_ASAP7_75t_L g678 ( .A(n_512), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g750 ( .A(n_512), .Y(n_750) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
OR2x2_ASAP7_75t_L g545 ( .A(n_513), .B(n_523), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_513), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_513), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g609 ( .A(n_513), .Y(n_609) );
AND2x2_ASAP7_75t_L g636 ( .A(n_513), .B(n_523), .Y(n_636) );
BUFx3_ASAP7_75t_L g639 ( .A(n_513), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_513), .B(n_614), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_513), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
AND2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_588), .Y(n_608) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g619 ( .A(n_523), .B(n_533), .Y(n_619) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_523), .Y(n_632) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_532), .B(n_639), .Y(n_689) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g560 ( .A(n_533), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_533), .B(n_608), .C(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g615 ( .A(n_533), .B(n_588), .Y(n_615) );
AND2x2_ASAP7_75t_L g635 ( .A(n_533), .B(n_588), .Y(n_635) );
AND2x2_ASAP7_75t_L g679 ( .A(n_533), .B(n_548), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_558), .B(n_561), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g754 ( .A(n_544), .B(n_679), .Y(n_754) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_545), .A2(n_652), .B1(n_694), .B2(n_696), .Y(n_693) );
OR2x2_ASAP7_75t_L g700 ( .A(n_545), .B(n_615), .Y(n_700) );
OR2x2_ASAP7_75t_L g724 ( .A(n_545), .B(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_545), .B(n_644), .Y(n_737) );
AND2x2_ASAP7_75t_L g630 ( .A(n_546), .B(n_631), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_546), .A2(n_703), .B(n_718), .Y(n_717) );
AOI32xp33_ASAP7_75t_L g738 ( .A1(n_546), .A2(n_628), .A3(n_739), .B1(n_741), .B2(n_742), .Y(n_738) );
OR2x2_ASAP7_75t_L g749 ( .A(n_546), .B(n_750), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g617 ( .A(n_547), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_547), .B(n_631), .Y(n_696) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g588 ( .A(n_548), .Y(n_588) );
AND2x2_ASAP7_75t_L g654 ( .A(n_548), .B(n_619), .Y(n_654) );
AND3x2_ASAP7_75t_L g663 ( .A(n_548), .B(n_559), .C(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g589 ( .A(n_560), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_560), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_560), .B(n_588), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g584 ( .A(n_562), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g624 ( .A(n_562), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g642 ( .A(n_562), .B(n_574), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_564), .Y(n_660) );
OR2x2_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g720 ( .A(n_562), .B(n_648), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_563), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_574), .Y(n_563) );
AND2x2_ASAP7_75t_L g621 ( .A(n_564), .B(n_599), .Y(n_621) );
OR2x2_ASAP7_75t_L g675 ( .A(n_564), .B(n_599), .Y(n_675) );
AND2x2_ASAP7_75t_L g728 ( .A(n_564), .B(n_585), .Y(n_728) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
AND2x2_ASAP7_75t_L g648 ( .A(n_565), .B(n_574), .Y(n_648) );
INVx2_ASAP7_75t_L g585 ( .A(n_574), .Y(n_585) );
INVx1_ASAP7_75t_L g605 ( .A(n_574), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .B(n_591), .C(n_603), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_584), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g747 ( .A(n_584), .Y(n_747) );
AND2x2_ASAP7_75t_L g625 ( .A(n_585), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_588), .B(n_589), .Y(n_597) );
INVx1_ASAP7_75t_L g682 ( .A(n_588), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_588), .B(n_609), .Y(n_706) );
AND2x2_ASAP7_75t_L g722 ( .A(n_588), .B(n_636), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_589), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g613 ( .A(n_590), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_594), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_595), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g620 ( .A(n_596), .B(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_SL g685 ( .A1(n_596), .A2(n_638), .B1(n_686), .B2(n_691), .C(n_693), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_596), .B(n_659), .Y(n_692) );
INVx1_ASAP7_75t_L g752 ( .A(n_598), .Y(n_752) );
BUFx3_ASAP7_75t_L g659 ( .A(n_599), .Y(n_659) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_605), .B(n_659), .Y(n_712) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_606), .B(n_659), .Y(n_670) );
INVxp67_ASAP7_75t_L g690 ( .A(n_608), .Y(n_690) );
AND2x2_ASAP7_75t_L g631 ( .A(n_609), .B(n_632), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_616), .B(n_620), .C(n_622), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_SL g645 ( .A(n_613), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_614), .B(n_645), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_614), .B(n_636), .Y(n_687) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_617), .A2(n_623), .B1(n_627), .B2(n_629), .Y(n_622) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g638 ( .A(n_619), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g683 ( .A(n_619), .B(n_684), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_621), .A2(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_625), .A2(n_634), .B1(n_637), .B2(n_638), .C(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_625), .B(n_659), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_625), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g741 ( .A(n_631), .Y(n_741) );
INVxp67_ASAP7_75t_L g664 ( .A(n_632), .Y(n_664) );
INVx1_ASAP7_75t_L g671 ( .A(n_634), .Y(n_671) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g710 ( .A(n_635), .B(n_639), .Y(n_710) );
INVx1_ASAP7_75t_L g684 ( .A(n_639), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_639), .B(n_654), .Y(n_714) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .A3(n_645), .B1(n_646), .B2(n_647), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g653 ( .A(n_648), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_648), .B(n_680), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_648), .B(n_709), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_648), .B(n_659), .Y(n_748) );
NAND5xp2_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .C(n_685), .D(n_697), .E(n_698), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_655), .B2(n_657), .C(n_661), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g676 ( .A(n_656), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_659), .B(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_660), .A2(n_673), .B1(n_676), .B2(n_680), .Y(n_672) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_663), .A2(n_668), .B(n_669), .C(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g695 ( .A(n_675), .Y(n_695) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_684), .B(n_733), .Y(n_743) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_703), .B2(n_707), .C1(n_710), .C2(n_711), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_726), .Y(n_721) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g733 ( .A(n_725), .Y(n_733) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_734), .B2(n_736), .C(n_738), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_749), .C(n_751), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B(n_754), .Y(n_751) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
endmodule