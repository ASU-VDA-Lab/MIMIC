module real_jpeg_4624_n_19 (n_17, n_8, n_116, n_0, n_2, n_10, n_114, n_9, n_12, n_6, n_121, n_11, n_14, n_120, n_7, n_117, n_18, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_16, n_15, n_13, n_113, n_19);

input n_17;
input n_8;
input n_116;
input n_0;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_120;
input n_7;
input n_117;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_1),
.B(n_34),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_2),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_4),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_5),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_94),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_7),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_8),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_48),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_13),
.B(n_38),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_14),
.B(n_44),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_15),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_17),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_18),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_18),
.B(n_107),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_111),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_50),
.B(n_97),
.C(n_106),
.Y(n_31)
);

NOR4xp25_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.C(n_43),
.D(n_47),
.Y(n_32)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_79),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_93),
.B(n_96),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_85),
.B(n_92),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_61),
.B1(n_82),
.B2(n_83),
.C(n_84),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_81),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_77),
.B(n_80),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B(n_76),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_91),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_103),
.C(n_104),
.D(n_105),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_113),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_114),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_115),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_116),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_117),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_118),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_119),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_120),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_121),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_122),
.Y(n_95)
);


endmodule