module real_aes_15894_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_147;
wire n_150;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_0), .Y(n_228) );
AND2x4_ASAP7_75t_L g879 ( .A(n_1), .B(n_880), .Y(n_879) );
BUFx3_ASAP7_75t_L g169 ( .A(n_2), .Y(n_169) );
INVx1_ASAP7_75t_L g880 ( .A(n_3), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_4), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g859 ( .A(n_4), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_5), .B(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g110 ( .A(n_6), .B(n_20), .Y(n_110) );
BUFx2_ASAP7_75t_L g875 ( .A(n_6), .Y(n_875) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_7), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_8), .B(n_163), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_9), .B(n_163), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_10), .B(n_188), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_11), .A2(n_79), .B1(n_138), .B2(n_163), .Y(n_237) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_12), .A2(n_34), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_13), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_14), .B(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_15), .Y(n_524) );
AO32x2_ASAP7_75t_L g234 ( .A1(n_16), .A2(n_155), .A3(n_156), .B1(n_235), .B2(n_238), .Y(n_234) );
AO32x1_ASAP7_75t_L g272 ( .A1(n_16), .A2(n_155), .A3(n_156), .B1(n_235), .B2(n_238), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_17), .B(n_509), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_18), .B(n_155), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_19), .Y(n_537) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_20), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_21), .A2(n_40), .B1(n_166), .B2(n_178), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_22), .A2(n_87), .B1(n_138), .B2(n_146), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_23), .B(n_145), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_24), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_25), .B(n_201), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_26), .A2(n_59), .B1(n_146), .B2(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_27), .B(n_163), .Y(n_579) );
INVx2_ASAP7_75t_L g844 ( .A(n_28), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_29), .B(n_142), .Y(n_610) );
INVx1_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
BUFx3_ASAP7_75t_L g847 ( .A(n_30), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_31), .A2(n_100), .B1(n_869), .B2(n_881), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_32), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_33), .B(n_515), .Y(n_616) );
AND2x2_ASAP7_75t_L g530 ( .A(n_35), .B(n_515), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_36), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_37), .B(n_200), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_38), .B(n_509), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_39), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_41), .B(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_42), .A2(n_73), .B1(n_200), .B2(n_201), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_43), .B(n_243), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_44), .A2(n_179), .B(n_226), .C(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_45), .A2(n_75), .B1(n_138), .B2(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g134 ( .A(n_46), .Y(n_134) );
AND2x4_ASAP7_75t_L g152 ( .A(n_47), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_48), .A2(n_49), .B1(n_146), .B2(n_166), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_50), .B(n_155), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_51), .B(n_515), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_52), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_53), .B(n_146), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_54), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g153 ( .A(n_55), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_56), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_57), .A2(n_226), .B(n_227), .C(n_229), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g150 ( .A(n_58), .B(n_138), .C(n_148), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_60), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_61), .B(n_155), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_62), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g231 ( .A(n_63), .B(n_232), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_64), .Y(n_247) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_65), .B(n_142), .C(n_178), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_66), .A2(n_91), .B1(n_163), .B2(n_200), .Y(n_204) );
INVx2_ASAP7_75t_L g143 ( .A(n_67), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_68), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_69), .B(n_507), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_70), .B(n_163), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_71), .B(n_203), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_72), .A2(n_849), .B1(n_860), .B2(n_864), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_74), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_76), .B(n_182), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_77), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_78), .A2(n_86), .B1(n_509), .B2(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_80), .B(n_163), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_81), .B(n_148), .Y(n_147) );
NAND2xp33_ASAP7_75t_SL g553 ( .A(n_82), .B(n_141), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_83), .B(n_176), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_84), .A2(n_98), .B1(n_146), .B2(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_85), .B(n_201), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g112 ( .A1(n_88), .A2(n_113), .B1(n_838), .B2(n_839), .Y(n_112) );
INVx1_ASAP7_75t_SL g839 ( .A(n_88), .Y(n_839) );
INVx1_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_89), .B(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_90), .B(n_188), .Y(n_264) );
NAND2xp33_ASAP7_75t_L g562 ( .A(n_92), .B(n_141), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_93), .B(n_515), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_94), .B(n_141), .C(n_203), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_95), .B(n_507), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_96), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_97), .B(n_509), .Y(n_512) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_111), .Y(n_100) );
AOI31xp33_ASAP7_75t_L g858 ( .A1(n_101), .A2(n_119), .A3(n_851), .B(n_859), .Y(n_858) );
NOR2x1_ASAP7_75t_SL g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx4_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND3x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .C(n_109), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_105), .B(n_877), .Y(n_876) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g855 ( .A(n_106), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_107), .B(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g117 ( .A(n_108), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_109), .B(n_846), .Y(n_845) );
AND2x6_ASAP7_75t_SL g853 ( .A(n_109), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_L g868 ( .A(n_110), .B(n_847), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_840), .B(n_848), .Y(n_111) );
INVx1_ASAP7_75t_L g838 ( .A(n_113), .Y(n_838) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_494), .Y(n_113) );
INVx8_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx12f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
BUFx8_ASAP7_75t_SL g837 ( .A(n_117), .Y(n_837) );
AND2x2_ASAP7_75t_L g867 ( .A(n_117), .B(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g857 ( .A(n_118), .Y(n_857) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_404), .Y(n_119) );
NAND4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_309), .C(n_336), .D(n_372), .Y(n_120) );
AOI221x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_214), .B1(n_248), .B2(n_284), .C(n_288), .Y(n_121) );
NAND3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_190), .C(n_212), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_157), .Y(n_125) );
INVx2_ASAP7_75t_L g249 ( .A(n_126), .Y(n_249) );
AND2x2_ASAP7_75t_L g422 ( .A(n_126), .B(n_366), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_126), .B(n_213), .Y(n_431) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g437 ( .A(n_127), .Y(n_437) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g282 ( .A(n_128), .Y(n_282) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g365 ( .A(n_129), .B(n_211), .Y(n_365) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B(n_154), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_130), .A2(n_135), .B(n_154), .Y(n_294) );
OAI21x1_ASAP7_75t_L g503 ( .A1(n_130), .A2(n_504), .B(n_514), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_130), .A2(n_535), .B(n_543), .Y(n_534) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_130), .A2(n_535), .B(n_543), .Y(n_633) );
OAI21xp33_ASAP7_75t_SL g724 ( .A1(n_130), .A2(n_504), .B(n_514), .Y(n_724) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g515 ( .A(n_131), .Y(n_515) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
INVx2_ASAP7_75t_L g209 ( .A(n_132), .Y(n_209) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_133), .Y(n_156) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_144), .B(n_151), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B(n_142), .Y(n_136) );
INVx2_ASAP7_75t_SL g201 ( .A(n_138), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_138), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_139), .Y(n_141) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx1_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx1_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
INVx1_ASAP7_75t_L g226 ( .A(n_139), .Y(n_226) );
INVx3_ASAP7_75t_L g507 ( .A(n_139), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_139), .Y(n_510) );
INVx2_ASAP7_75t_L g542 ( .A(n_141), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_142), .A2(n_162), .B1(n_164), .B2(n_165), .Y(n_161) );
INVx6_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_142), .A2(n_179), .B1(n_236), .B2(n_237), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_L g536 ( .A1(n_142), .A2(n_175), .B(n_537), .C(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_142), .A2(n_581), .B(n_582), .Y(n_580) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_150), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_146), .A2(n_507), .B1(n_528), .B2(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g587 ( .A(n_146), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_146), .A2(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
AOI31xp67_ASAP7_75t_L g159 ( .A1(n_151), .A2(n_160), .A3(n_161), .B(n_167), .Y(n_159) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_173), .B(n_180), .Y(n_172) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_151), .A2(n_505), .B(n_511), .Y(n_504) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_151), .A2(n_536), .B(n_539), .Y(n_535) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_151), .A2(n_548), .B(n_551), .Y(n_547) );
AND2x4_ASAP7_75t_SL g567 ( .A(n_151), .B(n_156), .Y(n_567) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_151), .A2(n_577), .B(n_580), .Y(n_576) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_151), .A2(n_609), .B(n_612), .Y(n_608) );
BUFx10_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_152), .A2(n_197), .A3(n_241), .B(n_246), .Y(n_240) );
BUFx10_ASAP7_75t_L g520 ( .A(n_152), .Y(n_520) );
INVx2_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_156), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
BUFx3_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_156), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_SL g255 ( .A(n_156), .Y(n_255) );
INVx1_ASAP7_75t_SL g546 ( .A(n_156), .Y(n_546) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_157), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_157), .B(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g435 ( .A(n_157), .Y(n_435) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_170), .Y(n_157) );
AND2x2_ASAP7_75t_L g213 ( .A(n_158), .B(n_196), .Y(n_213) );
INVx2_ASAP7_75t_L g291 ( .A(n_158), .Y(n_291) );
AND2x2_ASAP7_75t_L g356 ( .A(n_158), .B(n_294), .Y(n_356) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
INVx3_ASAP7_75t_L g263 ( .A(n_163), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_163), .A2(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g615 ( .A(n_163), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_199), .B1(n_202), .B2(n_204), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_164), .A2(n_242), .B1(n_244), .B2(n_245), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_164), .A2(n_261), .B(n_262), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_164), .A2(n_526), .B1(n_586), .B2(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g185 ( .A(n_166), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_166), .A2(n_178), .B1(n_222), .B2(n_223), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g283 ( .A(n_170), .Y(n_283) );
AND2x2_ASAP7_75t_L g293 ( .A(n_170), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g355 ( .A(n_170), .B(n_196), .Y(n_355) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_187), .Y(n_170) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_171), .A2(n_172), .B(n_187), .Y(n_193) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_171), .A2(n_576), .B(n_583), .Y(n_575) );
OAI21x1_ASAP7_75t_L g607 ( .A1(n_171), .A2(n_608), .B(n_616), .Y(n_607) );
OA21x2_ASAP7_75t_L g619 ( .A1(n_171), .A2(n_608), .B(n_616), .Y(n_619) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_171), .A2(n_576), .B(n_583), .Y(n_622) );
O2A1O1Ixp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_177), .C(n_179), .Y(n_173) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_179), .A2(n_506), .B(n_508), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_179), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_179), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_179), .A2(n_578), .B(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B1(n_185), .B2(n_186), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_182), .A2(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_183), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx3_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
INVx2_ASAP7_75t_L g218 ( .A(n_188), .Y(n_218) );
NOR2xp67_ASAP7_75t_SL g518 ( .A(n_188), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_189), .A2(n_520), .A3(n_585), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g320 ( .A(n_190), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_192), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_192), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_192), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_192), .B(n_390), .Y(n_397) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g366 ( .A(n_193), .B(n_341), .Y(n_366) );
OR2x2_ASAP7_75t_L g368 ( .A(n_193), .B(n_294), .Y(n_368) );
INVx1_ASAP7_75t_L g427 ( .A(n_193), .Y(n_427) );
BUFx2_ASAP7_75t_L g441 ( .A(n_193), .Y(n_441) );
OR2x2_ASAP7_75t_L g469 ( .A(n_193), .B(n_196), .Y(n_469) );
INVx1_ASAP7_75t_L g488 ( .A(n_194), .Y(n_488) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g335 ( .A(n_195), .Y(n_335) );
OR2x2_ASAP7_75t_L g348 ( .A(n_195), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g367 ( .A(n_195), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
INVx2_ASAP7_75t_L g287 ( .A(n_196), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_196), .B(n_210), .Y(n_303) );
INVx1_ASAP7_75t_L g341 ( .A(n_196), .Y(n_341) );
INVx1_ASAP7_75t_L g384 ( .A(n_196), .Y(n_384) );
AND2x2_ASAP7_75t_L g426 ( .A(n_196), .B(n_427), .Y(n_426) );
AO31x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .A3(n_205), .B(n_207), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_200), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g224 ( .A(n_203), .Y(n_224) );
INVx2_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_SL g238 ( .A(n_206), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx2_ASAP7_75t_L g232 ( .A(n_209), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_209), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g482 ( .A(n_212), .Y(n_482) );
AND2x4_ASAP7_75t_L g420 ( .A(n_213), .B(n_280), .Y(n_420) );
INVx2_ASAP7_75t_L g449 ( .A(n_213), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_213), .B(n_441), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_214), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_233), .Y(n_214) );
AND2x2_ASAP7_75t_L g360 ( .A(n_215), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g381 ( .A(n_215), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g252 ( .A(n_216), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g276 ( .A(n_216), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g307 ( .A(n_216), .Y(n_307) );
AND2x2_ASAP7_75t_L g347 ( .A(n_216), .B(n_239), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_216), .B(n_331), .Y(n_388) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g300 ( .A(n_217), .Y(n_300) );
AOI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_231), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_225), .B(n_230), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_224), .Y(n_220) );
AOI21x1_ASAP7_75t_L g612 ( .A1(n_224), .A2(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g565 ( .A(n_226), .Y(n_565) );
INVx2_ASAP7_75t_L g245 ( .A(n_229), .Y(n_245) );
INVx2_ASAP7_75t_L g526 ( .A(n_229), .Y(n_526) );
INVx3_ASAP7_75t_L g266 ( .A(n_233), .Y(n_266) );
AND2x2_ASAP7_75t_L g311 ( .A(n_233), .B(n_306), .Y(n_311) );
AND2x2_ASAP7_75t_L g466 ( .A(n_233), .B(n_270), .Y(n_466) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_239), .Y(n_233) );
INVx1_ASAP7_75t_L g317 ( .A(n_234), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_234), .B(n_253), .Y(n_345) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_238), .A2(n_257), .B(n_260), .Y(n_256) );
AND2x4_ASAP7_75t_L g298 ( .A(n_239), .B(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g271 ( .A(n_240), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g308 ( .A(n_240), .B(n_272), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_240), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_240), .B(n_253), .Y(n_370) );
AND2x2_ASAP7_75t_L g376 ( .A(n_240), .B(n_300), .Y(n_376) );
AOI21x1_ASAP7_75t_L g257 ( .A1(n_245), .A2(n_258), .B(n_259), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_245), .A2(n_512), .B(n_513), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_267), .Y(n_248) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_249), .A2(n_410), .B(n_414), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_249), .B(n_440), .Y(n_487) );
NAND2x1_ASAP7_75t_SL g250 ( .A(n_251), .B(n_265), .Y(n_250) );
INVx1_ASAP7_75t_L g493 ( .A(n_251), .Y(n_493) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g270 ( .A(n_253), .Y(n_270) );
INVx2_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
INVxp67_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
AND2x2_ASAP7_75t_L g316 ( .A(n_253), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g327 ( .A(n_253), .B(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g331 ( .A(n_253), .Y(n_331) );
INVx1_ASAP7_75t_L g349 ( .A(n_253), .Y(n_349) );
OR2x2_ASAP7_75t_L g382 ( .A(n_253), .B(n_317), .Y(n_382) );
INVx1_ASAP7_75t_L g453 ( .A(n_253), .Y(n_453) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_264), .Y(n_254) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_273), .B(n_278), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_269), .A2(n_392), .B1(n_394), .B2(n_397), .Y(n_391) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_270), .B(n_318), .Y(n_352) );
BUFx2_ASAP7_75t_L g411 ( .A(n_270), .Y(n_411) );
INVx2_ASAP7_75t_L g361 ( .A(n_271), .Y(n_361) );
OR2x2_ASAP7_75t_L g445 ( .A(n_271), .B(n_275), .Y(n_445) );
INVx1_ASAP7_75t_L g277 ( .A(n_272), .Y(n_277) );
INVx1_ASAP7_75t_L g326 ( .A(n_272), .Y(n_326) );
NOR2x1p5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_275), .Y(n_396) );
OR2x2_ASAP7_75t_L g480 ( .A(n_275), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g483 ( .A(n_275), .B(n_318), .Y(n_483) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_276), .Y(n_446) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_280), .B(n_340), .Y(n_402) );
AND2x2_ASAP7_75t_L g492 ( .A(n_280), .B(n_290), .Y(n_492) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g401 ( .A(n_281), .B(n_290), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g358 ( .A(n_282), .B(n_291), .Y(n_358) );
AND2x2_ASAP7_75t_L g393 ( .A(n_282), .B(n_287), .Y(n_393) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_293), .Y(n_312) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g452 ( .A(n_287), .B(n_453), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_295), .B1(n_301), .B2(n_304), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_289), .A2(n_490), .B(n_491), .C(n_493), .Y(n_489) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g340 ( .A(n_291), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g408 ( .A(n_291), .Y(n_408) );
OR2x2_ASAP7_75t_L g455 ( .A(n_292), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g310 ( .A(n_296), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g413 ( .A(n_299), .Y(n_413) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
INVx1_ASAP7_75t_L g400 ( .A(n_300), .Y(n_400) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g456 ( .A(n_303), .Y(n_456) );
AND2x2_ASAP7_75t_L g478 ( .A(n_303), .B(n_441), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_304), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g330 ( .A(n_308), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g386 ( .A(n_308), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g481 ( .A(n_308), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_313), .B2(n_320), .C(n_321), .Y(n_309) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx2_ASAP7_75t_L g403 ( .A(n_316), .Y(n_403) );
BUFx2_ASAP7_75t_L g423 ( .A(n_318), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_329), .B(n_332), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
AND2x2_ASAP7_75t_L g465 ( .A(n_324), .B(n_387), .Y(n_465) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
AND2x2_ASAP7_75t_L g461 ( .A(n_326), .B(n_331), .Y(n_461) );
INVx1_ASAP7_75t_L g344 ( .A(n_328), .Y(n_344) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_350), .C(n_362), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_346), .B2(n_348), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
BUFx2_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
AND2x2_ASAP7_75t_L g471 ( .A(n_345), .B(n_413), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_346), .A2(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B1(n_357), .B2(n_359), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_353), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g425 ( .A(n_358), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g412 ( .A(n_361), .B(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_361), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B(n_369), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
AND2x2_ASAP7_75t_L g439 ( .A(n_364), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g476 ( .A(n_364), .B(n_441), .Y(n_476) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
OR2x2_ASAP7_75t_L g468 ( .A(n_365), .B(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g383 ( .A(n_368), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
OR2x2_ASAP7_75t_L g448 ( .A(n_368), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_391), .C(n_398), .Y(n_372) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .A3(n_379), .B1(n_381), .B2(n_383), .C1(n_385), .C2(n_389), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_375), .A2(n_415), .B(n_451), .C(n_454), .Y(n_450) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_376), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g432 ( .A(n_376), .Y(n_432) );
AND2x4_ASAP7_75t_L g460 ( .A(n_376), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g429 ( .A1(n_378), .A2(n_416), .A3(n_430), .B1(n_432), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_384), .B(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_402), .C(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_405), .B(n_462), .Y(n_404) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_417), .C(n_442), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_410), .A2(n_485), .B(n_486), .C(n_488), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g464 ( .A1(n_412), .A2(n_465), .A3(n_466), .B(n_467), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
NAND4xp25_ASAP7_75t_SL g417 ( .A(n_418), .B(n_421), .C(n_429), .D(n_438), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AOI32xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .A3(n_424), .B1(n_425), .B2(n_428), .Y(n_421) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g485 ( .A(n_428), .Y(n_485) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_450), .C(n_457), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_446), .B(n_447), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_451), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_474), .C(n_484), .D(n_489), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_470), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_465), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_482), .B2(n_483), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_481), .Y(n_490) );
INVxp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_837), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_496), .B(n_732), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_497), .B(n_667), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_591), .C(n_640), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_531), .B(n_555), .C(n_572), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g806 ( .A(n_500), .B(n_725), .Y(n_806) );
OR2x2_ASAP7_75t_L g817 ( .A(n_500), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_501), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g708 ( .A(n_501), .B(n_598), .Y(n_708) );
AND2x2_ASAP7_75t_L g829 ( .A(n_501), .B(n_639), .Y(n_829) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_516), .Y(n_501) );
INVx2_ASAP7_75t_L g659 ( .A(n_502), .Y(n_659) );
AND2x2_ASAP7_75t_L g674 ( .A(n_502), .B(n_626), .Y(n_674) );
AND2x2_ASAP7_75t_L g683 ( .A(n_502), .B(n_557), .Y(n_683) );
AND2x2_ASAP7_75t_L g752 ( .A(n_502), .B(n_638), .Y(n_752) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g723 ( .A(n_516), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g571 ( .A(n_517), .B(n_545), .Y(n_571) );
INVx2_ASAP7_75t_L g596 ( .A(n_517), .Y(n_596) );
AOI21x1_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .B(n_530), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g760 ( .A(n_531), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_544), .Y(n_532) );
INVx1_ASAP7_75t_L g780 ( .A(n_533), .Y(n_780) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g618 ( .A(n_534), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g701 ( .A(n_534), .B(n_607), .Y(n_701) );
AND2x2_ASAP7_75t_L g627 ( .A(n_544), .B(n_570), .Y(n_627) );
INVxp67_ASAP7_75t_L g776 ( .A(n_544), .Y(n_776) );
OR2x2_ASAP7_75t_L g818 ( .A(n_544), .B(n_557), .Y(n_818) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_554), .Y(n_545) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_568), .Y(n_555) );
INVx1_ASAP7_75t_L g673 ( .A(n_556), .Y(n_673) );
AND2x2_ASAP7_75t_L g827 ( .A(n_556), .B(n_723), .Y(n_827) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g599 ( .A(n_557), .Y(n_599) );
INVx4_ASAP7_75t_L g638 ( .A(n_557), .Y(n_638) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B(n_567), .Y(n_559) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g654 ( .A(n_569), .B(n_637), .Y(n_654) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g691 ( .A(n_570), .B(n_639), .Y(n_691) );
INVx2_ASAP7_75t_L g657 ( .A(n_571), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_571), .B(n_662), .Y(n_825) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_574), .B(n_738), .Y(n_737) );
BUFx2_ASAP7_75t_L g810 ( .A(n_574), .Y(n_810) );
AND2x2_ASAP7_75t_L g824 ( .A(n_574), .B(n_646), .Y(n_824) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_584), .Y(n_574) );
INVx1_ASAP7_75t_L g605 ( .A(n_575), .Y(n_605) );
AND2x2_ASAP7_75t_L g759 ( .A(n_575), .B(n_666), .Y(n_759) );
OR2x2_ASAP7_75t_L g796 ( .A(n_575), .B(n_584), .Y(n_796) );
AND2x2_ASAP7_75t_L g606 ( .A(n_584), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g620 ( .A(n_584), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
OR2x2_ASAP7_75t_L g679 ( .A(n_584), .B(n_619), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_584), .B(n_619), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_601), .B(n_623), .Y(n_591) );
INVxp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI31xp33_ASAP7_75t_L g669 ( .A1(n_593), .A2(n_670), .A3(n_672), .B(n_675), .Y(n_669) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
AND2x2_ASAP7_75t_L g682 ( .A(n_594), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g692 ( .A(n_595), .Y(n_692) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_595), .Y(n_698) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g626 ( .A(n_596), .Y(n_626) );
AND2x2_ASAP7_75t_L g655 ( .A(n_596), .B(n_639), .Y(n_655) );
INVx2_ASAP7_75t_L g705 ( .A(n_596), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_597), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g730 ( .A(n_598), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g779 ( .A(n_598), .B(n_780), .Y(n_779) );
AOI33xp33_ASAP7_75t_L g834 ( .A1(n_598), .A2(n_664), .A3(n_674), .B1(n_701), .B2(n_810), .B3(n_835), .Y(n_834) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
INVx1_ASAP7_75t_L g726 ( .A(n_600), .Y(n_726) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_617), .Y(n_602) );
INVx2_ASAP7_75t_L g634 ( .A(n_603), .Y(n_634) );
AND2x2_ASAP7_75t_L g715 ( .A(n_603), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g677 ( .A(n_604), .Y(n_677) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g745 ( .A(n_605), .B(n_632), .Y(n_745) );
AND2x2_ASAP7_75t_L g695 ( .A(n_606), .B(n_689), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_606), .B(n_713), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_606), .B(n_745), .Y(n_794) );
AND2x2_ASAP7_75t_L g631 ( .A(n_607), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g650 ( .A(n_607), .B(n_645), .Y(n_650) );
INVx1_ASAP7_75t_L g665 ( .A(n_607), .Y(n_665) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g720 ( .A(n_618), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_618), .B(n_813), .Y(n_815) );
AND2x2_ASAP7_75t_L g828 ( .A(n_618), .B(n_644), .Y(n_828) );
AND2x2_ASAP7_75t_L g646 ( .A(n_619), .B(n_632), .Y(n_646) );
INVx2_ASAP7_75t_L g628 ( .A(n_620), .Y(n_628) );
AND2x2_ASAP7_75t_L g742 ( .A(n_620), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g801 ( .A(n_620), .B(n_713), .Y(n_801) );
BUFx2_ASAP7_75t_L g783 ( .A(n_621), .Y(n_783) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx3_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
OAI32xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_628), .A3(n_629), .B1(n_634), .B2(n_635), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_L g731 ( .A(n_626), .Y(n_731) );
AND2x2_ASAP7_75t_L g761 ( .A(n_626), .B(n_683), .Y(n_761) );
AND2x2_ASAP7_75t_L g703 ( .A(n_627), .B(n_704), .Y(n_703) );
AND3x2_ASAP7_75t_L g710 ( .A(n_627), .B(n_637), .C(n_705), .Y(n_710) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_630), .A2(n_652), .B1(n_661), .B2(n_663), .Y(n_660) );
OAI322xp33_ASAP7_75t_L g808 ( .A1(n_630), .A2(n_729), .A3(n_809), .B1(n_810), .B2(n_811), .C1(n_812), .C2(n_815), .Y(n_808) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g830 ( .A(n_631), .B(n_813), .Y(n_830) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_632), .Y(n_649) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_632), .Y(n_689) );
BUFx3_ASAP7_75t_L g713 ( .A(n_632), .Y(n_713) );
INVx1_ASAP7_75t_L g739 ( .A(n_632), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_632), .Y(n_743) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g697 ( .A(n_636), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g748 ( .A(n_637), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g799 ( .A(n_637), .B(n_705), .Y(n_799) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_638), .B(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g662 ( .A(n_638), .Y(n_662) );
AND2x2_ASAP7_75t_L g704 ( .A(n_638), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g725 ( .A(n_638), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_639), .B(n_752), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_647), .B(n_651), .C(n_660), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI31xp33_ASAP7_75t_L g802 ( .A1(n_642), .A2(n_803), .A3(n_805), .B(n_806), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
AND2x4_ASAP7_75t_L g755 ( .A(n_643), .B(n_664), .Y(n_755) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_644), .Y(n_687) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp67_ASAP7_75t_L g771 ( .A(n_645), .B(n_665), .Y(n_771) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .Y(n_651) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g811 ( .A(n_654), .Y(n_811) );
AND2x2_ASAP7_75t_L g671 ( .A(n_655), .B(n_662), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_656), .A2(n_741), .B1(n_744), .B2(n_746), .Y(n_740) );
OR2x6_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_SL g798 ( .A(n_659), .Y(n_798) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g768 ( .A(n_664), .B(n_713), .Y(n_768) );
INVx2_ASAP7_75t_L g814 ( .A(n_664), .Y(n_814) );
AND2x4_ASAP7_75t_L g822 ( .A(n_664), .B(n_743), .Y(n_822) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_684), .C(n_714), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_680), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_671), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AND2x4_ASAP7_75t_L g735 ( .A(n_673), .B(n_690), .Y(n_735) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_676), .B(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_L g766 ( .A(n_678), .B(n_745), .Y(n_766) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_679), .Y(n_686) );
INVx1_ASAP7_75t_L g804 ( .A(n_679), .Y(n_804) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g833 ( .A(n_682), .Y(n_833) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_683), .Y(n_718) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_690), .B(n_693), .C(n_706), .Y(n_684) );
NOR3x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .Y(n_685) );
NAND2x1_ASAP7_75t_L g754 ( .A(n_688), .B(n_755), .Y(n_754) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2x1p5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_692), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_699), .B2(n_702), .Y(n_693) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g787 ( .A(n_698), .Y(n_787) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g782 ( .A(n_701), .B(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g836 ( .A(n_704), .Y(n_836) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_711), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g790 ( .A(n_711), .Y(n_790) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx2_ASAP7_75t_L g717 ( .A(n_713), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_713), .B(n_771), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_719), .Y(n_714) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_717), .B(n_804), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_727), .B2(n_729), .Y(n_719) );
OR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g772 ( .A(n_722), .Y(n_772) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g747 ( .A(n_723), .B(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g764 ( .A(n_724), .Y(n_764) );
INVx1_ASAP7_75t_L g784 ( .A(n_725), .Y(n_784) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_788), .Y(n_732) );
NAND3xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_749), .C(n_762), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_740), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g795 ( .A(n_738), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_747), .B(n_775), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B1(n_756), .B2(n_760), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g805 ( .A(n_755), .Y(n_805) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI21xp33_ASAP7_75t_L g777 ( .A1(n_757), .A2(n_778), .B(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_773), .B1(n_777), .B2(n_785), .Y(n_762) );
OAI21xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B(n_767), .Y(n_763) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g832 ( .A(n_768), .Y(n_832) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g821 ( .A(n_771), .Y(n_821) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
INVx2_ASAP7_75t_L g813 ( .A(n_783), .Y(n_813) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_807), .Y(n_788) );
AOI211xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B(n_793), .C(n_802), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_795), .B(n_797), .C(n_800), .Y(n_793) );
OR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_816), .C(n_831), .Y(n_807) );
OR2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
OAI221xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .B1(n_823), .B2(n_825), .C(n_826), .Y(n_816) );
NOR2xp67_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_828), .B1(n_829), .B2(n_830), .Y(n_826) );
OAI21xp33_ASAP7_75t_SL g831 ( .A1(n_832), .A2(n_833), .B(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
BUFx12f_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AND2x6_ASAP7_75t_SL g842 ( .A(n_843), .B(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx3_ASAP7_75t_L g863 ( .A(n_844), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_844), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI21x1_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_856), .B(n_858), .Y(n_849) );
INVx5_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
CKINVDCx11_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx10_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx3_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OR2x6_ASAP7_75t_L g870 ( .A(n_871), .B(n_876), .Y(n_870) );
OR2x6_ASAP7_75t_L g883 ( .A(n_871), .B(n_876), .Y(n_883) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR2x1p5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
CKINVDCx6p67_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
CKINVDCx12_ASAP7_75t_R g882 ( .A(n_883), .Y(n_882) );
endmodule