module fake_netlist_6_4948_n_1713 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1713);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1713;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_12),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_26),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_21),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_89),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_26),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_1),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_118),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_39),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_58),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_61),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_51),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_22),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_50),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_11),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_34),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_36),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_16),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_8),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_53),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_101),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_81),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_85),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_42),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_35),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_123),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_27),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_88),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_32),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_20),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_14),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_80),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_152),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_106),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_105),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_90),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_71),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_69),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_56),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_87),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_149),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_70),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_134),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_109),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_5),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_76),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_74),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_114),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_57),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_28),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_13),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_84),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_77),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_29),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_145),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_31),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_16),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_147),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_68),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_31),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_29),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_27),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_120),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_92),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_122),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_97),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_127),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_82),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_65),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_5),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_42),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_72),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_4),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_143),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_17),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_47),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_47),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_124),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_132),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_136),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_55),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_91),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_12),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_24),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_11),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_168),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_289),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_191),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_160),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_168),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_192),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_168),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_255),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_193),
.B(n_0),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_168),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_287),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_181),
.B(n_2),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_200),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_R g325 ( 
.A(n_164),
.B(n_6),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_171),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_198),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_226),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_200),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_205),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_170),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_203),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_200),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_208),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_193),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_159),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_212),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_179),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_213),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_214),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_216),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_156),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_221),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_222),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

BUFx6f_ASAP7_75t_SL g353 ( 
.A(n_157),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_250),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_159),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_156),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_183),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_224),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_230),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_277),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_232),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_233),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_162),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_159),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_235),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_187),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_195),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_157),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_237),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_239),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_290),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_240),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_181),
.B(n_196),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_226),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_162),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_207),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_194),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_241),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_159),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_242),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_196),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_253),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_164),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_326),
.A2(n_274),
.B1(n_165),
.B2(n_190),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_328),
.B(n_169),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_194),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_253),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g412 ( 
.A(n_364),
.B(n_163),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_331),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_280),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_337),
.B(n_292),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_320),
.B(n_157),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_292),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_317),
.B(n_322),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_177),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_319),
.B(n_307),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_169),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_323),
.B(n_175),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_175),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_395),
.B(n_311),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_395),
.B(n_315),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_424),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_413),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_444),
.B(n_327),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_408),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_333),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_335),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_159),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_444),
.B(n_340),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_413),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_436),
.A2(n_310),
.B1(n_375),
.B2(n_370),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_342),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_409),
.B(n_351),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_409),
.B(n_369),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_423),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_388),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_402),
.B(n_345),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_443),
.B(n_349),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_387),
.B(n_280),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_423),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_438),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_452),
.B(n_369),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_449),
.B(n_350),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_359),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_408),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g504 ( 
.A1(n_412),
.A2(n_325),
.B1(n_312),
.B2(n_319),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_441),
.A2(n_312),
.B1(n_249),
.B2(n_215),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_360),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

INVx4_ASAP7_75t_SL g510 ( 
.A(n_400),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_452),
.B(n_374),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_430),
.B(n_158),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_417),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_394),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_362),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_R g520 ( 
.A(n_417),
.B(n_308),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_407),
.B(n_166),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_SL g522 ( 
.A1(n_430),
.A2(n_227),
.B(n_225),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_363),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_438),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_437),
.B(n_366),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_374),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_401),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_437),
.B(n_371),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_387),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_403),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_430),
.B(n_372),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_404),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_429),
.B(n_381),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_429),
.A2(n_373),
.B1(n_383),
.B2(n_219),
.Y(n_540)
);

INVx4_ASAP7_75t_SL g541 ( 
.A(n_424),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_404),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_408),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_412),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g545 ( 
.A(n_407),
.B(n_166),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_410),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_417),
.B(n_246),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_410),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_415),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_437),
.B(n_189),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_419),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_419),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_387),
.A2(n_161),
.B(n_155),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_389),
.B(n_173),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_391),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_389),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_447),
.B(n_353),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_389),
.A2(n_252),
.B1(n_275),
.B2(n_288),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_SL g566 ( 
.A(n_399),
.B(n_223),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_389),
.B(n_166),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_448),
.B(n_178),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_448),
.B(n_178),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_447),
.B(n_353),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_433),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_434),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_446),
.B(n_379),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_434),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_399),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_440),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_424),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_448),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_391),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_437),
.B(n_218),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_448),
.B(n_180),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_384),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_389),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_384),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_447),
.B(n_353),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_384),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_428),
.A2(n_278),
.B1(n_294),
.B2(n_353),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_385),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_428),
.Y(n_598)
);

OAI22x1_ASAP7_75t_L g599 ( 
.A1(n_451),
.A2(n_163),
.B1(n_306),
.B2(n_305),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_451),
.B(n_379),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_466),
.B(n_166),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_477),
.B(n_332),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_480),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_498),
.B(n_447),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_243),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_R g607 ( 
.A(n_544),
.B(n_343),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_480),
.Y(n_608)
);

BUFx6f_ASAP7_75t_SL g609 ( 
.A(n_532),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_591),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_497),
.B(n_447),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_SL g613 ( 
.A(n_496),
.B(n_354),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_465),
.B(n_341),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_474),
.B(n_440),
.C(n_199),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_454),
.B(n_180),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_535),
.A2(n_361),
.B1(n_254),
.B2(n_260),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_497),
.B(n_448),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_531),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_511),
.B(n_448),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_511),
.B(n_450),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_457),
.B(n_166),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_485),
.B(n_450),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_591),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_524),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_502),
.B(n_450),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_507),
.B(n_450),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_592),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_495),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_517),
.B(n_450),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_509),
.B(n_229),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_559),
.B(n_450),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_598),
.B(n_186),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_593),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_598),
.B(n_450),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_522),
.A2(n_428),
.B(n_176),
.C(n_174),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_478),
.B(n_450),
.Y(n_639)
);

OR2x2_ASAP7_75t_SL g640 ( 
.A(n_566),
.B(n_262),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_479),
.B(n_336),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_524),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_504),
.B(n_229),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_478),
.B(n_428),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_593),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

AND2x6_ASAP7_75t_SL g648 ( 
.A(n_539),
.B(n_547),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_336),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_495),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_509),
.B(n_186),
.Y(n_651)
);

INVx8_ASAP7_75t_L g652 ( 
.A(n_547),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_509),
.B(n_186),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_582),
.B(n_186),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_524),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_553),
.B(n_428),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_523),
.B(n_186),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_527),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_463),
.A2(n_264),
.B1(n_248),
.B2(n_245),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_456),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_587),
.B(n_420),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_456),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_526),
.B(n_271),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_487),
.B(n_231),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_579),
.B(n_451),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_420),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_470),
.A2(n_272),
.B1(n_247),
.B2(n_269),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_471),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_530),
.B(n_271),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_477),
.B(n_231),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_536),
.B(n_558),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_536),
.B(n_271),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_482),
.B(n_420),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_482),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_597),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_536),
.B(n_558),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_473),
.B(n_281),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_460),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_490),
.B(n_420),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_462),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_490),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_496),
.B(n_380),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_495),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_506),
.B(n_211),
.C(n_210),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_460),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_540),
.B(n_380),
.C(n_256),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_462),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_505),
.B(n_508),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_566),
.B(n_209),
.C(n_259),
.Y(n_691)
);

AND2x6_ASAP7_75t_SL g692 ( 
.A(n_547),
.B(n_185),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_558),
.B(n_568),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_547),
.B(n_281),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_467),
.A2(n_263),
.B1(n_285),
.B2(n_271),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_514),
.B(n_286),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_505),
.B(n_286),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_512),
.B(n_461),
.C(n_581),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_491),
.B(n_271),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_495),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_516),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_491),
.B(n_293),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_516),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_579),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_568),
.B(n_586),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_467),
.A2(n_261),
.B1(n_197),
.B2(n_204),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_568),
.B(n_206),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_586),
.B(n_217),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_532),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_586),
.B(n_220),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_518),
.B(n_420),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_512),
.B(n_276),
.C(n_188),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_518),
.B(n_442),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_599),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_557),
.B(n_228),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_528),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_468),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_528),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_529),
.B(n_442),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_529),
.B(n_442),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_542),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_491),
.B(n_293),
.Y(n_724)
);

AOI221xp5_ASAP7_75t_L g725 ( 
.A1(n_599),
.A2(n_167),
.B1(n_306),
.B2(n_305),
.C(n_172),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_468),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_491),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_546),
.B(n_442),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_546),
.B(n_442),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_548),
.B(n_391),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_557),
.B(n_489),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_548),
.B(n_408),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_601),
.B(n_234),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_550),
.B(n_408),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_550),
.B(n_414),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_554),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_554),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_581),
.A2(n_284),
.B1(n_172),
.B2(n_182),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_469),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_555),
.B(n_295),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_469),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_476),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_601),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_555),
.B(n_295),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_564),
.B(n_414),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_564),
.B(n_414),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_565),
.B(n_414),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_557),
.B(n_236),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_491),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_565),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_532),
.B(n_201),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_472),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_570),
.B(n_414),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_455),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_573),
.A2(n_304),
.B1(n_302),
.B2(n_300),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_570),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_561),
.B(n_300),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_520),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_489),
.B(n_244),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_574),
.A2(n_304),
.B1(n_302),
.B2(n_301),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_577),
.B(n_418),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_577),
.B(n_238),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_476),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_580),
.B(n_418),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_455),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_493),
.B(n_251),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_588),
.A2(n_268),
.B(n_303),
.C(n_258),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_580),
.B(n_418),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_521),
.A2(n_297),
.B1(n_182),
.B2(n_279),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_572),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_472),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_584),
.B(n_431),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_493),
.B(n_431),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_612),
.A2(n_464),
.B(n_543),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_700),
.B(n_749),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_627),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_618),
.B(n_534),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_614),
.B(n_584),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_619),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_673),
.A2(n_503),
.B(n_513),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_614),
.B(n_743),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_743),
.B(n_589),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_673),
.A2(n_693),
.B(n_678),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_616),
.B(n_589),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_616),
.B(n_499),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_641),
.B(n_167),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_678),
.A2(n_571),
.B(n_513),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_605),
.B(n_499),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_661),
.B(n_500),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_663),
.B(n_500),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_758),
.B(n_682),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_629),
.Y(n_792)
);

OAI321xp33_ASAP7_75t_L g793 ( 
.A1(n_679),
.A2(n_596),
.A3(n_563),
.B1(n_556),
.B2(n_519),
.C(n_525),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_705),
.A2(n_575),
.B1(n_594),
.B2(n_501),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_649),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_689),
.B(n_633),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_705),
.A2(n_521),
.B1(n_545),
.B2(n_515),
.Y(n_797)
);

AOI21x1_ASAP7_75t_L g798 ( 
.A1(n_674),
.A2(n_556),
.B(n_501),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_603),
.B(n_534),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_693),
.A2(n_513),
.B(n_590),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_670),
.B(n_515),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_680),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_684),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_714),
.A2(n_545),
.B1(n_562),
.B2(n_560),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_706),
.A2(n_459),
.B(n_590),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_687),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_714),
.A2(n_537),
.B1(n_525),
.B2(n_533),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_676),
.B(n_519),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_643),
.A2(n_537),
.B(n_578),
.C(n_576),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_706),
.A2(n_458),
.B(n_590),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_683),
.B(n_533),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_642),
.B(n_534),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_620),
.A2(n_453),
.B(n_492),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_621),
.A2(n_571),
.B(n_459),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_623),
.A2(n_571),
.B(n_459),
.Y(n_815)
);

AO21x1_ASAP7_75t_L g816 ( 
.A1(n_602),
.A2(n_551),
.B(n_538),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_701),
.B(n_538),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_626),
.A2(n_583),
.B(n_458),
.Y(n_818)
);

BUFx12f_ASAP7_75t_L g819 ( 
.A(n_771),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_628),
.A2(n_583),
.B(n_458),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_702),
.B(n_704),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_619),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_679),
.A2(n_551),
.B(n_578),
.C(n_576),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_631),
.A2(n_657),
.B(n_662),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_731),
.A2(n_639),
.B(n_644),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_602),
.A2(n_560),
.B1(n_549),
.B2(n_552),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_731),
.A2(n_583),
.B(n_455),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_666),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_634),
.A2(n_455),
.B(n_585),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_718),
.B(n_549),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_720),
.B(n_552),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_700),
.B(n_562),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_700),
.B(n_567),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_666),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_723),
.B(n_567),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_645),
.B(n_510),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_700),
.B(n_455),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_637),
.A2(n_600),
.B(n_585),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_607),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_736),
.B(n_453),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_632),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_737),
.B(n_453),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_633),
.B(n_492),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_665),
.A2(n_299),
.B(n_298),
.C(n_297),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_716),
.B(n_492),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_630),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_651),
.A2(n_488),
.B(n_486),
.C(n_421),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_672),
.B(n_279),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_699),
.A2(n_600),
.B(n_585),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_607),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_750),
.B(n_486),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_756),
.B(n_488),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_674),
.A2(n_569),
.B(n_421),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_770),
.A2(n_600),
.B(n_585),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_659),
.B(n_572),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_770),
.A2(n_600),
.B(n_585),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_730),
.A2(n_600),
.B(n_572),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_690),
.B(n_572),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_672),
.B(n_572),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_697),
.B(n_569),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_754),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_630),
.Y(n_862)
);

O2A1O1Ixp5_ASAP7_75t_L g863 ( 
.A1(n_651),
.A2(n_653),
.B(n_671),
.C(n_658),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_754),
.B(n_765),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_754),
.B(n_765),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_708),
.A2(n_711),
.B(n_709),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_604),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_SL g868 ( 
.A(n_609),
.B(n_283),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_695),
.B(n_431),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_727),
.A2(n_665),
.B1(n_695),
.B2(n_608),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_696),
.B(n_265),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_708),
.A2(n_475),
.B(n_481),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_709),
.A2(n_475),
.B(n_481),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_751),
.B(n_284),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_710),
.B(n_283),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_754),
.B(n_510),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_711),
.A2(n_475),
.B(n_481),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_765),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_697),
.B(n_569),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_765),
.B(n_510),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_719),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_749),
.A2(n_475),
.B(n_481),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_752),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_740),
.B(n_569),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_652),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_749),
.A2(n_475),
.B(n_481),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_615),
.B(n_98),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_611),
.A2(n_569),
.B1(n_421),
.B2(n_431),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_650),
.A2(n_483),
.B(n_484),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_726),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_650),
.A2(n_483),
.B(n_484),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_625),
.B(n_298),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_609),
.B(n_299),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_617),
.B(n_266),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_715),
.A2(n_722),
.B(n_721),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_727),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_685),
.A2(n_483),
.B(n_484),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_655),
.B(n_270),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_685),
.A2(n_483),
.B(n_484),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_728),
.A2(n_569),
.B(n_411),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_761),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_613),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_606),
.A2(n_483),
.B(n_484),
.Y(n_903)
);

NOR2x1p5_ASAP7_75t_L g904 ( 
.A(n_713),
.B(n_273),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_740),
.B(n_510),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_653),
.B(n_411),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_739),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_667),
.A2(n_411),
.B(n_406),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_654),
.A2(n_406),
.B(n_405),
.C(n_396),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_660),
.B(n_151),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_729),
.A2(n_406),
.B(n_405),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_744),
.B(n_541),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_744),
.B(n_541),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_762),
.B(n_541),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_762),
.B(n_541),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_764),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_733),
.B(n_431),
.Y(n_918)
);

AOI33xp33_ASAP7_75t_L g919 ( 
.A1(n_738),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_14),
.B3(n_15),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_768),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_733),
.B(n_431),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_675),
.B(n_431),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_694),
.B(n_738),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_681),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_654),
.B(n_712),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_742),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_763),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_757),
.B(n_405),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_652),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_769),
.A2(n_396),
.B(n_385),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_732),
.A2(n_396),
.B(n_385),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_610),
.B(n_18),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_734),
.A2(n_148),
.B(n_146),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_652),
.Y(n_934)
);

OAI22xp33_ASAP7_75t_L g935 ( 
.A1(n_725),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_624),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_694),
.B(n_23),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_636),
.B(n_23),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_646),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_658),
.A2(n_137),
.B(n_131),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_735),
.A2(n_126),
.B(n_125),
.Y(n_941)
);

OAI21xp33_ASAP7_75t_L g942 ( 
.A1(n_769),
.A2(n_686),
.B(n_688),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_745),
.A2(n_112),
.B(n_108),
.Y(n_943)
);

AND2x6_ASAP7_75t_L g944 ( 
.A(n_647),
.B(n_103),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_656),
.B(n_25),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_772),
.B(n_102),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_669),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_677),
.B(n_25),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_664),
.A2(n_83),
.B(n_79),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_746),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_638),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_622),
.B(n_33),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_668),
.B(n_67),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_747),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_622),
.A2(n_66),
.B1(n_63),
.B2(n_37),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_753),
.A2(n_34),
.B(n_36),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_698),
.B(n_37),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_759),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_755),
.B(n_640),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_664),
.A2(n_38),
.B(n_43),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_671),
.A2(n_38),
.B(n_43),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_691),
.B(n_49),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_703),
.A2(n_44),
.B(n_45),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_796),
.B(n_648),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_803),
.B(n_760),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_824),
.A2(n_724),
.B(n_748),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_836),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_792),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_796),
.B(n_767),
.Y(n_969)
);

CKINVDCx10_ASAP7_75t_R g970 ( 
.A(n_839),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_836),
.Y(n_971)
);

NOR2x1_ASAP7_75t_R g972 ( 
.A(n_819),
.B(n_692),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_846),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_866),
.A2(n_717),
.B(n_748),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_SL g975 ( 
.A1(n_777),
.A2(n_946),
.B(n_766),
.C(n_759),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_776),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_846),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_923),
.A2(n_707),
.B(n_717),
.C(n_635),
.Y(n_978)
);

CKINVDCx14_ASAP7_75t_R g979 ( 
.A(n_850),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_SL g980 ( 
.A(n_935),
.B(n_766),
.C(n_635),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_869),
.A2(n_707),
.B1(n_773),
.B2(n_49),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_778),
.B(n_773),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_781),
.B(n_46),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_SL g984 ( 
.A1(n_923),
.A2(n_48),
.B1(n_937),
.B2(n_869),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_942),
.A2(n_48),
.B1(n_937),
.B2(n_894),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_791),
.B(n_795),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_825),
.A2(n_858),
.B(n_818),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_791),
.B(n_803),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_799),
.B(n_784),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_902),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_802),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_815),
.A2(n_820),
.B(n_788),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_870),
.A2(n_785),
.B1(n_896),
.B2(n_859),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_894),
.B(n_848),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_845),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_814),
.A2(n_783),
.B(n_813),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_901),
.B(n_917),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_959),
.A2(n_777),
.B1(n_834),
.B2(n_828),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_878),
.Y(n_999)
);

AOI22x1_ASAP7_75t_L g1000 ( 
.A1(n_920),
.A2(n_954),
.B1(n_950),
.B2(n_924),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_821),
.B(n_841),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_896),
.A2(n_843),
.B1(n_860),
.B2(n_884),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_874),
.B(n_875),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_774),
.A2(n_800),
.B(n_787),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_806),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_828),
.B(n_959),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_871),
.B(n_935),
.C(n_962),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_883),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_SL g1010 ( 
.A1(n_871),
.A2(n_957),
.B1(n_893),
.B2(n_868),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_805),
.A2(n_810),
.B(n_775),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_827),
.A2(n_780),
.B(n_905),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_892),
.A2(n_898),
.B1(n_963),
.B2(n_929),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_952),
.A2(n_944),
.B1(n_940),
.B2(n_949),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_837),
.A2(n_916),
.B(n_915),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_846),
.B(n_862),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_851),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_845),
.B(n_867),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_837),
.A2(n_895),
.B(n_925),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_806),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_786),
.A2(n_904),
.B1(n_934),
.B2(n_958),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_862),
.B(n_779),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_878),
.Y(n_1023)
);

CKINVDCx10_ASAP7_75t_R g1024 ( 
.A(n_812),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_843),
.B(n_782),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_863),
.A2(n_823),
.B(n_879),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_844),
.B(n_779),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_822),
.B(n_789),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_822),
.A2(n_912),
.B1(n_914),
.B2(n_794),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_918),
.A2(n_921),
.B(n_829),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_857),
.A2(n_838),
.B(n_903),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_862),
.B(n_878),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_885),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_910),
.A2(n_953),
.B1(n_881),
.B2(n_907),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_854),
.A2(n_856),
.B(n_833),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_823),
.A2(n_844),
.B(n_951),
.C(n_835),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_862),
.B(n_878),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_934),
.B(n_790),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_832),
.A2(n_833),
.B(n_864),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_809),
.A2(n_793),
.B(n_831),
.C(n_801),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_852),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_SL g1042 ( 
.A(n_885),
.B(n_887),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_832),
.A2(n_865),
.B(n_864),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_808),
.A2(n_830),
.B1(n_817),
.B2(n_811),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_927),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_926),
.B(n_927),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_797),
.A2(n_804),
.B1(n_855),
.B2(n_826),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_947),
.B(n_913),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_951),
.A2(n_938),
.B(n_945),
.C(n_948),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_890),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_890),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_947),
.B(n_936),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_939),
.B(n_861),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_865),
.A2(n_849),
.B(n_886),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_936),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_861),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_960),
.A2(n_961),
.B(n_855),
.C(n_930),
.Y(n_1057)
);

NOR2x1_ASAP7_75t_L g1058 ( 
.A(n_932),
.B(n_946),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_956),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_840),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_842),
.B(n_826),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_807),
.B(n_928),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_876),
.B(n_880),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_876),
.B(n_880),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_900),
.A2(n_847),
.B(n_922),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_798),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_922),
.B(n_816),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_944),
.A2(n_955),
.B1(n_906),
.B2(n_943),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_933),
.B(n_941),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_944),
.B(n_853),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_944),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_909),
.A2(n_911),
.B(n_908),
.C(n_931),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_919),
.B(n_944),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_919),
.A2(n_888),
.B(n_873),
.C(n_877),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_882),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_872),
.A2(n_889),
.B(n_891),
.C(n_897),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_899),
.A2(n_869),
.B1(n_784),
.B2(n_870),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_824),
.A2(n_678),
.B(n_673),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_869),
.A2(n_784),
.B1(n_870),
.B2(n_923),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_828),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_923),
.A2(n_942),
.B(n_937),
.C(n_466),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_846),
.B(n_630),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_836),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_778),
.A2(n_781),
.B(n_937),
.C(n_784),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_803),
.B(n_603),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_796),
.B(n_544),
.Y(n_1086)
);

BUFx2_ASAP7_75t_SL g1087 ( 
.A(n_934),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_863),
.A2(n_825),
.B(n_783),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_869),
.A2(n_923),
.B1(n_937),
.B2(n_942),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_796),
.B(n_544),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_923),
.A2(n_869),
.B1(n_942),
.B2(n_937),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_923),
.A2(n_942),
.B(n_937),
.C(n_466),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_846),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_878),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_792),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_792),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_824),
.A2(n_678),
.B(n_673),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_869),
.A2(n_923),
.B1(n_937),
.B2(n_942),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_824),
.A2(n_678),
.B(n_673),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_796),
.B(n_544),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_836),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_792),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_824),
.A2(n_678),
.B(n_673),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_923),
.A2(n_942),
.B(n_937),
.C(n_466),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_878),
.Y(n_1105)
);

CKINVDCx11_ASAP7_75t_R g1106 ( 
.A(n_819),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_803),
.B(n_603),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1005),
.A2(n_966),
.B(n_996),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1081),
.A2(n_1104),
.B(n_1092),
.C(n_994),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_SL g1110 ( 
.A1(n_969),
.A2(n_1079),
.B(n_1100),
.C(n_1090),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_997),
.B(n_1086),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1077),
.A2(n_1029),
.A3(n_1047),
.B(n_993),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1091),
.A2(n_1008),
.B(n_1098),
.C(n_1089),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1009),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1011),
.A2(n_987),
.B(n_992),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_976),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_990),
.A2(n_1002),
.B1(n_998),
.B2(n_964),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_1084),
.A2(n_1008),
.B(n_1049),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1017),
.B(n_1041),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1089),
.A2(n_1098),
.B(n_1084),
.C(n_985),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_1033),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_984),
.A2(n_1010),
.B1(n_1007),
.B2(n_1085),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_989),
.A2(n_983),
.B(n_995),
.C(n_978),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1078),
.A2(n_1099),
.B(n_1103),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1067),
.A2(n_1003),
.A3(n_1015),
.B(n_1012),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_973),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1107),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1004),
.B(n_1080),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_968),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1095),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1097),
.A2(n_1088),
.B(n_1019),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_974),
.A2(n_1025),
.B(n_1031),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1054),
.A2(n_1030),
.B(n_1035),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1062),
.A2(n_1026),
.B(n_1040),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1057),
.A2(n_1074),
.A3(n_1066),
.B(n_981),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_1106),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1069),
.A2(n_1049),
.B(n_1058),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_975),
.A2(n_1036),
.B(n_1065),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_995),
.B(n_988),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_965),
.B(n_1018),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_982),
.B(n_1060),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_980),
.A2(n_1010),
.B(n_1027),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1080),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_973),
.B(n_972),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1039),
.A2(n_1014),
.B(n_1043),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_1001),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_1102),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1013),
.B(n_967),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1069),
.A2(n_1014),
.B(n_1076),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1096),
.B(n_1048),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1076),
.A2(n_1072),
.B(n_1000),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_1068),
.A2(n_1061),
.B(n_1073),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1028),
.B(n_967),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1063),
.A2(n_1064),
.A3(n_1050),
.B(n_1051),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1072),
.A2(n_1036),
.B(n_1068),
.Y(n_1156)
);

BUFx10_ASAP7_75t_L g1157 ( 
.A(n_1056),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_991),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1006),
.Y(n_1159)
);

NOR4xp25_ASAP7_75t_L g1160 ( 
.A(n_1059),
.B(n_1034),
.C(n_1071),
.D(n_1052),
.Y(n_1160)
);

AO32x2_ASAP7_75t_L g1161 ( 
.A1(n_977),
.A2(n_1001),
.A3(n_1093),
.B1(n_1071),
.B2(n_1069),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_SL g1162 ( 
.A(n_1087),
.B(n_1093),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1070),
.A2(n_1055),
.B(n_1020),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1070),
.A2(n_1042),
.B(n_1046),
.C(n_1045),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1053),
.A2(n_1022),
.B(n_1032),
.Y(n_1165)
);

AND3x2_ASAP7_75t_L g1166 ( 
.A(n_1023),
.B(n_1024),
.C(n_970),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_971),
.A2(n_1101),
.B(n_1083),
.C(n_1075),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1021),
.A2(n_1075),
.A3(n_1023),
.B(n_1037),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1075),
.A2(n_1016),
.B(n_1082),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_999),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_SL g1171 ( 
.A1(n_971),
.A2(n_1101),
.B(n_1083),
.C(n_1105),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_979),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1056),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1056),
.B(n_999),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_999),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1094),
.B(n_1105),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1094),
.A2(n_1081),
.B(n_1104),
.C(n_1092),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1094),
.A2(n_1008),
.B1(n_984),
.B2(n_923),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1094),
.A2(n_1089),
.B1(n_1098),
.B2(n_1091),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1105),
.B(n_461),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1026),
.A2(n_1088),
.B(n_1015),
.Y(n_1181)
);

AO21x2_ASAP7_75t_L g1182 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_1088),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_1081),
.A2(n_1104),
.B(n_1092),
.C(n_994),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_994),
.B(n_997),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_997),
.B(n_1081),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.Y(n_1186)
);

BUFx4_ASAP7_75t_SL g1187 ( 
.A(n_1033),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1008),
.A2(n_984),
.B1(n_923),
.B2(n_994),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1009),
.Y(n_1189)
);

NAND3x1_ASAP7_75t_L g1190 ( 
.A(n_1008),
.B(n_923),
.C(n_994),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1056),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_990),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1077),
.A2(n_1079),
.A3(n_1092),
.B(n_1081),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1077),
.A2(n_1079),
.A3(n_1092),
.B(n_1081),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1089),
.A2(n_1098),
.B1(n_1091),
.B2(n_1092),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.C(n_994),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_994),
.A2(n_544),
.B1(n_444),
.B2(n_696),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1085),
.B(n_1107),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1026),
.A2(n_1088),
.B(n_1015),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1077),
.A2(n_1079),
.A3(n_1092),
.B(n_1081),
.Y(n_1203)
);

AOI31xp67_ASAP7_75t_L g1204 ( 
.A1(n_1062),
.A2(n_602),
.A3(n_794),
.B(n_664),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_1088),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1011),
.A2(n_1054),
.B(n_1030),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.C(n_978),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.C(n_978),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_994),
.B(n_1008),
.C(n_1081),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1033),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_997),
.B(n_1081),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1033),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_986),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1085),
.B(n_1107),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_968),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1026),
.A2(n_1088),
.B(n_1015),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_997),
.B(n_1081),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_994),
.B(n_997),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1106),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1077),
.A2(n_1079),
.A3(n_1092),
.B(n_1081),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1009),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_1088),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1026),
.A2(n_1088),
.B(n_1015),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1077),
.A2(n_1079),
.A3(n_1092),
.B(n_1081),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1104),
.C(n_994),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1085),
.B(n_461),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_SL g1229 ( 
.A(n_984),
.B(n_869),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_L g1230 ( 
.A1(n_994),
.A2(n_923),
.B1(n_1008),
.B2(n_985),
.C(n_1104),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_968),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_973),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1005),
.A2(n_966),
.B(n_824),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1011),
.A2(n_1054),
.B(n_1030),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1230),
.A2(n_1209),
.B1(n_1188),
.B2(n_1142),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1188),
.A2(n_1142),
.B1(n_1197),
.B2(n_1229),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1136),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1229),
.A2(n_1178),
.B1(n_1218),
.B2(n_1184),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1190),
.A2(n_1140),
.B1(n_1117),
.B2(n_1200),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1114),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1189),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1219),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1111),
.A2(n_1122),
.B1(n_1144),
.B2(n_1178),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1157),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1172),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1195),
.A2(n_1196),
.B(n_1235),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1197),
.A2(n_1199),
.B1(n_1186),
.B2(n_1118),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1186),
.A2(n_1199),
.B1(n_1179),
.B2(n_1134),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1179),
.A2(n_1139),
.B1(n_1119),
.B2(n_1185),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1192),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1156),
.A2(n_1182),
.B1(n_1224),
.B2(n_1205),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1213),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1119),
.A2(n_1217),
.B1(n_1185),
.B2(n_1211),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1223),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1121),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1157),
.Y(n_1258)
);

INVx6_ASAP7_75t_L g1259 ( 
.A(n_1126),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1126),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1211),
.A2(n_1217),
.B1(n_1127),
.B2(n_1214),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_SL g1262 ( 
.A(n_1212),
.Y(n_1262)
);

INVx8_ASAP7_75t_L g1263 ( 
.A(n_1173),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1201),
.B(n_1141),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1130),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1143),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1210),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1109),
.A2(n_1198),
.B(n_1227),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1182),
.A2(n_1205),
.B1(n_1224),
.B2(n_1150),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1120),
.A2(n_1113),
.B1(n_1148),
.B2(n_1228),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1128),
.A2(n_1151),
.B1(n_1145),
.B2(n_1154),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1138),
.A2(n_1153),
.B1(n_1149),
.B2(n_1137),
.Y(n_1272)
);

INVx8_ASAP7_75t_L g1273 ( 
.A(n_1191),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1180),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1233),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_1187),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1164),
.A2(n_1177),
.B1(n_1167),
.B2(n_1123),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1145),
.A2(n_1138),
.B1(n_1153),
.B2(n_1215),
.Y(n_1278)
);

CKINVDCx8_ASAP7_75t_R g1279 ( 
.A(n_1166),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1213),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1232),
.A2(n_1158),
.B1(n_1159),
.B2(n_1183),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1174),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1175),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1162),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1155),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1181),
.A2(n_1225),
.B1(n_1216),
.B2(n_1202),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1181),
.A2(n_1202),
.B1(n_1216),
.B2(n_1225),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1176),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1168),
.Y(n_1289)
);

BUFx2_ASAP7_75t_SL g1290 ( 
.A(n_1170),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1163),
.A2(n_1165),
.B1(n_1169),
.B2(n_1147),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1163),
.A2(n_1165),
.B1(n_1146),
.B2(n_1131),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1110),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1161),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1207),
.A2(n_1208),
.B1(n_1146),
.B2(n_1152),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1160),
.B(n_1194),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1171),
.Y(n_1298)
);

INVx8_ASAP7_75t_L g1299 ( 
.A(n_1160),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1135),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1193),
.A2(n_1226),
.B1(n_1222),
.B2(n_1203),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1132),
.Y(n_1302)
);

BUFx8_ASAP7_75t_SL g1303 ( 
.A(n_1204),
.Y(n_1303)
);

OAI21xp33_ASAP7_75t_L g1304 ( 
.A1(n_1108),
.A2(n_1234),
.B(n_1231),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1193),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1124),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1193),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1125),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1133),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1220),
.A2(n_1221),
.B1(n_1226),
.B2(n_1194),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1206),
.B(n_1236),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1125),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1194),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1115),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1203),
.A2(n_1222),
.B1(n_1226),
.B2(n_1112),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1203),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1222),
.A2(n_1229),
.B1(n_1188),
.B2(n_937),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1112),
.A2(n_1008),
.B1(n_1230),
.B2(n_984),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1112),
.A2(n_1008),
.B1(n_1230),
.B2(n_984),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1114),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1114),
.Y(n_1321)
);

BUFx2_ASAP7_75t_R g1322 ( 
.A(n_1172),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1201),
.B(n_1214),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1229),
.A2(n_984),
.B1(n_869),
.B2(n_923),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1114),
.Y(n_1325)
);

INVx6_ASAP7_75t_L g1326 ( 
.A(n_1126),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1188),
.A2(n_994),
.B1(n_1092),
.B2(n_1081),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1230),
.A2(n_1008),
.B1(n_984),
.B2(n_1209),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1230),
.A2(n_1008),
.B1(n_984),
.B2(n_1209),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1129),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1126),
.B(n_1233),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1201),
.B(n_1214),
.Y(n_1332)
);

OAI22x1_ASAP7_75t_L g1333 ( 
.A1(n_1188),
.A2(n_1178),
.B1(n_923),
.B2(n_994),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1229),
.A2(n_1188),
.B1(n_1178),
.B2(n_923),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_L g1335 ( 
.A(n_1136),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1136),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1116),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1136),
.Y(n_1338)
);

CKINVDCx6p67_ASAP7_75t_R g1339 ( 
.A(n_1136),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1285),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1300),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1238),
.B(n_1305),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1265),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1239),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1307),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1313),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1266),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1316),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1294),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1248),
.A2(n_1311),
.B(n_1310),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1297),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1306),
.B(n_1289),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1288),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1328),
.A2(n_1329),
.B1(n_1324),
.B2(n_1334),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1266),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1309),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1301),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1308),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1308),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1311),
.A2(n_1310),
.B(n_1287),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1282),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1312),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1312),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1274),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1327),
.A2(n_1268),
.B(n_1329),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1314),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1296),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1287),
.A2(n_1292),
.B(n_1304),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1328),
.B(n_1237),
.C(n_1241),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1278),
.A2(n_1255),
.B(n_1251),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1323),
.B(n_1332),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1280),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1272),
.A2(n_1249),
.B(n_1269),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1269),
.A2(n_1291),
.B(n_1315),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1337),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1238),
.B(n_1305),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1284),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1255),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1315),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1333),
.A2(n_1245),
.B(n_1270),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1237),
.B(n_1249),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1302),
.A2(n_1250),
.B(n_1240),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1299),
.B(n_1275),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1253),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_1257),
.Y(n_1388)
);

INVx6_ASAP7_75t_L g1389 ( 
.A(n_1259),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1324),
.A2(n_1334),
.B1(n_1240),
.B2(n_1299),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1250),
.B(n_1272),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_SL g1393 ( 
.A(n_1279),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1281),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1264),
.B(n_1261),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1303),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1251),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1286),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1278),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1261),
.B(n_1325),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1295),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1295),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1256),
.B(n_1320),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1298),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1280),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1317),
.A2(n_1293),
.B(n_1330),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1271),
.A2(n_1331),
.B(n_1284),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1271),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1284),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1293),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1284),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1276),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1242),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1242),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1243),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1290),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1383),
.B(n_1243),
.Y(n_1417)
);

OAI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1365),
.A2(n_1254),
.B(n_1321),
.C(n_1239),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1383),
.B(n_1321),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1280),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1409),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1344),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1407),
.A2(n_1267),
.B(n_1263),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1369),
.A2(n_1263),
.B(n_1335),
.C(n_1273),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1350),
.A2(n_1283),
.B(n_1246),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1354),
.A2(n_1262),
.B1(n_1326),
.B2(n_1260),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1391),
.A2(n_1260),
.B1(n_1326),
.B2(n_1259),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1384),
.A2(n_1258),
.B(n_1246),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1382),
.A2(n_1335),
.B(n_1258),
.C(n_1259),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1398),
.B(n_1380),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1392),
.B(n_1339),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1340),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1358),
.B(n_1252),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1368),
.A2(n_1322),
.B(n_1247),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1358),
.B(n_1338),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1359),
.B(n_1336),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1392),
.B(n_1244),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1381),
.A2(n_1382),
.B(n_1372),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1344),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1368),
.A2(n_1375),
.B(n_1350),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1351),
.B(n_1349),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1370),
.A2(n_1366),
.B(n_1372),
.Y(n_1442)
);

AO32x2_ASAP7_75t_L g1443 ( 
.A1(n_1353),
.A2(n_1378),
.A3(n_1367),
.B1(n_1373),
.B2(n_1410),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_SL g1444 ( 
.A(n_1342),
.B(n_1377),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1375),
.A2(n_1360),
.B(n_1399),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1361),
.B(n_1395),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1396),
.A2(n_1372),
.B1(n_1390),
.B2(n_1385),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1385),
.A2(n_1390),
.B(n_1342),
.C(n_1377),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1376),
.B(n_1374),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1347),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1381),
.A2(n_1357),
.B(n_1400),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1355),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1372),
.A2(n_1397),
.B(n_1408),
.C(n_1410),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1360),
.A2(n_1404),
.B(n_1370),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1374),
.B(n_1343),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1372),
.B(n_1386),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1408),
.A2(n_1397),
.B(n_1366),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1379),
.A2(n_1357),
.B1(n_1371),
.B2(n_1401),
.C(n_1402),
.Y(n_1459)
);

AND2x2_ASAP7_75t_SL g1460 ( 
.A(n_1374),
.B(n_1352),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1374),
.B(n_1343),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1403),
.B(n_1388),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1396),
.A2(n_1352),
.B(n_1379),
.C(n_1394),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1459),
.A2(n_1370),
.B1(n_1402),
.B2(n_1401),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1455),
.B(n_1348),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1443),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_L g1468 ( 
.A(n_1425),
.B(n_1411),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1346),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1448),
.B(n_1406),
.C(n_1416),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1346),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1455),
.B(n_1461),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1460),
.B(n_1348),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1450),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1432),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1346),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1456),
.B(n_1356),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1460),
.B(n_1345),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1451),
.A2(n_1437),
.B1(n_1431),
.B2(n_1446),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1445),
.B(n_1345),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1430),
.B(n_1458),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1445),
.B(n_1341),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1406),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1431),
.B(n_1413),
.Y(n_1484)
);

AOI33xp33_ASAP7_75t_L g1485 ( 
.A1(n_1465),
.A2(n_1437),
.A3(n_1417),
.B1(n_1419),
.B2(n_1453),
.B3(n_1420),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1472),
.B(n_1454),
.Y(n_1486)
);

AND2x2_ASAP7_75t_SL g1487 ( 
.A(n_1467),
.B(n_1352),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1482),
.Y(n_1488)
);

OAI31xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1470),
.A2(n_1447),
.A3(n_1438),
.B(n_1418),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1482),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1465),
.A2(n_1451),
.B1(n_1444),
.B2(n_1442),
.C(n_1457),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1475),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1475),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1480),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1477),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1469),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1479),
.A2(n_1388),
.B1(n_1439),
.B2(n_1422),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1477),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1479),
.A2(n_1464),
.B1(n_1424),
.B2(n_1428),
.C(n_1429),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1456),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1469),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1476),
.B(n_1443),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1463),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1466),
.B(n_1441),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1492),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1501),
.B(n_1471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1492),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1492),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1496),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1421),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1487),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1500),
.B(n_1483),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1496),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1490),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1483),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1487),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1496),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1508),
.B(n_1476),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1495),
.B(n_1422),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1478),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1508),
.B(n_1478),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1498),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1503),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1503),
.B(n_1506),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1494),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1490),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1495),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1520),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1520),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1519),
.B(n_1506),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1519),
.B(n_1506),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1534),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1540),
.A2(n_1505),
.B(n_1491),
.C(n_1470),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1487),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1536),
.B(n_1511),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1536),
.B(n_1506),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1534),
.Y(n_1550)
);

NOR2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1527),
.B(n_1439),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1540),
.B(n_1485),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1504),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1502),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1531),
.B(n_1485),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1538),
.A2(n_1489),
.B(n_1491),
.Y(n_1557)
);

NOR2x1p5_ASAP7_75t_SL g1558 ( 
.A(n_1534),
.B(n_1488),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1513),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1489),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1515),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1516),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1516),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1514),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1530),
.B(n_1512),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1517),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1536),
.B(n_1511),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1517),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1523),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1523),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1535),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1529),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1578)
);

AOI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1518),
.A2(n_1505),
.B(n_1423),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1518),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1518),
.A2(n_1406),
.B1(n_1434),
.B2(n_1352),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1529),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1555),
.B(n_1575),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1556),
.B(n_1412),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1575),
.A2(n_1433),
.B1(n_1436),
.B2(n_1462),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1552),
.B(n_1557),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1532),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1541),
.B(n_1538),
.Y(n_1589)
);

NAND4xp25_ASAP7_75t_L g1590 ( 
.A(n_1562),
.B(n_1420),
.C(n_1426),
.D(n_1419),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1551),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1542),
.B(n_1532),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1555),
.B(n_1536),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1554),
.B(n_1533),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1577),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1533),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1577),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1555),
.B(n_1533),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1582),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1572),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1545),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1578),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_1514),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1548),
.B(n_1499),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1514),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1572),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1559),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1535),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1560),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1499),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1576),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1567),
.B(n_1509),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1561),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1547),
.B(n_1509),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1549),
.B(n_1499),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1549),
.B(n_1535),
.Y(n_1617)
);

AOI222xp33_ASAP7_75t_L g1618 ( 
.A1(n_1587),
.A2(n_1558),
.B1(n_1581),
.B2(n_1580),
.C1(n_1493),
.C2(n_1497),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1588),
.A2(n_1579),
.B1(n_1581),
.B2(n_1535),
.C(n_1550),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1598),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1596),
.B(n_1545),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1613),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1583),
.A2(n_1591),
.B(n_1584),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1543),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1595),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1595),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1585),
.A2(n_1544),
.B1(n_1543),
.B2(n_1549),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1593),
.B(n_1544),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1611),
.Y(n_1632)
);

OAI21xp33_ASAP7_75t_L g1633 ( 
.A1(n_1592),
.A2(n_1550),
.B(n_1484),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1609),
.B(n_1486),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1614),
.B(n_1486),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1597),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1593),
.A2(n_1433),
.B(n_1436),
.C(n_1393),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1602),
.A2(n_1589),
.B1(n_1600),
.B2(n_1606),
.C(n_1586),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1608),
.A2(n_1576),
.B1(n_1503),
.B2(n_1506),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1600),
.B(n_1606),
.C(n_1602),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1620),
.A2(n_1589),
.B1(n_1586),
.B2(n_1594),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1639),
.B(n_1618),
.C(n_1619),
.Y(n_1644)
);

AND2x4_ASAP7_75t_SL g1645 ( 
.A(n_1623),
.B(n_1433),
.Y(n_1645)
);

OAI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1621),
.A2(n_1616),
.B(n_1612),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1642),
.A2(n_1607),
.B1(n_1601),
.B2(n_1608),
.C(n_1605),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1624),
.A2(n_1608),
.B(n_1601),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1637),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1632),
.B(n_1607),
.Y(n_1650)
);

OAI211xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1630),
.A2(n_1605),
.B(n_1603),
.C(n_1615),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

INVxp33_ASAP7_75t_L g1653 ( 
.A(n_1630),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1629),
.B(n_1616),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1638),
.A2(n_1603),
.B1(n_1617),
.B2(n_1535),
.C(n_1610),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1622),
.B(n_1604),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1638),
.B(n_1576),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1627),
.B(n_1604),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1631),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1631),
.A2(n_1434),
.B1(n_1436),
.B2(n_1406),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_1625),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1653),
.B(n_1636),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1660),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1645),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1644),
.A2(n_1633),
.B1(n_1641),
.B2(n_1640),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1654),
.B(n_1610),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1647),
.B(n_1634),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1643),
.A2(n_1635),
.B(n_1617),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1657),
.B(n_1521),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1651),
.A2(n_1435),
.B(n_1506),
.Y(n_1671)
);

OAI321xp33_ASAP7_75t_L g1672 ( 
.A1(n_1655),
.A2(n_1427),
.A3(n_1386),
.B1(n_1570),
.B2(n_1566),
.C(n_1574),
.Y(n_1672)
);

OAI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1663),
.A2(n_1650),
.B(n_1648),
.C(n_1659),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1664),
.B(n_1659),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1662),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1666),
.B(n_1658),
.C(n_1646),
.D(n_1652),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1664),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1667),
.B(n_1656),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1665),
.B(n_1521),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1670),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1669),
.Y(n_1681)
);

AOI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1673),
.A2(n_1668),
.B(n_1671),
.C(n_1672),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1681),
.A2(n_1661),
.B1(n_1573),
.B2(n_1565),
.C(n_1563),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1680),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1673),
.A2(n_1661),
.B1(n_1497),
.B2(n_1493),
.C(n_1537),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1676),
.A2(n_1497),
.B1(n_1493),
.B2(n_1537),
.C(n_1521),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1684),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1683),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1682),
.A2(n_1678),
.B1(n_1674),
.B2(n_1675),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1686),
.A2(n_1677),
.B(n_1679),
.C(n_1373),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1685),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1684),
.Y(n_1692)
);

NAND4xp75_ASAP7_75t_L g1693 ( 
.A(n_1687),
.B(n_1468),
.C(n_1434),
.D(n_1525),
.Y(n_1693)
);

XNOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1691),
.B(n_1435),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1692),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1692),
.B(n_1435),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_L g1697 ( 
.A(n_1688),
.B(n_1689),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1690),
.B(n_1405),
.C(n_1484),
.Y(n_1698)
);

NOR2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1695),
.B(n_1405),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1694),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1699),
.Y(n_1701)
);

OA22x2_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1700),
.B1(n_1698),
.B2(n_1696),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1702),
.B(n_1693),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1702),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1704),
.A2(n_1703),
.B1(n_1405),
.B2(n_1389),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1703),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1537),
.B1(n_1524),
.B2(n_1539),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1705),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1708),
.B(n_1537),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1709),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1710),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_R g1712 ( 
.A1(n_1711),
.A2(n_1707),
.B1(n_1528),
.B2(n_1539),
.C(n_1522),
.Y(n_1712)
);

AOI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1414),
.B(n_1415),
.C(n_1409),
.Y(n_1713)
);


endmodule