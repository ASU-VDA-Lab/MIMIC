module fake_ibex_434_n_1526 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_274, n_55, n_130, n_275, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1526);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_274;
input n_55;
input n_130;
input n_275;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1526;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1421;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g281 ( 
.A(n_39),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_44),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_85),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_224),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_174),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_259),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_239),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_200),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_220),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_1),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_76),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_171),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_107),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_63),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_232),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_147),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_133),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_37),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_129),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_152),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_93),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_210),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_16),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_36),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_129),
.B(n_21),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_103),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_144),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_29),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_45),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_214),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_66),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_219),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_172),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_176),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_158),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_6),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_183),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_43),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_95),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_53),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_257),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_225),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_108),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_209),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_142),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_167),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_177),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_47),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_132),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_237),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_270),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_83),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_189),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_182),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_100),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_4),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_92),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_81),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_156),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_274),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_163),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_207),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_52),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_248),
.B(n_244),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_115),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_47),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_202),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_271),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_223),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_245),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_50),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_234),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_121),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_18),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_221),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_184),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_54),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_263),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_66),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_80),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_256),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_162),
.Y(n_391)
);

BUFx2_ASAP7_75t_SL g392 ( 
.A(n_36),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_107),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_216),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_168),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_86),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_85),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_58),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_241),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_169),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_279),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_91),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_243),
.B(n_235),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_135),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_212),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_49),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_74),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_157),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_205),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_151),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_141),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_155),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_267),
.Y(n_414)
);

BUFx10_ASAP7_75t_L g415 ( 
.A(n_120),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_276),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_246),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_266),
.B(n_211),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_278),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_23),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_222),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_67),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_83),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_149),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_3),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_258),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_253),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_52),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_204),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_215),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_116),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_190),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_194),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_40),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_120),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_109),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_61),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_249),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_87),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_199),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_178),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_238),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_196),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_198),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_213),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_165),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_186),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_62),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_22),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_30),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_13),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_255),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_159),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_11),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_8),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_126),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_160),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_226),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_88),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_59),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_164),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_105),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_145),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_94),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_280),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_240),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_20),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_187),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_268),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_154),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_15),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_130),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_82),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_206),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_32),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_73),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_72),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_31),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_3),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_236),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_95),
.B(n_193),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_58),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_191),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_119),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_138),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_275),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_99),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_87),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_97),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_128),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_51),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_15),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_126),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_8),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_24),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_128),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_74),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_20),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_180),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_99),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_89),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_82),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_188),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_127),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_59),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_43),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_261),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_195),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_72),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_231),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_201),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_282),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_302),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_297),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_283),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_302),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_283),
.B(n_0),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_333),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_292),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_378),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_282),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_361),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_291),
.B(n_0),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_359),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_2),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_297),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_297),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_470),
.B(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_291),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_297),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_344),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_2),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_407),
.B(n_5),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_281),
.B(n_5),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_373),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_407),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_361),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_316),
.Y(n_541)
);

BUFx8_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_379),
.Y(n_543)
);

BUFx12f_ASAP7_75t_L g544 ( 
.A(n_359),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_344),
.B(n_7),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_425),
.B(n_7),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_415),
.B(n_9),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_425),
.B(n_9),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_415),
.B(n_359),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_385),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_10),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_379),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_444),
.A2(n_136),
.B(n_134),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_385),
.B(n_10),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_320),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_304),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_340),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_383),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_385),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_316),
.B(n_139),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_299),
.B(n_11),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_320),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_376),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_383),
.B(n_12),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_511),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_500),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_417),
.B(n_12),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_286),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_304),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_288),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_351),
.A2(n_19),
.B1(n_14),
.B2(n_17),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_388),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_376),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_289),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_290),
.A2(n_143),
.B(n_140),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_393),
.B(n_14),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_376),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_459),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_308),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_441),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_584)
);

BUFx12f_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_397),
.B(n_22),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_293),
.B(n_146),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_309),
.A2(n_150),
.B(n_148),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_475),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_23),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_397),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_483),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_458),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_398),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_492),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_458),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_398),
.B(n_24),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_506),
.B(n_25),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_358),
.B(n_25),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_403),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_403),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_458),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_306),
.B(n_29),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_310),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_458),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_315),
.B(n_153),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_471),
.Y(n_609)
);

BUFx12f_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_294),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_317),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_471),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_313),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_318),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_314),
.B(n_319),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_469),
.B(n_33),
.Y(n_617)
);

BUFx6f_ASAP7_75t_SL g618 ( 
.A(n_518),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_518),
.B(n_499),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_525),
.B(n_322),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_518),
.B(n_327),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_515),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_515),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_528),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_590),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_556),
.B(n_591),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_590),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_581),
.B(n_296),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_581),
.B(n_331),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_599),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_559),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_567),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_582),
.B(n_332),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_599),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_524),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_529),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_532),
.Y(n_648)
);

AO21x2_ASAP7_75t_L g649 ( 
.A1(n_588),
.A2(n_418),
.B(n_339),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_532),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_554),
.B(n_294),
.Y(n_651)
);

AO22x2_ASAP7_75t_L g652 ( 
.A1(n_602),
.A2(n_524),
.B1(n_546),
.B2(n_545),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_559),
.B(n_338),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_545),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_546),
.B(n_348),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_573),
.A2(n_324),
.B1(n_420),
.B2(n_307),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_551),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_551),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_549),
.B(n_300),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_556),
.B(n_307),
.Y(n_660)
);

CKINVDCx6p67_ASAP7_75t_R g661 ( 
.A(n_544),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_555),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_559),
.B(n_350),
.Y(n_665)
);

INVx11_ASAP7_75t_L g666 ( 
.A(n_544),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_567),
.B(n_303),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_560),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_562),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_604),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_571),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_562),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_591),
.B(n_301),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_531),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_562),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_563),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_569),
.B(n_352),
.Y(n_677)
);

BUFx6f_ASAP7_75t_SL g678 ( 
.A(n_520),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_570),
.B(n_354),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_594),
.A2(n_335),
.B1(n_353),
.B2(n_312),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_580),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_580),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_572),
.B(n_366),
.Y(n_683)
);

INVx11_ASAP7_75t_L g684 ( 
.A(n_550),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_550),
.B(n_392),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_607),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_575),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_594),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_575),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_576),
.B(n_368),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_616),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_577),
.A2(n_371),
.B(n_370),
.Y(n_694)
);

BUFx10_ASAP7_75t_L g695 ( 
.A(n_521),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_568),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_580),
.B(n_303),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_579),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_560),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_616),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_576),
.B(n_387),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_593),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_534),
.Y(n_703)
);

AND3x2_ASAP7_75t_L g704 ( 
.A(n_538),
.B(n_345),
.C(n_325),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_513),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_568),
.B(n_329),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_560),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_593),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_593),
.Y(n_709)
);

INVx6_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_514),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_514),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_527),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_517),
.Y(n_714)
);

AND2x2_ASAP7_75t_SL g715 ( 
.A(n_587),
.B(n_535),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_585),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_530),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_547),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_585),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_608),
.B(n_471),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_583),
.B(n_390),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_596),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_589),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_527),
.B(n_391),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_608),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_605),
.B(n_394),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_603),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_610),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_608),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_605),
.B(n_401),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_610),
.B(n_334),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_603),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_539),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_606),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_537),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_405),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_542),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_542),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_612),
.B(n_410),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_612),
.B(n_413),
.Y(n_742)
);

AND3x2_ASAP7_75t_L g743 ( 
.A(n_600),
.B(n_396),
.C(n_380),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_609),
.Y(n_744)
);

CKINVDCx11_ASAP7_75t_R g745 ( 
.A(n_615),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_609),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_609),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_615),
.B(n_522),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_609),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_566),
.B(n_414),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_608),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_541),
.B(n_399),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_519),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_703),
.B(n_537),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_692),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_670),
.B(n_537),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_705),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_687),
.B(n_526),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_685),
.B(n_706),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_671),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_713),
.B(n_542),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_619),
.A2(n_578),
.B1(n_598),
.B2(n_586),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_SL g764 ( 
.A(n_618),
.B(n_312),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

BUFx6f_ASAP7_75t_SL g766 ( 
.A(n_706),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_689),
.B(n_548),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_752),
.B(n_617),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_636),
.B(n_600),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_689),
.B(n_548),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_620),
.B(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_620),
.B(n_508),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_637),
.B(n_508),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_647),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_637),
.B(n_509),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_713),
.B(n_536),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_656),
.B(n_611),
.C(n_584),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_642),
.B(n_512),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_647),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_689),
.B(n_284),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_696),
.B(n_601),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_619),
.A2(n_353),
.B1(n_355),
.B2(n_335),
.Y(n_783)
);

BUFx6f_ASAP7_75t_SL g784 ( 
.A(n_706),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_678),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_641),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_651),
.B(n_374),
.C(n_367),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_717),
.B(n_566),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_659),
.B(n_724),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_731),
.B(n_685),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_668),
.B(n_285),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_724),
.B(n_595),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_653),
.B(n_595),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_651),
.B(n_498),
.C(n_423),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_720),
.B(n_553),
.C(n_523),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_733),
.B(n_639),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_695),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_644),
.B(n_519),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_645),
.B(n_523),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_654),
.B(n_540),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_653),
.B(n_595),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_729),
.B(n_287),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_657),
.B(n_543),
.Y(n_804)
);

BUFx6f_ASAP7_75t_SL g805 ( 
.A(n_731),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_665),
.B(n_557),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_707),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_638),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_662),
.B(n_558),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_652),
.A2(n_377),
.B1(n_412),
.B2(n_355),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_720),
.B(n_553),
.C(n_552),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_663),
.B(n_574),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_652),
.A2(n_412),
.B1(n_443),
.B2(n_377),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_695),
.B(n_592),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_677),
.B(n_305),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_597),
.Y(n_816)
);

BUFx5_ASAP7_75t_L g817 ( 
.A(n_725),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_638),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_718),
.B(n_295),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_674),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_685),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_631),
.B(n_298),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_686),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_623),
.B(n_400),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_711),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_712),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_714),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_745),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_751),
.B(n_311),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_655),
.B(n_421),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_677),
.B(n_330),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_621),
.B(n_336),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_622),
.B(n_337),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_655),
.B(n_504),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_745),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_753),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_719),
.B(n_321),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_629),
.B(n_341),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_323),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_635),
.B(n_342),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_666),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_643),
.Y(n_842)
);

AND2x4_ASAP7_75t_SL g843 ( 
.A(n_731),
.B(n_443),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_658),
.B(n_346),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_710),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_736),
.A2(n_741),
.B(n_742),
.C(n_748),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_710),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_716),
.B(n_326),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_R g849 ( 
.A(n_738),
.B(n_464),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_725),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_652),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_715),
.B(n_362),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_715),
.B(n_369),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_667),
.B(n_381),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_649),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_697),
.B(n_384),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_680),
.B(n_328),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_L g858 ( 
.A1(n_735),
.A2(n_420),
.B1(n_428),
.B2(n_324),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_649),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_641),
.B(n_395),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_641),
.B(n_402),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_681),
.B(n_406),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_SL g863 ( 
.A(n_728),
.B(n_409),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_679),
.B(n_347),
.C(n_343),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_682),
.B(n_411),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_723),
.B(n_416),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_750),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_736),
.B(n_349),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_SL g869 ( 
.A(n_684),
.B(n_424),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_750),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_704),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_678),
.A2(n_464),
.B1(n_357),
.B2(n_360),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_SL g873 ( 
.A(n_738),
.B(n_426),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_743),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_660),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_742),
.B(n_565),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_683),
.B(n_356),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_691),
.B(n_565),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_701),
.B(n_419),
.Y(n_879)
);

BUFx5_ASAP7_75t_L g880 ( 
.A(n_694),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_R g881 ( 
.A(n_721),
.B(n_428),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_726),
.A2(n_364),
.B1(n_365),
.B2(n_363),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_726),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_730),
.B(n_372),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_730),
.B(n_427),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_633),
.B(n_429),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_624),
.B(n_430),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_624),
.B(n_432),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_633),
.B(n_433),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_625),
.B(n_431),
.Y(n_890)
);

NOR2x1p5_ASAP7_75t_L g891 ( 
.A(n_625),
.B(n_375),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_627),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_628),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_633),
.B(n_438),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_630),
.A2(n_386),
.B1(n_389),
.B2(n_382),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_630),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_664),
.B(n_439),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_632),
.A2(n_437),
.B1(n_440),
.B2(n_436),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_634),
.B(n_442),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_664),
.B(n_445),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_640),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_846),
.A2(n_451),
.B(n_457),
.C(n_449),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_791),
.B(n_448),
.Y(n_903)
);

AND2x6_ASAP7_75t_L g904 ( 
.A(n_791),
.B(n_462),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_771),
.B(n_408),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_787),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_761),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_798),
.B(n_446),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_787),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_790),
.B(n_502),
.C(n_499),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_842),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_478),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_814),
.B(n_422),
.Y(n_913)
);

CKINVDCx8_ASAP7_75t_R g914 ( 
.A(n_821),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_816),
.B(n_434),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_760),
.B(n_767),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_796),
.A2(n_404),
.B(n_646),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_783),
.A2(n_491),
.B1(n_463),
.B2(n_465),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_807),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_760),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_828),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_776),
.A2(n_468),
.B(n_472),
.C(n_461),
.Y(n_922)
);

NOR2x1_ASAP7_75t_L g923 ( 
.A(n_760),
.B(n_473),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_821),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_758),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_477),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_839),
.B(n_435),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_851),
.A2(n_488),
.B1(n_494),
.B2(n_480),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_821),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_835),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_777),
.A2(n_501),
.B(n_503),
.C(n_496),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_754),
.B(n_447),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_766),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_843),
.B(n_450),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_780),
.B(n_452),
.Y(n_935)
);

AOI222xp33_ASAP7_75t_L g936 ( 
.A1(n_858),
.A2(n_510),
.B1(n_497),
.B2(n_493),
.C1(n_455),
.C2(n_456),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_796),
.A2(n_811),
.B(n_859),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_763),
.B(n_460),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_822),
.B(n_474),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_766),
.Y(n_940)
);

AND2x2_ASAP7_75t_SL g941 ( 
.A(n_810),
.B(n_499),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_755),
.A2(n_485),
.B1(n_489),
.B2(n_476),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_765),
.B(n_490),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_768),
.B(n_453),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_756),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_811),
.A2(n_650),
.B(n_648),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_781),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_820),
.A2(n_499),
.B(n_502),
.C(n_471),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_774),
.B(n_454),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_868),
.B(n_466),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_769),
.A2(n_823),
.B1(n_782),
.B2(n_818),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_757),
.B(n_772),
.Y(n_952)
);

NOR4xp25_ASAP7_75t_SL g953 ( 
.A(n_764),
.B(n_481),
.C(n_484),
.D(n_467),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_757),
.B(n_486),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_774),
.B(n_487),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_773),
.B(n_34),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_808),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_779),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_775),
.B(n_34),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_778),
.B(n_35),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_809),
.A2(n_613),
.B(n_749),
.C(n_669),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_762),
.A2(n_35),
.B(n_37),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_841),
.B(n_38),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_812),
.A2(n_747),
.B(n_675),
.C(n_676),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_789),
.A2(n_676),
.B(n_672),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_877),
.B(n_39),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_799),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_799),
.A2(n_801),
.B(n_800),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_800),
.Y(n_969)
);

AOI21xp33_ASAP7_75t_L g970 ( 
.A1(n_819),
.A2(n_40),
.B(n_41),
.Y(n_970)
);

NOR2x1_ASAP7_75t_R g971 ( 
.A(n_874),
.B(n_42),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_852),
.A2(n_853),
.B1(n_795),
.B2(n_788),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_837),
.B(n_44),
.Y(n_974)
);

BUFx4f_ASAP7_75t_L g975 ( 
.A(n_871),
.Y(n_975)
);

AOI33xp33_ASAP7_75t_L g976 ( 
.A1(n_898),
.A2(n_746),
.A3(n_744),
.B1(n_740),
.B2(n_739),
.B3(n_734),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_793),
.A2(n_690),
.B(n_688),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_884),
.B(n_46),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_L g979 ( 
.A(n_864),
.B(n_698),
.C(n_693),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_844),
.A2(n_702),
.B(n_698),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_826),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_891),
.B(n_786),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_824),
.B(n_49),
.Y(n_983)
);

NOR2x2_ASAP7_75t_L g984 ( 
.A(n_849),
.B(n_784),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_857),
.A2(n_702),
.B(n_708),
.C(n_709),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_L g986 ( 
.A(n_875),
.B(n_874),
.C(n_872),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_830),
.B(n_50),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_883),
.A2(n_870),
.B(n_867),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_832),
.A2(n_838),
.B(n_833),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_825),
.A2(n_722),
.B1(n_734),
.B2(n_732),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_834),
.B(n_51),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_806),
.B(n_53),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_840),
.A2(n_709),
.B(n_708),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_836),
.A2(n_722),
.B1(n_732),
.B2(n_727),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_797),
.B(n_784),
.Y(n_995)
);

NOR2x2_ASAP7_75t_L g996 ( 
.A(n_805),
.B(n_54),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_881),
.Y(n_997)
);

OA22x2_ASAP7_75t_L g998 ( 
.A1(n_805),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_848),
.B(n_55),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_827),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_873),
.B(n_60),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_794),
.B(n_62),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_882),
.B(n_64),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_SL g1004 ( 
.A(n_817),
.B(n_161),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_802),
.B(n_65),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_876),
.B(n_65),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_879),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_862),
.B(n_68),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_831),
.B(n_69),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_879),
.A2(n_70),
.B(n_71),
.C(n_73),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_873),
.B(n_71),
.Y(n_1011)
);

OAI321xp33_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_75),
.A3(n_76),
.B1(n_77),
.B2(n_78),
.C(n_79),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_878),
.A2(n_75),
.B(n_78),
.C(n_79),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_890),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_888),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_885),
.B(n_81),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_845),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_895),
.B(n_84),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_866),
.B(n_84),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_890),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_886),
.A2(n_897),
.B(n_829),
.C(n_856),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_815),
.A2(n_86),
.B(n_89),
.Y(n_1022)
);

AND2x2_ASAP7_75t_SL g1023 ( 
.A(n_860),
.B(n_90),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_854),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_869),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_850),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_L g1027 ( 
.A(n_865),
.B(n_90),
.C(n_92),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_861),
.A2(n_93),
.B(n_94),
.C(n_96),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_893),
.A2(n_896),
.B(n_901),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_847),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_889),
.A2(n_894),
.B(n_900),
.C(n_899),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_863),
.B(n_96),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_803),
.A2(n_203),
.B(n_264),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_792),
.A2(n_197),
.B(n_262),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_L g1035 ( 
.A(n_817),
.B(n_173),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_785),
.B(n_98),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_892),
.A2(n_98),
.B(n_100),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_880),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_912),
.B(n_907),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_924),
.B(n_101),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_914),
.Y(n_1041)
);

AOI211x1_ASAP7_75t_L g1042 ( 
.A1(n_1022),
.A2(n_102),
.B(n_104),
.C(n_105),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_997),
.Y(n_1043)
);

BUFx8_ASAP7_75t_L g1044 ( 
.A(n_1025),
.Y(n_1044)
);

NAND2x2_ASAP7_75t_L g1045 ( 
.A(n_945),
.B(n_106),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_951),
.B(n_110),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_971),
.B(n_110),
.C(n_111),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_926),
.B(n_112),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_941),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_924),
.B(n_113),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_938),
.A2(n_114),
.B(n_115),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_924),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_916),
.B(n_116),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_951),
.B(n_117),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_902),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_931),
.A2(n_118),
.B(n_121),
.C(n_122),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_905),
.B(n_122),
.Y(n_1057)
);

BUFx2_ASAP7_75t_SL g1058 ( 
.A(n_933),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_922),
.B(n_123),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_1014),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_988),
.A2(n_123),
.B(n_124),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1038),
.A2(n_124),
.B(n_125),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_926),
.B(n_125),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_927),
.B(n_935),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_903),
.B(n_127),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1006),
.A2(n_130),
.B(n_131),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_933),
.B(n_131),
.Y(n_1067)
);

AND2x2_ASAP7_75t_SL g1068 ( 
.A(n_920),
.B(n_181),
.Y(n_1068)
);

AOI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_939),
.A2(n_966),
.B(n_934),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_940),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

AOI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_950),
.A2(n_985),
.B(n_954),
.Y(n_1072)
);

AOI221x1_ASAP7_75t_L g1073 ( 
.A1(n_910),
.A2(n_1027),
.B1(n_962),
.B2(n_970),
.C(n_1037),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_974),
.A2(n_959),
.B(n_956),
.C(n_960),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1020),
.A2(n_972),
.B1(n_992),
.B2(n_978),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1000),
.Y(n_1076)
);

AND2x6_ASAP7_75t_L g1077 ( 
.A(n_906),
.B(n_909),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_903),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1031),
.A2(n_977),
.B(n_1029),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_975),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_983),
.A2(n_987),
.B(n_991),
.C(n_1007),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_904),
.B(n_972),
.Y(n_1082)
);

BUFx2_ASAP7_75t_SL g1083 ( 
.A(n_940),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1000),
.A2(n_944),
.B1(n_1005),
.B2(n_1002),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_929),
.B(n_916),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_977),
.A2(n_993),
.B(n_980),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1023),
.B(n_936),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1010),
.A2(n_1028),
.B(n_1013),
.C(n_1016),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_1004),
.A2(n_1035),
.B(n_1036),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_923),
.B(n_1024),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_930),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_965),
.A2(n_915),
.B(n_913),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_975),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_947),
.Y(n_1094)
);

AND3x1_ASAP7_75t_SL g1095 ( 
.A(n_984),
.B(n_996),
.C(n_986),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_995),
.A2(n_943),
.B(n_932),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_919),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_904),
.B(n_928),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_942),
.A2(n_999),
.B1(n_921),
.B2(n_982),
.C(n_1018),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1008),
.B(n_1019),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1003),
.A2(n_979),
.B(n_976),
.C(n_957),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1008),
.B(n_1019),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_982),
.B(n_1017),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_925),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_998),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1001),
.B(n_1011),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_948),
.A2(n_1034),
.B(n_1033),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1032),
.A2(n_1009),
.B1(n_1021),
.B2(n_1012),
.C(n_908),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_953),
.Y(n_1109)
);

OAI22x1_ASAP7_75t_L g1110 ( 
.A1(n_1012),
.A2(n_953),
.B1(n_963),
.B2(n_1030),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_990),
.A2(n_994),
.B(n_961),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_958),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_949),
.B(n_955),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_937),
.A2(n_946),
.B(n_859),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_912),
.B(n_759),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_967),
.B(n_969),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_967),
.B(n_969),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_1027),
.B(n_910),
.C(n_917),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_989),
.A2(n_952),
.B(n_902),
.C(n_968),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_917),
.A2(n_937),
.B(n_910),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_967),
.B(n_969),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1026),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_924),
.B(n_920),
.Y(n_1123)
);

AND2x6_ASAP7_75t_SL g1124 ( 
.A(n_999),
.B(n_760),
.Y(n_1124)
);

AOI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_952),
.A2(n_754),
.B(n_737),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_912),
.B(n_759),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_967),
.B(n_969),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_967),
.B(n_969),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_903),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1022),
.A2(n_855),
.A3(n_859),
.B(n_964),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_L g1131 ( 
.A(n_1027),
.B(n_910),
.C(n_917),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_967),
.B(n_969),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_907),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_967),
.A2(n_969),
.B1(n_973),
.B2(n_1015),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1027),
.B(n_910),
.C(n_917),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_912),
.B(n_759),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_967),
.B(n_969),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_952),
.B(n_902),
.C(n_968),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_907),
.B(n_798),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_967),
.A2(n_969),
.B1(n_973),
.B2(n_1015),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_967),
.B(n_969),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_907),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_969),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_902),
.A2(n_931),
.B1(n_922),
.B2(n_968),
.C(n_846),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_L g1145 ( 
.A(n_903),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_924),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_907),
.Y(n_1147)
);

AND3x4_ASAP7_75t_L g1148 ( 
.A(n_986),
.B(n_777),
.C(n_791),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_967),
.A2(n_969),
.B1(n_973),
.B2(n_1015),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_967),
.B(n_969),
.Y(n_1150)
);

OA22x2_ASAP7_75t_L g1151 ( 
.A1(n_918),
.A2(n_810),
.B1(n_813),
.B2(n_680),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_945),
.Y(n_1152)
);

BUFx4f_ASAP7_75t_L g1153 ( 
.A(n_903),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_967),
.B(n_969),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_SL g1155 ( 
.A1(n_968),
.A2(n_798),
.B(n_1022),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_912),
.B(n_759),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_941),
.A2(n_777),
.B1(n_652),
.B2(n_952),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_907),
.B(n_798),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_924),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_907),
.B(n_761),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_981),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_941),
.A2(n_777),
.B1(n_912),
.B2(n_918),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_924),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_945),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_933),
.B(n_756),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_967),
.B(n_969),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_912),
.B(n_687),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_945),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1133),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1171)
);

AOI22x1_ASAP7_75t_L g1172 ( 
.A1(n_1110),
.A2(n_1109),
.B1(n_1155),
.B2(n_1092),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1079),
.A2(n_1086),
.B(n_1114),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1163),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1163),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1162),
.A2(n_1151),
.B1(n_1087),
.B2(n_1148),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1044),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1160),
.A2(n_1157),
.B1(n_1156),
.B2(n_1136),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1070),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1071),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1163),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1039),
.B(n_1064),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1133),
.B(n_1147),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1121),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_SL g1186 ( 
.A(n_1044),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1125),
.B(n_1167),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_1108),
.B(n_1042),
.C(n_1074),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1127),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_1142),
.B(n_1080),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1128),
.B(n_1132),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_SL g1192 ( 
.A(n_1041),
.Y(n_1192)
);

AO21x2_ASAP7_75t_L g1193 ( 
.A1(n_1120),
.A2(n_1111),
.B(n_1118),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1118),
.A2(n_1135),
.B(n_1131),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_1131),
.A2(n_1135),
.B(n_1101),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1145),
.B(n_1153),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1069),
.A2(n_1075),
.B(n_1084),
.C(n_1056),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1157),
.B1(n_1147),
.B2(n_1040),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1137),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1073),
.A2(n_1061),
.B(n_1062),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1055),
.A2(n_1140),
.B(n_1149),
.C(n_1057),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1141),
.B(n_1143),
.Y(n_1202)
);

NAND2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1145),
.B(n_1153),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1150),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1094),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1078),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1154),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1107),
.A2(n_1072),
.B(n_1061),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1123),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1078),
.B(n_1068),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1062),
.A2(n_1082),
.B(n_1066),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_1054),
.B(n_1046),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1052),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1166),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1152),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

OAI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1099),
.A2(n_1049),
.B1(n_1105),
.B2(n_1096),
.C(n_1144),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1164),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1098),
.A2(n_1065),
.B(n_1159),
.Y(n_1219)
);

BUFx2_ASAP7_75t_R g1220 ( 
.A(n_1093),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1063),
.B(n_1053),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1146),
.B(n_1043),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1051),
.A2(n_1106),
.B(n_1059),
.Y(n_1223)
);

NOR2x1_ASAP7_75t_R g1224 ( 
.A(n_1058),
.B(n_1083),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1076),
.A2(n_1161),
.B(n_1130),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1060),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1078),
.A2(n_1053),
.B1(n_1048),
.B2(n_1067),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1113),
.A2(n_1130),
.B(n_1165),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1067),
.A2(n_1085),
.B1(n_1040),
.B2(n_1050),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1050),
.A2(n_1090),
.B1(n_1095),
.B2(n_1067),
.Y(n_1230)
);

AND2x6_ASAP7_75t_L g1231 ( 
.A(n_1122),
.B(n_1112),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1130),
.A2(n_1112),
.B(n_1158),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_1047),
.B(n_1139),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1085),
.B(n_1168),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1091),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_R g1236 ( 
.A(n_1124),
.B(n_1103),
.Y(n_1236)
);

AOI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1097),
.A2(n_1090),
.B1(n_1060),
.B2(n_1103),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1085),
.B(n_1124),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1045),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1077),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1077),
.B(n_1116),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1077),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1163),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_SL g1245 ( 
.A(n_1163),
.B(n_914),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1134),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1108),
.B(n_1042),
.C(n_1074),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1116),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1163),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_SL g1251 ( 
.A1(n_1062),
.A2(n_1061),
.B(n_1134),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1108),
.B(n_1042),
.C(n_1074),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1163),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1078),
.B(n_1123),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1044),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1079),
.A2(n_1089),
.A3(n_1138),
.B(n_1119),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1116),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1163),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1071),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1163),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1088),
.A2(n_952),
.B(n_1081),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1044),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1116),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1163),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1116),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1115),
.B(n_1126),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1163),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1185),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1185),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1189),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1199),
.B(n_1204),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1204),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1171),
.B(n_1246),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1207),
.B(n_1249),
.Y(n_1279)
);

NAND2x1_ASAP7_75t_L g1280 ( 
.A(n_1219),
.B(n_1231),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1171),
.B(n_1256),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1258),
.B(n_1249),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1242),
.B(n_1175),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1266),
.B(n_1269),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1260),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

AOI221xp5_ASAP7_75t_L g1287 ( 
.A1(n_1187),
.A2(n_1177),
.B1(n_1217),
.B2(n_1259),
.C(n_1170),
.Y(n_1287)
);

AOI222xp33_ASAP7_75t_L g1288 ( 
.A1(n_1177),
.A2(n_1261),
.B1(n_1271),
.B2(n_1236),
.C1(n_1186),
.C2(n_1187),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1247),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1216),
.Y(n_1290)
);

BUFx2_ASAP7_75t_R g1291 ( 
.A(n_1178),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1173),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1175),
.B(n_1191),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1184),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_SL g1295 ( 
.A1(n_1251),
.A2(n_1229),
.B(n_1227),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1175),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1230),
.B(n_1221),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1198),
.A2(n_1210),
.B1(n_1179),
.B2(n_1191),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1268),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1205),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1268),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1268),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1174),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1270),
.B(n_1242),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1231),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1181),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_1265),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1202),
.A2(n_1247),
.B1(n_1214),
.B2(n_1206),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1264),
.B(n_1170),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1169),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1257),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1242),
.A2(n_1238),
.B1(n_1206),
.B2(n_1186),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1226),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1262),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1257),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1180),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1265),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1257),
.Y(n_1318)
);

BUFx2_ASAP7_75t_SL g1319 ( 
.A(n_1174),
.Y(n_1319)
);

CKINVDCx14_ASAP7_75t_R g1320 ( 
.A(n_1178),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1254),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1192),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1226),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1235),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1231),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1183),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1176),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1286),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1324),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1280),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1276),
.B(n_1194),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1276),
.B(n_1194),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1286),
.Y(n_1333)
);

OAI222xp33_ASAP7_75t_L g1334 ( 
.A1(n_1308),
.A2(n_1237),
.B1(n_1254),
.B2(n_1197),
.C1(n_1245),
.C2(n_1234),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1282),
.B(n_1193),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1283),
.B(n_1232),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1280),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1279),
.B(n_1284),
.Y(n_1338)
);

NOR2x1_ASAP7_75t_L g1339 ( 
.A(n_1305),
.B(n_1188),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1309),
.B(n_1287),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1317),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1274),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1288),
.A2(n_1233),
.B1(n_1248),
.B2(n_1252),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1309),
.B(n_1233),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1279),
.B(n_1239),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1326),
.B(n_1294),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1323),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1293),
.A2(n_1211),
.B1(n_1212),
.B2(n_1223),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1293),
.B(n_1194),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1295),
.A2(n_1319),
.B1(n_1321),
.B2(n_1283),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1290),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1298),
.A2(n_1254),
.B1(n_1222),
.B2(n_1240),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1323),
.Y(n_1354)
);

INVx5_ASAP7_75t_SL g1355 ( 
.A(n_1316),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1273),
.B(n_1195),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1289),
.B(n_1228),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1313),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1275),
.B(n_1195),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1275),
.B(n_1211),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1295),
.A2(n_1240),
.B1(n_1172),
.B2(n_1176),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1319),
.A2(n_1244),
.B1(n_1272),
.B2(n_1182),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1277),
.B(n_1208),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1344),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1328),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1340),
.A2(n_1283),
.B1(n_1297),
.B2(n_1299),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1328),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1333),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1348),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1338),
.B(n_1300),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1350),
.B(n_1331),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1350),
.B(n_1315),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1358),
.Y(n_1374)
);

AOI222xp33_ASAP7_75t_L g1375 ( 
.A1(n_1343),
.A2(n_1224),
.B1(n_1281),
.B2(n_1278),
.C1(n_1317),
.C2(n_1314),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1331),
.B(n_1315),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1332),
.B(n_1318),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1332),
.B(n_1318),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1351),
.A2(n_1312),
.B1(n_1307),
.B2(n_1321),
.C(n_1234),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1341),
.B(n_1322),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1338),
.B(n_1296),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1335),
.B(n_1310),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1341),
.B(n_1316),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1354),
.B(n_1277),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1330),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1354),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1352),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1347),
.B(n_1300),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1329),
.B(n_1306),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1342),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1352),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1383),
.B(n_1360),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1391),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1387),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1372),
.B(n_1356),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1365),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1383),
.B(n_1357),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1375),
.B(n_1362),
.C(n_1339),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1366),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1366),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1368),
.B(n_1356),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1377),
.B(n_1336),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1372),
.B(n_1359),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1377),
.B(n_1355),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1368),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1380),
.B(n_1339),
.C(n_1346),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1364),
.B(n_1357),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1373),
.B(n_1359),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1373),
.B(n_1363),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1387),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1369),
.B(n_1363),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1367),
.A2(n_1299),
.B1(n_1301),
.B2(n_1302),
.Y(n_1413)
);

AND2x4_ASAP7_75t_SL g1414 ( 
.A(n_1382),
.B(n_1330),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1369),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1396),
.B(n_1374),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1397),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1396),
.B(n_1376),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1410),
.B(n_1371),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1409),
.B(n_1378),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1399),
.A2(n_1341),
.B1(n_1381),
.B2(n_1353),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1400),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1399),
.B(n_1390),
.C(n_1384),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1409),
.B(n_1370),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1400),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1414),
.B(n_1378),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1408),
.B(n_1364),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1414),
.B(n_1379),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1401),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1407),
.A2(n_1334),
.B(n_1190),
.Y(n_1433)
);

NOR3xp33_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1361),
.C(n_1201),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1414),
.B(n_1379),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1424),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1425),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1423),
.A2(n_1405),
.B1(n_1341),
.B2(n_1395),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1429),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1434),
.A2(n_1413),
.B1(n_1336),
.B2(n_1403),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1417),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1429),
.B(n_1419),
.Y(n_1442)
);

INVx3_ASAP7_75t_SL g1443 ( 
.A(n_1428),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1428),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1416),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1418),
.B(n_1395),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1435),
.B(n_1403),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1417),
.Y(n_1448)
);

OAI221xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1426),
.A2(n_1413),
.B1(n_1398),
.B2(n_1408),
.C(n_1393),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_SL g1450 ( 
.A(n_1433),
.B(n_1255),
.C(n_1398),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1424),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1418),
.B(n_1394),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1427),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1403),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1420),
.B(n_1403),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1430),
.A2(n_1412),
.B1(n_1393),
.B2(n_1402),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1443),
.A2(n_1435),
.B1(n_1421),
.B2(n_1420),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1443),
.A2(n_1444),
.B1(n_1454),
.B2(n_1449),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1437),
.A2(n_1386),
.B(n_1285),
.Y(n_1459)
);

OA222x2_ASAP7_75t_L g1460 ( 
.A1(n_1442),
.A2(n_1411),
.B1(n_1387),
.B2(n_1337),
.C1(n_1385),
.C2(n_1355),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1450),
.A2(n_1422),
.B1(n_1431),
.B2(n_1427),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1440),
.A2(n_1422),
.B1(n_1432),
.B2(n_1431),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_R g1463 ( 
.A1(n_1442),
.A2(n_1389),
.B(n_1412),
.C(n_1402),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1451),
.Y(n_1464)
);

OAI31xp33_ASAP7_75t_L g1465 ( 
.A1(n_1438),
.A2(n_1411),
.A3(n_1432),
.B(n_1304),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1445),
.A2(n_1415),
.B1(n_1406),
.B2(n_1392),
.C(n_1388),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1439),
.A2(n_1444),
.B1(n_1452),
.B2(n_1456),
.C(n_1446),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1446),
.A2(n_1320),
.B(n_1255),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1457),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1464),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1466),
.B(n_1467),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1461),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1458),
.A2(n_1447),
.B1(n_1455),
.B2(n_1355),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1462),
.A2(n_1455),
.B(n_1447),
.Y(n_1474)
);

NAND4xp25_ASAP7_75t_L g1475 ( 
.A(n_1465),
.B(n_1215),
.C(n_1218),
.D(n_1213),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1460),
.A2(n_1411),
.B1(n_1349),
.B2(n_1436),
.C(n_1453),
.Y(n_1476)
);

XNOR2xp5_ASAP7_75t_L g1477 ( 
.A(n_1468),
.B(n_1447),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1459),
.A2(n_1436),
.B(n_1337),
.C(n_1327),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1463),
.A2(n_1355),
.B1(n_1448),
.B2(n_1441),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1464),
.Y(n_1480)
);

AOI211xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1458),
.A2(n_1192),
.B(n_1337),
.C(n_1325),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1470),
.Y(n_1482)
);

NOR2x1_ASAP7_75t_L g1483 ( 
.A(n_1475),
.B(n_1182),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1480),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1469),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1476),
.A2(n_1291),
.B1(n_1377),
.B2(n_1304),
.Y(n_1486)
);

AND4x1_ASAP7_75t_L g1487 ( 
.A(n_1481),
.B(n_1180),
.C(n_1220),
.D(n_1241),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1477),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1473),
.B(n_1180),
.C(n_1215),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1472),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_L g1491 ( 
.A(n_1475),
.B(n_1244),
.Y(n_1491)
);

AOI211xp5_ASAP7_75t_L g1492 ( 
.A1(n_1486),
.A2(n_1471),
.B(n_1474),
.C(n_1478),
.Y(n_1492)
);

AND2x2_ASAP7_75t_SL g1493 ( 
.A(n_1487),
.B(n_1479),
.Y(n_1493)
);

AOI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1486),
.A2(n_1218),
.B(n_1272),
.C(n_1267),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_SL g1495 ( 
.A(n_1488),
.B(n_1203),
.C(n_1196),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1485),
.B(n_1441),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1490),
.B(n_1448),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1489),
.A2(n_1263),
.B(n_1250),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1484),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1415),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1499),
.B(n_1483),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1496),
.Y(n_1502)
);

NOR4xp75_ASAP7_75t_L g1503 ( 
.A(n_1495),
.B(n_1491),
.C(n_1285),
.D(n_1209),
.Y(n_1503)
);

NOR2x1_ASAP7_75t_L g1504 ( 
.A(n_1497),
.B(n_1267),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1500),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1498),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1493),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1492),
.B(n_1406),
.Y(n_1508)
);

NAND4xp75_ASAP7_75t_L g1509 ( 
.A(n_1494),
.B(n_1223),
.C(n_1200),
.D(n_1243),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1502),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_L g1511 ( 
.A(n_1507),
.B(n_1253),
.C(n_1213),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_L g1512 ( 
.A(n_1506),
.B(n_1196),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1503),
.B(n_1234),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1501),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1510),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1514),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1511),
.B(n_1504),
.Y(n_1517)
);

XNOR2xp5_ASAP7_75t_L g1518 ( 
.A(n_1516),
.B(n_1513),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1518),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1518),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1520),
.A2(n_1517),
.B1(n_1512),
.B2(n_1513),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1521),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1522),
.B(n_1519),
.Y(n_1523)
);

OAI21xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1523),
.A2(n_1515),
.B(n_1505),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1524),
.B(n_1517),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1525),
.A2(n_1508),
.B1(n_1509),
.B2(n_1303),
.Y(n_1526)
);


endmodule