module fake_netlist_1_5728_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x2_ASAP7_75t_SL g3 ( .A(n_2), .B(n_0), .Y(n_3) );
CKINVDCx20_ASAP7_75t_R g4 ( .A(n_1), .Y(n_4) );
AOI21xp5_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
INVx2_ASAP7_75t_SL g6 ( .A(n_5), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_6), .B(n_3), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
OAI22x1_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_4), .B1(n_1), .B2(n_0), .Y(n_10) );
XNOR2x1_ASAP7_75t_L g11 ( .A(n_10), .B(n_2), .Y(n_11) );
endmodule