module real_aes_17901_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_18;
NOR3xp33_ASAP7_75t_SL g13 ( .A(n_0), .B(n_5), .C(n_14), .Y(n_13) );
NOR5xp2_ASAP7_75t_SL g11 ( .A(n_1), .B(n_7), .C(n_12), .D(n_16), .E(n_17), .Y(n_11) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_2), .B(n_19), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_4), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g10 ( .A(n_11), .B(n_18), .Y(n_10) );
NAND2xp33_ASAP7_75t_R g12 ( .A(n_13), .B(n_15), .Y(n_12) );
endmodule