module fake_jpeg_8048_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_32),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_18),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_58),
.B1(n_67),
.B2(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_59),
.B1(n_25),
.B2(n_24),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_64),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_19),
.B1(n_30),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_34),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_30),
.B1(n_23),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_30),
.B1(n_25),
.B2(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_35),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_106),
.B1(n_60),
.B2(n_68),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_27),
.B(n_45),
.C(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_89),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_87),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_47),
.B1(n_68),
.B2(n_22),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_82),
.Y(n_133)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_43),
.C(n_40),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_102),
.C(n_105),
.Y(n_132)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_90),
.B1(n_94),
.B2(n_97),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_93),
.Y(n_123)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_29),
.B(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_100),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_47),
.B1(n_31),
.B2(n_20),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_31),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_107),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_36),
.B(n_21),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_47),
.B1(n_21),
.B2(n_36),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_36),
.B1(n_21),
.B2(n_47),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_54),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_98),
.B1(n_80),
.B2(n_78),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_136),
.Y(n_148)
);

AO21x2_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_37),
.B(n_52),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_52),
.B(n_57),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_35),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_15),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_37),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_37),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_60),
.B1(n_83),
.B2(n_87),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_76),
.B1(n_102),
.B2(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_147),
.B1(n_158),
.B2(n_170),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_97),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_127),
.B(n_129),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_145),
.B(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_155),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_84),
.C(n_37),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_113),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_46),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_123),
.B(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_78),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_93),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_46),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_37),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_103),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_46),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_0),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_173),
.B(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_103),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_115),
.B(n_38),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_98),
.B1(n_46),
.B2(n_38),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_38),
.B1(n_57),
.B2(n_70),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_135),
.B1(n_100),
.B2(n_109),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_14),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_28),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_176),
.C(n_168),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_132),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_131),
.A3(n_127),
.B1(n_122),
.B2(n_133),
.C1(n_126),
.C2(n_135),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_186),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_178),
.A2(n_180),
.B(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_191),
.B1(n_192),
.B2(n_195),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_204),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_141),
.B1(n_130),
.B2(n_116),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_116),
.B1(n_126),
.B2(n_139),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_116),
.B1(n_124),
.B2(n_57),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_22),
.B(n_26),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_124),
.B1(n_70),
.B2(n_28),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_206),
.B1(n_169),
.B2(n_174),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_156),
.A2(n_22),
.B(n_26),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_143),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_124),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_28),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_207),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_35),
.B1(n_26),
.B2(n_99),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_213),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_215),
.C(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_188),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_159),
.B1(n_158),
.B2(n_167),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_231),
.B1(n_179),
.B2(n_195),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_142),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_197),
.B1(n_181),
.B2(n_173),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_201),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_162),
.CI(n_142),
.CON(n_220),
.SN(n_220)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_164),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_222),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_151),
.Y(n_222)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_233),
.C(n_196),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_163),
.C(n_145),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_230),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_172),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_179),
.A2(n_173),
.B1(n_165),
.B2(n_145),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_181),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_165),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_235),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_240),
.B1(n_250),
.B2(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_173),
.B1(n_187),
.B2(n_184),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_218),
.C(n_225),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_180),
.B1(n_198),
.B2(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_182),
.CI(n_184),
.CON(n_248),
.SN(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_234),
.B1(n_229),
.B2(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_202),
.B1(n_206),
.B2(n_199),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_200),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_234),
.A2(n_202),
.B1(n_199),
.B2(n_99),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_101),
.B1(n_35),
.B2(n_22),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_262),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_215),
.C(n_224),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_268),
.C(n_271),
.Y(n_282)
);

OAI322xp33_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_227),
.A3(n_210),
.B1(n_221),
.B2(n_212),
.C1(n_220),
.C2(n_211),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_272),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_210),
.B(n_216),
.C(n_8),
.D(n_9),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_270),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_7),
.C(n_12),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_6),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_1),
.C(n_2),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_6),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_8),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_274),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_1),
.C(n_2),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_237),
.B1(n_249),
.B2(n_246),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_285),
.B1(n_258),
.B2(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_269),
.B1(n_257),
.B2(n_255),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_236),
.B(n_242),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_279),
.B(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_241),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_239),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_5),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_273),
.B1(n_236),
.B2(n_264),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_288),
.B1(n_11),
.B2(n_5),
.Y(n_309)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_302),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_260),
.B1(n_248),
.B2(n_265),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_298),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_265),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_9),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_5),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_11),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_282),
.C(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_282),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_301),
.C(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_296),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_293),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_319),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_12),
.B(n_14),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_322),
.B(n_308),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_323),
.B(n_309),
.C(n_318),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_315),
.B(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_321),
.C(n_307),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_317),
.B(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_4),
.Y(n_331)
);


endmodule