module real_aes_2717_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_503;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_958;
wire n_677;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_1078;
wire n_1072;
wire n_744;
wire n_938;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_976;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_656;
wire n_532;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_860;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_455;
wire n_973;
wire n_504;
wire n_725;
wire n_1081;
wire n_1084;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_1031;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_703;
wire n_652;
wire n_601;
wire n_500;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1101;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_0), .A2(n_72), .B1(n_454), .B2(n_660), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_1), .A2(n_126), .B1(n_691), .B2(n_692), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_2), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_3), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_4), .A2(n_262), .B1(n_464), .B2(n_748), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_5), .A2(n_80), .B1(n_442), .B2(n_855), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_6), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_7), .A2(n_357), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_8), .A2(n_70), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_9), .A2(n_56), .B1(n_525), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_10), .A2(n_391), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_11), .A2(n_254), .B1(n_762), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_12), .A2(n_264), .B1(n_485), .B2(n_488), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_13), .A2(n_268), .B1(n_660), .B2(n_715), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_14), .A2(n_315), .B1(n_497), .B2(n_597), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g1053 ( .A1(n_15), .A2(n_331), .B1(n_576), .B2(n_747), .Y(n_1053) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_16), .A2(n_85), .B1(n_509), .B2(n_512), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_17), .A2(n_137), .B1(n_454), .B2(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_18), .A2(n_190), .B1(n_464), .B2(n_521), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_19), .A2(n_346), .B1(n_414), .B2(n_430), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_20), .A2(n_196), .B1(n_751), .B2(n_810), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_21), .A2(n_267), .B1(n_414), .B2(n_430), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_22), .B(n_584), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_23), .A2(n_97), .B1(n_576), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_24), .A2(n_227), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_25), .A2(n_296), .B1(n_827), .B2(n_860), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_26), .A2(n_146), .B1(n_802), .B2(n_803), .Y(n_998) );
INVx1_ASAP7_75t_SL g425 ( .A(n_27), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_27), .B(n_45), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_28), .A2(n_282), .B1(n_501), .B2(n_505), .Y(n_500) );
AOI22xp5_ASAP7_75t_SL g1056 ( .A1(n_29), .A2(n_271), .B1(n_488), .B2(n_638), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g878 ( .A1(n_30), .A2(n_324), .B1(n_363), .B2(n_434), .C1(n_728), .C2(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_31), .B(n_675), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_32), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_33), .A2(n_356), .B1(n_568), .B2(n_635), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_34), .A2(n_38), .B1(n_523), .B2(n_576), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_35), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_36), .A2(n_225), .B1(n_630), .B2(n_633), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_37), .A2(n_313), .B1(n_503), .B2(n_620), .Y(n_619) );
XNOR2x1_ASAP7_75t_SL g972 ( .A(n_39), .B(n_973), .Y(n_972) );
AOI22xp5_ASAP7_75t_SL g1006 ( .A1(n_39), .A2(n_973), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
INVx1_ASAP7_75t_L g1008 ( .A(n_39), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_40), .A2(n_276), .B1(n_510), .B2(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_41), .A2(n_107), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_42), .A2(n_103), .B1(n_695), .B2(n_696), .Y(n_694) );
OA21x2_ASAP7_75t_L g890 ( .A1(n_43), .A2(n_891), .B(n_910), .Y(n_890) );
INVx1_ASAP7_75t_L g912 ( .A(n_43), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_44), .A2(n_101), .B1(n_638), .B2(n_699), .Y(n_813) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_45), .A2(n_368), .B1(n_417), .B2(n_429), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_46), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_47), .A2(n_309), .B1(n_477), .B2(n_478), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_48), .A2(n_108), .B1(n_699), .B2(n_1004), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_49), .B(n_1098), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_50), .A2(n_195), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_51), .A2(n_95), .B1(n_477), .B2(n_478), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_52), .A2(n_292), .B1(n_494), .B2(n_869), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_53), .A2(n_114), .B1(n_574), .B2(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_54), .A2(n_295), .B1(n_800), .B2(n_853), .Y(n_996) );
INVx1_ASAP7_75t_L g426 ( .A(n_55), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_57), .A2(n_358), .B1(n_588), .B2(n_678), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_58), .A2(n_197), .B1(n_352), .B2(n_529), .C1(n_532), .C2(n_535), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_59), .A2(n_260), .B1(n_475), .B2(n_668), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_60), .A2(n_116), .B1(n_509), .B2(n_512), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_61), .B(n_552), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_62), .A2(n_285), .B1(n_622), .B2(n_623), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_63), .A2(n_337), .B1(n_477), .B2(n_478), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_64), .A2(n_99), .B1(n_520), .B2(n_523), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_65), .A2(n_118), .B1(n_832), .B2(n_833), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_66), .A2(n_141), .B1(n_591), .B2(n_761), .Y(n_760) );
AO222x2_ASAP7_75t_SL g935 ( .A1(n_67), .A2(n_121), .B1(n_170), .B2(n_414), .C1(n_430), .C2(n_435), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_68), .A2(n_394), .B1(n_512), .B2(n_622), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_69), .A2(n_310), .B1(n_442), .B2(n_505), .Y(n_964) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_71), .A2(n_203), .B1(n_417), .B2(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_73), .A2(n_338), .B1(n_526), .B2(n_860), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_74), .A2(n_78), .B1(n_470), .B2(n_790), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_75), .B(n_764), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_76), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_77), .A2(n_163), .B1(n_475), .B2(n_668), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_79), .A2(n_294), .B1(n_660), .B2(n_715), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_81), .A2(n_128), .B1(n_497), .B2(n_598), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_82), .A2(n_202), .B1(n_503), .B2(n_620), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_83), .A2(n_278), .B1(n_464), .B2(n_527), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_84), .B(n_434), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_86), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_87), .A2(n_290), .B1(n_470), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_88), .A2(n_300), .B1(n_492), .B2(n_497), .Y(n_491) );
AO22x1_ASAP7_75t_L g897 ( .A1(n_89), .A2(n_263), .B1(n_587), .B2(n_591), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_90), .A2(n_396), .B1(n_475), .B2(n_668), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_91), .A2(n_259), .B1(n_758), .B2(n_766), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_92), .A2(n_272), .B1(n_464), .B2(n_471), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_93), .A2(n_344), .B1(n_809), .B2(n_810), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g977 ( .A1(n_94), .A2(n_314), .B1(n_536), .B2(n_978), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_96), .A2(n_139), .B1(n_464), .B2(n_468), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_98), .A2(n_246), .B1(n_523), .B2(n_526), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_100), .A2(n_327), .B1(n_656), .B2(n_731), .Y(n_780) );
AO22x2_ASAP7_75t_L g818 ( .A1(n_102), .A2(n_819), .B1(n_839), .B2(n_840), .Y(n_818) );
INVx1_ASAP7_75t_L g840 ( .A(n_102), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_104), .A2(n_371), .B1(n_588), .B2(n_678), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_105), .A2(n_383), .B1(n_535), .B2(n_587), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_106), .A2(n_347), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_109), .A2(n_145), .B1(n_442), .B2(n_682), .Y(n_917) );
OAI22x1_ASAP7_75t_L g846 ( .A1(n_110), .A2(n_847), .B1(n_848), .B2(n_863), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_110), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_111), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_112), .A2(n_265), .B1(n_488), .B2(n_574), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_113), .A2(n_283), .B1(n_758), .B2(n_798), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_115), .A2(n_191), .B1(n_576), .B2(n_985), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_117), .A2(n_348), .B1(n_517), .B2(n_520), .Y(n_516) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_119), .A2(n_301), .B1(n_417), .B2(n_418), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_120), .A2(n_237), .B1(n_459), .B2(n_715), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_122), .A2(n_209), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_123), .A2(n_349), .B1(n_526), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_124), .A2(n_152), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_125), .A2(n_218), .B1(n_1004), .B2(n_1023), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_127), .A2(n_392), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_129), .A2(n_181), .B1(n_414), .B2(n_430), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_130), .A2(n_364), .B1(n_471), .B2(n_789), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_131), .A2(n_153), .B1(n_510), .B2(n_512), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_132), .A2(n_281), .B1(n_497), .B2(n_635), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_133), .A2(n_161), .B1(n_685), .B2(n_832), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_134), .A2(n_173), .B1(n_656), .B2(n_731), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_135), .A2(n_362), .B1(n_747), .B2(n_748), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_136), .A2(n_151), .B1(n_526), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_138), .A2(n_244), .B1(n_519), .B2(n_901), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_140), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g649 ( .A(n_142), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_143), .A2(n_217), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_144), .A2(n_156), .B1(n_587), .B2(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_147), .A2(n_329), .B1(n_414), .B2(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_148), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_149), .A2(n_312), .B1(n_474), .B2(n_475), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_150), .A2(n_378), .B1(n_681), .B2(n_682), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_154), .A2(n_330), .B1(n_475), .B2(n_668), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_155), .A2(n_188), .B1(n_526), .B2(n_1084), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_157), .Y(n_440) );
AO22x1_ASAP7_75t_L g554 ( .A1(n_158), .A2(n_229), .B1(n_536), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_159), .A2(n_178), .B1(n_798), .B2(n_961), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_160), .B(n_529), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_162), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_164), .A2(n_238), .B1(n_477), .B2(n_478), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_165), .A2(n_184), .B1(n_789), .B2(n_790), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_166), .Y(n_1068) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_167), .A2(n_370), .B1(n_656), .B2(n_731), .Y(n_730) );
OA22x2_ASAP7_75t_L g914 ( .A1(n_168), .A2(n_915), .B1(n_929), .B2(n_930), .Y(n_914) );
INVx1_ASAP7_75t_L g929 ( .A(n_168), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_169), .A2(n_306), .B1(n_696), .B2(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_171), .A2(n_270), .B1(n_632), .B2(n_752), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_172), .A2(n_376), .B1(n_442), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_174), .A2(n_211), .B1(n_622), .B2(n_623), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_175), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_176), .A2(n_252), .B1(n_695), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_177), .A2(n_221), .B1(n_632), .B2(n_692), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_179), .A2(n_302), .B1(n_571), .B2(n_809), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_180), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_182), .B(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_183), .A2(n_365), .B1(n_470), .B2(n_471), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_185), .A2(n_226), .B1(n_477), .B2(n_478), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_186), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_187), .A2(n_245), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_189), .A2(n_256), .B1(n_752), .B2(n_809), .Y(n_1001) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_192), .B(n_529), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_193), .A2(n_258), .B1(n_574), .B2(n_740), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_194), .A2(n_243), .B1(n_520), .B2(n_523), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_198), .A2(n_343), .B1(n_873), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_199), .A2(n_305), .B1(n_533), .B2(n_678), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_200), .A2(n_284), .B1(n_470), .B2(n_527), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_201), .A2(n_253), .B1(n_632), .B2(n_1020), .Y(n_1059) );
INVx1_ASAP7_75t_L g1041 ( .A(n_203), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_204), .A2(n_280), .B1(n_459), .B2(n_715), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_205), .A2(n_273), .B1(n_517), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_206), .A2(n_374), .B1(n_474), .B2(n_475), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_207), .A2(n_249), .B1(n_571), .B2(n_1081), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_208), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_210), .A2(n_235), .B1(n_638), .B2(n_1023), .Y(n_1085) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_212), .A2(n_387), .B1(n_567), .B2(n_568), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_213), .A2(n_321), .B1(n_478), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_214), .A2(n_388), .B1(n_568), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_215), .A2(n_380), .B1(n_636), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_216), .A2(n_255), .B1(n_475), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_219), .A2(n_393), .B1(n_615), .B2(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_220), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_222), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_223), .A2(n_389), .B1(n_414), .B2(n_430), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_224), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_228), .A2(n_397), .B1(n_598), .B2(n_869), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_230), .A2(n_261), .B1(n_492), .B2(n_498), .Y(n_1082) );
INVx2_ASAP7_75t_L g1096 ( .A(n_231), .Y(n_1096) );
XOR2x2_ASAP7_75t_L g957 ( .A(n_232), .B(n_958), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_233), .A2(n_250), .B1(n_747), .B2(n_748), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_234), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g1046 ( .A1(n_236), .A2(n_1047), .B1(n_1060), .B2(n_1061), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_236), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_239), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_240), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_241), .A2(n_266), .B1(n_470), .B2(n_471), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_242), .A2(n_248), .B1(n_532), .B2(n_645), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_247), .A2(n_335), .B1(n_603), .B2(n_752), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_251), .A2(n_345), .B1(n_459), .B2(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_257), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_269), .A2(n_279), .B1(n_689), .B2(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_274), .B(n_795), .Y(n_1075) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_275), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_277), .B(n_795), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_286), .A2(n_336), .B1(n_532), .B2(n_644), .Y(n_963) );
OA22x2_ASAP7_75t_L g864 ( .A1(n_287), .A2(n_865), .B1(n_866), .B2(n_881), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_287), .Y(n_865) );
AO21x2_ASAP7_75t_L g884 ( .A1(n_287), .A2(n_866), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g814 ( .A(n_288), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_289), .B(n_773), .Y(n_772) );
AOI22x1_ASAP7_75t_L g932 ( .A1(n_291), .A2(n_933), .B1(n_946), .B2(n_947), .Y(n_932) );
INVx1_ASAP7_75t_L g947 ( .A(n_291), .Y(n_947) );
XNOR2x1_ASAP7_75t_L g993 ( .A(n_293), .B(n_994), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_297), .A2(n_303), .B1(n_505), .B2(n_510), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_298), .A2(n_354), .B1(n_638), .B2(n_1020), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_299), .B(n_795), .Y(n_1050) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_301), .B(n_1040), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_304), .A2(n_326), .B1(n_464), .B2(n_471), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_307), .B(n_585), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_308), .A2(n_381), .B1(n_656), .B2(n_657), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_311), .A2(n_351), .B1(n_695), .B2(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_316), .A2(n_390), .B1(n_567), .B2(n_568), .Y(n_858) );
OA22x2_ASAP7_75t_L g408 ( .A1(n_317), .A2(n_409), .B1(n_410), .B2(n_480), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_317), .Y(n_409) );
AND2x2_ASAP7_75t_L g551 ( .A(n_318), .B(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_319), .A2(n_334), .B1(n_689), .B2(n_926), .Y(n_925) );
INVx3_ASAP7_75t_L g417 ( .A(n_320), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_322), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_323), .A2(n_359), .B1(n_587), .B2(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_325), .A2(n_340), .B1(n_797), .B2(n_833), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_328), .A2(n_339), .B1(n_536), .B2(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_332), .A2(n_382), .B1(n_503), .B2(n_803), .Y(n_877) );
INVx1_ASAP7_75t_L g546 ( .A(n_333), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_341), .Y(n_624) );
AND2x2_ASAP7_75t_L g894 ( .A(n_342), .B(n_895), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_350), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_353), .A2(n_361), .B1(n_492), .B2(n_807), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_355), .A2(n_360), .B1(n_689), .B2(n_903), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_366), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_367), .B(n_675), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_369), .A2(n_377), .B1(n_622), .B2(n_1052), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_372), .B(n_764), .Y(n_962) );
INVx1_ASAP7_75t_L g1036 ( .A(n_373), .Y(n_1036) );
NAND2xp5_ASAP7_75t_SL g1095 ( .A(n_373), .B(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1037 ( .A(n_375), .Y(n_1037) );
AND2x2_ASAP7_75t_R g1063 ( .A(n_375), .B(n_1036), .Y(n_1063) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_379), .Y(n_1094) );
XNOR2xp5_ASAP7_75t_L g743 ( .A(n_384), .B(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_385), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g1078 ( .A(n_386), .B(n_1052), .Y(n_1078) );
XOR2x2_ASAP7_75t_L g670 ( .A(n_395), .B(n_671), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_1043), .B(n_1044), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_842), .B(n_1033), .Y(n_399) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_400), .B(n_842), .Y(n_1043) );
XOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_703), .Y(n_400) );
OAI22xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_403), .B1(n_625), .B2(n_701), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_542), .B2(n_543), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
AO22x2_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_481), .B1(n_538), .B2(n_541), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g540 ( .A(n_408), .Y(n_540) );
AO22x2_ASAP7_75t_L g1013 ( .A1(n_408), .A2(n_540), .B1(n_992), .B2(n_993), .Y(n_1013) );
INVx1_ASAP7_75t_L g480 ( .A(n_410), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_461), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_439), .C(n_451), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_433), .Y(n_412) );
INVx1_ASAP7_75t_SL g880 ( .A(n_414), .Y(n_880) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_422), .Y(n_414) );
AND2x2_ASAP7_75t_L g454 ( .A(n_415), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g468 ( .A(n_415), .B(n_467), .Y(n_468) );
AND2x4_ASAP7_75t_L g511 ( .A(n_415), .B(n_455), .Y(n_511) );
AND2x2_ASAP7_75t_L g534 ( .A(n_415), .B(n_422), .Y(n_534) );
AND2x2_ASAP7_75t_L g715 ( .A(n_415), .B(n_455), .Y(n_715) );
AND2x2_ASAP7_75t_L g790 ( .A(n_415), .B(n_467), .Y(n_790) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
AND2x2_ASAP7_75t_L g432 ( .A(n_416), .B(n_420), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_416), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
INVx2_ASAP7_75t_L g418 ( .A(n_417), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
OAI22x1_ASAP7_75t_L g423 ( .A1(n_417), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_417), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_417), .Y(n_429) );
AND2x4_ASAP7_75t_L g437 ( .A(n_419), .B(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_420), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g443 ( .A(n_422), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g474 ( .A(n_422), .B(n_437), .Y(n_474) );
AND2x4_ASAP7_75t_L g525 ( .A(n_422), .B(n_437), .Y(n_525) );
AND2x4_ASAP7_75t_L g656 ( .A(n_422), .B(n_444), .Y(n_656) );
AND2x2_ASAP7_75t_L g668 ( .A(n_422), .B(n_437), .Y(n_668) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_423), .Y(n_431) );
AND2x2_ASAP7_75t_L g436 ( .A(n_423), .B(n_428), .Y(n_436) );
INVx2_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
AND2x4_ASAP7_75t_L g467 ( .A(n_427), .B(n_456), .Y(n_467) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g455 ( .A(n_428), .B(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g479 ( .A(n_428), .Y(n_479) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g537 ( .A(n_431), .B(n_432), .Y(n_537) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_431), .B(n_432), .Y(n_728) );
AND2x4_ASAP7_75t_L g475 ( .A(n_432), .B(n_467), .Y(n_475) );
AND2x4_ASAP7_75t_L g478 ( .A(n_432), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g498 ( .A(n_432), .B(n_479), .Y(n_498) );
AND2x4_ASAP7_75t_L g521 ( .A(n_432), .B(n_467), .Y(n_521) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g776 ( .A(n_435), .Y(n_776) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AND2x4_ASAP7_75t_L g448 ( .A(n_436), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g459 ( .A(n_436), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g514 ( .A(n_436), .B(n_460), .Y(n_514) );
AND2x2_ASAP7_75t_L g531 ( .A(n_436), .B(n_437), .Y(n_531) );
AND2x2_ASAP7_75t_L g657 ( .A(n_436), .B(n_449), .Y(n_657) );
AND2x2_ASAP7_75t_L g660 ( .A(n_436), .B(n_460), .Y(n_660) );
AND2x2_ASAP7_75t_L g731 ( .A(n_436), .B(n_449), .Y(n_731) );
AND2x4_ASAP7_75t_L g466 ( .A(n_437), .B(n_467), .Y(n_466) );
AND2x6_ASAP7_75t_L g470 ( .A(n_437), .B(n_455), .Y(n_470) );
AND2x2_ASAP7_75t_L g487 ( .A(n_437), .B(n_455), .Y(n_487) );
AND2x2_ASAP7_75t_L g789 ( .A(n_437), .B(n_467), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_446), .B2(n_447), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_SL g758 ( .A(n_442), .Y(n_758) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_443), .Y(n_802) );
AND2x6_ASAP7_75t_L g471 ( .A(n_444), .B(n_467), .Y(n_471) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_444), .B(n_455), .Y(n_477) );
AND2x4_ASAP7_75t_L g490 ( .A(n_444), .B(n_467), .Y(n_490) );
AND2x2_ASAP7_75t_L g496 ( .A(n_444), .B(n_455), .Y(n_496) );
AND2x2_ASAP7_75t_L g664 ( .A(n_444), .B(n_455), .Y(n_664) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
INVx2_ASAP7_75t_SL g620 ( .A(n_447), .Y(n_620) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
BUFx6f_ASAP7_75t_SL g682 ( .A(n_448), .Y(n_682) );
BUFx3_ASAP7_75t_L g803 ( .A(n_448), .Y(n_803) );
BUFx4f_ASAP7_75t_L g855 ( .A(n_448), .Y(n_855) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_457), .B2(n_458), .Y(n_451) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_469), .Y(n_462) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
INVx2_ASAP7_75t_SL g615 ( .A(n_465), .Y(n_615) );
INVx2_ASAP7_75t_L g638 ( .A(n_465), .Y(n_638) );
INVx3_ASAP7_75t_SL g751 ( .A(n_465), .Y(n_751) );
INVx2_ASAP7_75t_SL g837 ( .A(n_465), .Y(n_837) );
INVx8_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_468), .Y(n_527) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_468), .Y(n_699) );
INVx2_ASAP7_75t_L g741 ( .A(n_468), .Y(n_741) );
BUFx3_ASAP7_75t_L g827 ( .A(n_468), .Y(n_827) );
INVx1_ASAP7_75t_L g924 ( .A(n_470), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
NAND4xp75_ASAP7_75t_L g482 ( .A(n_483), .B(n_499), .C(n_515), .D(n_528), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_491), .Y(n_483) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g574 ( .A(n_486), .Y(n_574) );
INVx2_ASAP7_75t_L g604 ( .A(n_486), .Y(n_604) );
INVx2_ASAP7_75t_L g691 ( .A(n_486), .Y(n_691) );
INVx3_ASAP7_75t_L g809 ( .A(n_486), .Y(n_809) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g632 ( .A(n_487), .Y(n_632) );
BUFx2_ASAP7_75t_L g754 ( .A(n_487), .Y(n_754) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_489), .A2(n_601), .B1(n_602), .B2(n_605), .Y(n_600) );
INVx2_ASAP7_75t_L g633 ( .A(n_489), .Y(n_633) );
INVx2_ASAP7_75t_L g692 ( .A(n_489), .Y(n_692) );
INVx2_ASAP7_75t_L g752 ( .A(n_489), .Y(n_752) );
INVx2_ASAP7_75t_SL g810 ( .A(n_489), .Y(n_810) );
INVx1_ASAP7_75t_SL g861 ( .A(n_489), .Y(n_861) );
INVx2_ASAP7_75t_SL g991 ( .A(n_489), .Y(n_991) );
INVx8_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_494), .Y(n_987) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g636 ( .A(n_495), .Y(n_636) );
INVx1_ASAP7_75t_L g926 ( .A(n_495), .Y(n_926) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_496), .Y(n_598) );
BUFx3_ASAP7_75t_L g806 ( .A(n_496), .Y(n_806) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx5_ASAP7_75t_SL g569 ( .A(n_498), .Y(n_569) );
BUFx2_ASAP7_75t_L g689 ( .A(n_498), .Y(n_689) );
BUFx3_ASAP7_75t_L g807 ( .A(n_498), .Y(n_807) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_502), .A2(n_506), .B1(n_558), .B2(n_559), .Y(n_557) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g681 ( .A(n_504), .Y(n_681) );
INVx1_ASAP7_75t_L g1074 ( .A(n_504), .Y(n_1074) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g759 ( .A(n_507), .Y(n_759) );
BUFx4f_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g562 ( .A(n_510), .Y(n_562) );
BUFx2_ASAP7_75t_L g622 ( .A(n_510), .Y(n_622) );
BUFx2_ASAP7_75t_L g961 ( .A(n_510), .Y(n_961) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g684 ( .A(n_511), .Y(n_684) );
BUFx2_ASAP7_75t_L g797 ( .A(n_511), .Y(n_797) );
BUFx3_ASAP7_75t_L g832 ( .A(n_511), .Y(n_832) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_513), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g623 ( .A(n_513), .Y(n_623) );
INVx2_ASAP7_75t_L g685 ( .A(n_513), .Y(n_685) );
INVx2_ASAP7_75t_SL g766 ( .A(n_513), .Y(n_766) );
INVx2_ASAP7_75t_L g798 ( .A(n_513), .Y(n_798) );
INVx2_ASAP7_75t_SL g833 ( .A(n_513), .Y(n_833) );
INVx6_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_519), .Y(n_860) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_SL g576 ( .A(n_521), .Y(n_576) );
INVx2_ASAP7_75t_L g697 ( .A(n_521), .Y(n_697) );
BUFx3_ASAP7_75t_L g748 ( .A(n_521), .Y(n_748) );
BUFx3_ASAP7_75t_L g812 ( .A(n_521), .Y(n_812) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_524), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g640 ( .A(n_524), .Y(n_640) );
INVx2_ASAP7_75t_L g747 ( .A(n_524), .Y(n_747) );
INVx2_ASAP7_75t_L g985 ( .A(n_524), .Y(n_985) );
INVx3_ASAP7_75t_L g1004 ( .A(n_524), .Y(n_1004) );
INVx6_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g695 ( .A(n_525), .Y(n_695) );
BUFx3_ASAP7_75t_L g1084 ( .A(n_525), .Y(n_1084) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g617 ( .A(n_527), .Y(n_617) );
BUFx2_ASAP7_75t_L g764 ( .A(n_529), .Y(n_764) );
INVx4_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g553 ( .A(n_530), .Y(n_553) );
INVx3_ASAP7_75t_SL g585 ( .A(n_530), .Y(n_585) );
INVx4_ASAP7_75t_SL g675 ( .A(n_530), .Y(n_675) );
INVx3_ASAP7_75t_L g795 ( .A(n_530), .Y(n_795) );
INVx3_ASAP7_75t_L g896 ( .A(n_530), .Y(n_896) );
INVx6_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g556 ( .A(n_534), .Y(n_556) );
BUFx3_ASAP7_75t_L g588 ( .A(n_534), .Y(n_588) );
BUFx5_ASAP7_75t_L g978 ( .A(n_534), .Y(n_978) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g592 ( .A(n_536), .Y(n_592) );
BUFx12f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g646 ( .A(n_537), .Y(n_646) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_578), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_577), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_546), .B(n_549), .Y(n_577) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_564), .Y(n_549) );
NOR4xp75_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .C(n_557), .D(n_560), .Y(n_550) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g762 ( .A(n_556), .Y(n_762) );
INVx2_ASAP7_75t_L g853 ( .A(n_556), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_572), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_569), .A2(n_595), .B1(n_596), .B2(n_599), .Y(n_594) );
INVx2_ASAP7_75t_L g869 ( .A(n_569), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g610 ( .A(n_576), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_624), .Y(n_578) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_580), .B(n_593), .C(n_606), .D(n_618), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_586), .B2(n_589), .C(n_590), .Y(n_581) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g822 ( .A(n_585), .Y(n_822) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_616), .B2(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g901 ( .A(n_617), .Y(n_901) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
BUFx2_ASAP7_75t_L g702 ( .A(n_625), .Y(n_702) );
OA22x2_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_650), .B1(n_651), .B2(n_700), .Y(n_625) );
INVx1_ASAP7_75t_L g700 ( .A(n_626), .Y(n_700) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_649), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_641), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .C(n_637), .D(n_639), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .C(n_647), .D(n_648), .Y(n_641) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g678 ( .A(n_646), .Y(n_678) );
INVx2_ASAP7_75t_L g800 ( .A(n_646), .Y(n_800) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
XNOR2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_670), .Y(n_651) );
XNOR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_669), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_662), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_658), .C(n_659), .D(n_661), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .C(n_666), .D(n_667), .Y(n_662) );
NAND2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_686), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_679), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_676), .B(n_677), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g975 ( .A1(n_674), .A2(n_976), .B(n_977), .Y(n_975) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
BUFx2_ASAP7_75t_SL g909 ( .A(n_682), .Y(n_909) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_693), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .Y(n_693) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_699), .Y(n_755) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_768), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OA22x2_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_743), .B2(n_767), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
XNOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_722), .Y(n_707) );
XNOR2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_717), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .C(n_714), .D(n_716), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .C(n_720), .D(n_721), .Y(n_717) );
AO22x2_ASAP7_75t_L g770 ( .A1(n_722), .A2(n_771), .B1(n_815), .B2(n_816), .Y(n_770) );
INVx1_ASAP7_75t_L g815 ( .A(n_722), .Y(n_815) );
XOR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_742), .Y(n_722) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_733), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_729), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g873 ( .A(n_741), .Y(n_873) );
INVx2_ASAP7_75t_SL g767 ( .A(n_743), .Y(n_767) );
NOR2xp67_ASAP7_75t_L g744 ( .A(n_745), .B(n_756), .Y(n_744) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .C(n_750), .D(n_753), .Y(n_745) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_754), .Y(n_1081) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .C(n_763), .D(n_765), .Y(n_756) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_817), .B2(n_841), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g816 ( .A(n_771), .Y(n_816) );
XOR2x1_ASAP7_75t_SL g771 ( .A(n_772), .B(n_791), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_774), .B(n_782), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
OAI21xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_777), .B(n_778), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_786), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
XNOR2x1_ASAP7_75t_L g791 ( .A(n_792), .B(n_814), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_804), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .C(n_799), .D(n_801), .Y(n_793) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_800), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_802), .Y(n_908) );
BUFx6f_ASAP7_75t_SL g1052 ( .A(n_803), .Y(n_1052) );
NAND4xp25_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .C(n_811), .D(n_813), .Y(n_804) );
BUFx2_ASAP7_75t_L g903 ( .A(n_806), .Y(n_903) );
BUFx6f_ASAP7_75t_L g1023 ( .A(n_812), .Y(n_1023) );
INVx1_ASAP7_75t_L g841 ( .A(n_817), .Y(n_841) );
INVx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_SL g839 ( .A(n_819), .Y(n_839) );
AND2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_829), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_825), .Y(n_820) );
OAI21xp33_ASAP7_75t_SL g821 ( .A1(n_822), .A2(n_823), .B(n_824), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_835), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_838), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_952), .B1(n_1031), .B2(n_1032), .Y(n_842) );
INVx1_ASAP7_75t_L g1031 ( .A(n_843), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_887), .B2(n_888), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
OA22x2_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_864), .B1(n_882), .B2(n_883), .Y(n_845) );
INVx1_ASAP7_75t_SL g882 ( .A(n_846), .Y(n_882) );
INVx2_ASAP7_75t_SL g863 ( .A(n_848), .Y(n_863) );
OR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_856), .Y(n_848) );
NAND4xp25_ASAP7_75t_SL g849 ( .A(n_850), .B(n_851), .C(n_852), .D(n_854), .Y(n_849) );
NAND4xp25_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .C(n_859), .D(n_862), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_865), .Y(n_886) );
INVx1_ASAP7_75t_L g881 ( .A(n_866), .Y(n_881) );
NOR2x1_ASAP7_75t_SL g885 ( .A(n_866), .B(n_886), .Y(n_885) );
NAND4xp75_ASAP7_75t_L g866 ( .A(n_867), .B(n_871), .C(n_875), .D(n_878), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_870), .Y(n_867) );
AND2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_874), .Y(n_871) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_873), .Y(n_1020) );
AND2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AO22x2_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_913), .B1(n_950), .B2(n_951), .Y(n_889) );
INVx1_ASAP7_75t_L g950 ( .A(n_890), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_891), .B(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_905), .Y(n_892) );
NOR3xp33_ASAP7_75t_SL g893 ( .A(n_894), .B(n_897), .C(n_898), .Y(n_893) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND4xp25_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .C(n_902), .D(n_904), .Y(n_898) );
AND2x2_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g951 ( .A(n_913), .Y(n_951) );
AOI22x1_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_931), .B1(n_948), .B2(n_949), .Y(n_913) );
INVx2_ASAP7_75t_L g949 ( .A(n_914), .Y(n_949) );
INVx1_ASAP7_75t_L g930 ( .A(n_915), .Y(n_930) );
NOR2x1_ASAP7_75t_L g915 ( .A(n_916), .B(n_921), .Y(n_915) );
NAND4xp25_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .C(n_919), .D(n_920), .Y(n_916) );
NAND4xp25_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_927), .D(n_928), .Y(n_921) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_SL g948 ( .A(n_931), .Y(n_948) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g946 ( .A(n_933), .Y(n_946) );
NAND2x1_ASAP7_75t_SL g933 ( .A(n_934), .B(n_939), .Y(n_933) );
NOR2xp67_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
NOR2x1_ASAP7_75t_L g939 ( .A(n_940), .B(n_943), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_953), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_1010), .B2(n_1011), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_970), .B1(n_971), .B2(n_1009), .Y(n_956) );
INVx5_ASAP7_75t_L g1009 ( .A(n_957), .Y(n_1009) );
NOR2x1_ASAP7_75t_L g958 ( .A(n_959), .B(n_965), .Y(n_958) );
NAND4xp25_ASAP7_75t_L g959 ( .A(n_960), .B(n_962), .C(n_963), .D(n_964), .Y(n_959) );
NAND4xp25_ASAP7_75t_L g965 ( .A(n_966), .B(n_967), .C(n_968), .D(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_992), .B1(n_993), .B2(n_1006), .Y(n_971) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_973), .Y(n_1007) );
AND2x2_ASAP7_75t_L g973 ( .A(n_974), .B(n_982), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_979), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_983), .B(n_988), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_986), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_990), .Y(n_988) );
INVx1_ASAP7_75t_SL g992 ( .A(n_993), .Y(n_992) );
OR2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_1000), .Y(n_994) );
NAND4xp25_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .C(n_998), .D(n_999), .Y(n_995) );
NAND4xp25_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .C(n_1003), .D(n_1005), .Y(n_1000) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
OA22x2_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
XNOR2x1_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1030), .Y(n_1015) );
NOR2xp67_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1024), .Y(n_1016) );
NAND4xp25_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .C(n_1021), .D(n_1022), .Y(n_1017) );
NAND4xp25_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1026), .C(n_1028), .D(n_1029), .Y(n_1024) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1035), .B(n_1039), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1037), .Y(n_1092) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
NAND2xp5_ASAP7_75t_SL g1044 ( .A(n_1045), .B(n_1097), .Y(n_1044) );
OA222x2_ASAP7_75t_SL g1045 ( .A1(n_1046), .A2(n_1062), .B1(n_1064), .B2(n_1068), .C1(n_1086), .C2(n_1089), .Y(n_1045) );
CKINVDCx16_ASAP7_75t_R g1061 ( .A(n_1047), .Y(n_1061) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
NOR2x1_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1055), .Y(n_1048) );
NAND4xp25_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .C(n_1053), .D(n_1054), .Y(n_1049) );
NAND4xp25_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .C(n_1058), .D(n_1059), .Y(n_1055) );
INVx1_ASAP7_75t_SL g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
XNOR2x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1079), .Y(n_1069) );
NAND4xp25_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1076), .C(n_1077), .D(n_1078), .Y(n_1070) );
OA21x2_ASAP7_75t_SL g1071 ( .A1(n_1072), .A2(n_1073), .B(n_1075), .Y(n_1071) );
INVxp33_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NAND4xp25_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .C(n_1083), .D(n_1085), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1086 ( .A(n_1087), .Y(n_1086) );
CKINVDCx6p67_ASAP7_75t_R g1087 ( .A(n_1088), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_1090), .Y(n_1089) );
CKINVDCx20_ASAP7_75t_R g1090 ( .A(n_1091), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1092), .Y(n_1101) );
AND2x4_ASAP7_75t_SL g1100 ( .A(n_1093), .B(n_1101), .Y(n_1100) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_1100), .Y(n_1099) );
endmodule