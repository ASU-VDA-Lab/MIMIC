module fake_netlist_5_1869_n_763 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_763);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_763;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_142;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_144;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_35),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_53),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_20),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_2),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_57),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_9),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_32),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_78),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_3),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_81),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_L g166 ( 
.A(n_60),
.B(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_42),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_74),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_75),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_94),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_0),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_55),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_130),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_46),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_2),
.Y(n_209)
);

OAI22x1_ASAP7_75t_R g210 ( 
.A1(n_159),
.A2(n_163),
.B1(n_184),
.B2(n_164),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_3),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_14),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_15),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_149),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_150),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_194),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_216),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_206),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_153),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_191),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_205),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_205),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_190),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_210),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_211),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_211),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_234),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_262),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_209),
.B1(n_222),
.B2(n_225),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_206),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_222),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_206),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_206),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_223),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_215),
.C(n_209),
.Y(n_300)
);

AND2x4_ASAP7_75t_SL g301 ( 
.A(n_240),
.B(n_225),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_219),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_269),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_229),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_217),
.C(n_212),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_269),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_237),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_239),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_241),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_203),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_203),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_203),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_213),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

BUFx6f_ASAP7_75t_SL g326 ( 
.A(n_277),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_242),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_245),
.B(n_229),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_229),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_247),
.B(n_219),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_249),
.B(n_229),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_213),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_250),
.B(n_199),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_267),
.B(n_229),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_275),
.B(n_219),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_235),
.B(n_219),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_213),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_236),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_253),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_266),
.B(n_219),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_255),
.B(n_201),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_246),
.A2(n_202),
.B1(n_208),
.B2(n_204),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_255),
.B(n_201),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_333),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_289),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_201),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_303),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_220),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_196),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_220),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_284),
.B(n_154),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_220),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_334),
.B(n_158),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_208),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_305),
.B(n_162),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_165),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

BUFx6f_ASAP7_75t_SL g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_300),
.B(n_283),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_220),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_338),
.A2(n_202),
.B1(n_188),
.B2(n_185),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_292),
.B(n_175),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_319),
.B(n_178),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_292),
.B(n_179),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_299),
.B(n_7),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_180),
.Y(n_388)
);

OR2x6_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_7),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_181),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_291),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_309),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_310),
.B(n_183),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_293),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_294),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_8),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_295),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_292),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_302),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_331),
.B(n_16),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_338),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_292),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_292),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_306),
.B(n_17),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_336),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_288),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_349),
.A2(n_335),
.B(n_344),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_SL g417 ( 
.A(n_377),
.B(n_304),
.C(n_298),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_329),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_L g419 ( 
.A1(n_346),
.A2(n_296),
.B1(n_342),
.B2(n_330),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_361),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_8),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_346),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_18),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_19),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_349),
.A2(n_370),
.B(n_365),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_326),
.B1(n_86),
.B2(n_87),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_352),
.A2(n_84),
.B(n_139),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_408),
.B(n_21),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_380),
.B1(n_390),
.B2(n_391),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_375),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_408),
.B(n_395),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_326),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_389),
.A2(n_12),
.B1(n_13),
.B2(n_23),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_13),
.Y(n_439)
);

CKINVDCx8_ASAP7_75t_R g440 ( 
.A(n_389),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_24),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_352),
.A2(n_25),
.B(n_26),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_386),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_351),
.B(n_33),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_34),
.B(n_36),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_358),
.B(n_37),
.Y(n_447)
);

O2A1O1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_362),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_41),
.Y(n_449)
);

AO32x1_ASAP7_75t_L g450 ( 
.A1(n_401),
.A2(n_43),
.A3(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_365),
.B(n_48),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_379),
.A2(n_49),
.B(n_50),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_382),
.A2(n_51),
.B(n_52),
.C(n_54),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_367),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_410),
.A2(n_411),
.B(n_405),
.Y(n_459)
);

AO32x1_ASAP7_75t_L g460 ( 
.A1(n_402),
.A2(n_61),
.A3(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_388),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_SL g463 ( 
.A(n_368),
.B(n_73),
.C(n_76),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_383),
.A2(n_77),
.B(n_80),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_392),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_466)
);

O2A1O1Ixp5_ASAP7_75t_L g467 ( 
.A1(n_383),
.A2(n_90),
.B(n_92),
.C(n_93),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_398),
.A2(n_95),
.B(n_97),
.C(n_98),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_363),
.B(n_99),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_415),
.A2(n_385),
.B(n_412),
.Y(n_471)
);

AO21x2_ASAP7_75t_L g472 ( 
.A1(n_426),
.A2(n_385),
.B(n_407),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_404),
.B(n_403),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_413),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_434),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_428),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_347),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_435),
.B(n_384),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_434),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g482 ( 
.A1(n_451),
.A2(n_355),
.B(n_371),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_419),
.A2(n_354),
.B(n_373),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_437),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_440),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_441),
.A2(n_347),
.B(n_373),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_418),
.B(n_369),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_447),
.A2(n_406),
.B(n_348),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_467),
.A2(n_406),
.B(n_348),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_406),
.B(n_348),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_100),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_101),
.B(n_102),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_429),
.A2(n_103),
.B(n_105),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

BUFx2_ASAP7_75t_R g500 ( 
.A(n_430),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

NAND2x1_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_106),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_469),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_107),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_469),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_456),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_449),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_493),
.A2(n_495),
.B(n_490),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_494),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_494),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_476),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_486),
.Y(n_523)
);

BUFx2_ASAP7_75t_R g524 ( 
.A(n_488),
.Y(n_524)
);

CKINVDCx11_ASAP7_75t_R g525 ( 
.A(n_476),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_493),
.A2(n_442),
.B(n_452),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_445),
.B(n_425),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_414),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_516),
.A2(n_438),
.B1(n_427),
.B2(n_374),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_475),
.B(n_443),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_489),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_501),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_485),
.B(n_417),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_510),
.A2(n_423),
.B(n_461),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_501),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_514),
.A2(n_453),
.B(n_448),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_503),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_514),
.A2(n_468),
.B(n_466),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_516),
.A2(n_374),
.B1(n_432),
.B2(n_460),
.Y(n_544)
);

AOI222xp33_ASAP7_75t_L g545 ( 
.A1(n_479),
.A2(n_460),
.B1(n_111),
.B2(n_115),
.C1(n_116),
.C2(n_118),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_505),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_508),
.Y(n_547)
);

CKINVDCx11_ASAP7_75t_R g548 ( 
.A(n_511),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_504),
.Y(n_549)
);

CKINVDCx11_ASAP7_75t_R g550 ( 
.A(n_511),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_110),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_491),
.Y(n_552)
);

BUFx8_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_483),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_483),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_474),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_548),
.Y(n_560)
);

AO31x2_ASAP7_75t_L g561 ( 
.A1(n_536),
.A2(n_509),
.A3(n_515),
.B(n_512),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_R g562 ( 
.A(n_557),
.B(n_488),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_SL g563 ( 
.A(n_544),
.B(n_487),
.C(n_500),
.Y(n_563)
);

AND2x4_ASAP7_75t_SL g564 ( 
.A(n_535),
.B(n_480),
.Y(n_564)
);

NAND2x1_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_502),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_534),
.B(n_485),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_R g567 ( 
.A(n_534),
.B(n_487),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_531),
.B(n_504),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_508),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_554),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_529),
.A2(n_496),
.B1(n_506),
.B2(n_482),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_513),
.Y(n_572)
);

INVx8_ASAP7_75t_L g573 ( 
.A(n_555),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_508),
.Y(n_574)
);

AO31x2_ASAP7_75t_L g575 ( 
.A1(n_520),
.A2(n_515),
.A3(n_509),
.B(n_471),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_540),
.B(n_513),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_556),
.B(n_499),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_541),
.B(n_496),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_499),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_504),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_539),
.B(n_496),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_553),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_R g583 ( 
.A(n_550),
.B(n_489),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_553),
.B(n_489),
.Y(n_584)
);

AO31x2_ASAP7_75t_L g585 ( 
.A1(n_521),
.A2(n_532),
.A3(n_533),
.B(n_537),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_535),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_529),
.A2(n_506),
.B1(n_502),
.B2(n_484),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_523),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_R g589 ( 
.A(n_551),
.B(n_502),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_540),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_549),
.B(n_482),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_530),
.A2(n_484),
.B1(n_473),
.B2(n_482),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_518),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_SL g596 ( 
.A(n_519),
.B(n_497),
.C(n_498),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_522),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

OAI222xp33_ASAP7_75t_L g599 ( 
.A1(n_522),
.A2(n_497),
.B1(n_498),
.B2(n_473),
.C1(n_484),
.C2(n_124),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_524),
.B(n_473),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_524),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_549),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_538),
.B(n_542),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_538),
.B(n_472),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_559),
.B(n_542),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_595),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_604),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_593),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_472),
.Y(n_609)
);

NAND2x1_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_547),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_591),
.A2(n_545),
.B1(n_555),
.B2(n_471),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_570),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_472),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_595),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_585),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_545),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_562),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_575),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_597),
.A2(n_471),
.B1(n_492),
.B2(n_555),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_575),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_561),
.B(n_517),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_566),
.A2(n_492),
.B1(n_526),
.B2(n_527),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_561),
.B(n_492),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_561),
.B(n_120),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_602),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_581),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_574),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_578),
.Y(n_630)
);

CKINVDCx11_ASAP7_75t_R g631 ( 
.A(n_601),
.Y(n_631)
);

NOR2x1_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_121),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_577),
.B(n_122),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_594),
.B(n_138),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_574),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_569),
.B(n_123),
.Y(n_637)
);

INVx8_ASAP7_75t_L g638 ( 
.A(n_573),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_566),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_579),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_572),
.B(n_137),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_563),
.B(n_125),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_612),
.B(n_590),
.Y(n_643)
);

AND2x4_ASAP7_75t_SL g644 ( 
.A(n_640),
.B(n_558),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_606),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_615),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_587),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_611),
.B(n_571),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_605),
.B(n_576),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_618),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_607),
.B(n_576),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_639),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_609),
.B(n_558),
.Y(n_654)
);

OA21x2_ASAP7_75t_L g655 ( 
.A1(n_621),
.A2(n_599),
.B(n_596),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_618),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_628),
.B(n_598),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_616),
.B(n_568),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_639),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_621),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_629),
.B(n_583),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_622),
.Y(n_662)
);

AND2x4_ASAP7_75t_SL g663 ( 
.A(n_639),
.B(n_568),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_609),
.B(n_613),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_608),
.B(n_564),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_622),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_613),
.B(n_560),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_619),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_646),
.B(n_624),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_654),
.B(n_608),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_608),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_647),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_627),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_635),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_645),
.Y(n_676)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_643),
.B(n_626),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_R g678 ( 
.A(n_653),
.B(n_584),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_667),
.B(n_669),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_662),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_662),
.B(n_635),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_667),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_666),
.Y(n_683)
);

NAND2x1p5_ASAP7_75t_L g684 ( 
.A(n_655),
.B(n_610),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_648),
.B(n_624),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_644),
.B(n_639),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_676),
.B(n_648),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_674),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_685),
.B(n_670),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_672),
.B(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_682),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_673),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_677),
.B(n_632),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_680),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_684),
.A2(n_649),
.B(n_616),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_681),
.B(n_655),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_678),
.A2(n_649),
.B1(n_658),
.B2(n_589),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_692),
.Y(n_698)
);

OAI21xp33_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_658),
.B(n_670),
.Y(n_699)
);

AOI21xp33_ASAP7_75t_L g700 ( 
.A1(n_693),
.A2(n_567),
.B(n_657),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_687),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_691),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_688),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_698),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_702),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_699),
.Y(n_706)
);

AOI222xp33_ASAP7_75t_L g707 ( 
.A1(n_700),
.A2(n_642),
.B1(n_634),
.B2(n_631),
.C1(n_644),
.C2(n_689),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_697),
.B(n_617),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_704),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_SL g711 ( 
.A(n_707),
.B(n_657),
.C(n_650),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_709),
.B(n_705),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);

NAND2x1_ASAP7_75t_SL g714 ( 
.A(n_710),
.B(n_703),
.Y(n_714)
);

OAI221xp5_ASAP7_75t_L g715 ( 
.A1(n_714),
.A2(n_711),
.B1(n_696),
.B2(n_684),
.C(n_661),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_712),
.A2(n_696),
.B1(n_631),
.B2(n_686),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_713),
.B(n_582),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_712),
.A2(n_634),
.B(n_626),
.C(n_641),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_715),
.B(n_716),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_718),
.B(n_641),
.Y(n_720)
);

NOR2x1_ASAP7_75t_L g721 ( 
.A(n_717),
.B(n_633),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_717),
.B(n_694),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_717),
.A2(n_665),
.B1(n_683),
.B2(n_637),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_717),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_715),
.B(n_633),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_721),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_722),
.Y(n_728)
);

NAND5xp2_ASAP7_75t_L g729 ( 
.A(n_719),
.B(n_620),
.C(n_625),
.D(n_671),
.E(n_623),
.Y(n_729)
);

NOR2x1_ASAP7_75t_L g730 ( 
.A(n_725),
.B(n_637),
.Y(n_730)
);

AOI211x1_ASAP7_75t_L g731 ( 
.A1(n_720),
.A2(n_685),
.B(n_675),
.C(n_690),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_719),
.A2(n_655),
.B1(n_663),
.B2(n_659),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_R g733 ( 
.A(n_728),
.B(n_638),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_726),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_727),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_730),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_727),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_732),
.B(n_680),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_731),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_729),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_734),
.A2(n_580),
.B1(n_679),
.B2(n_637),
.Y(n_741)
);

XNOR2x1_ASAP7_75t_L g742 ( 
.A(n_737),
.B(n_129),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_735),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_736),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_739),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_738),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_740),
.A2(n_638),
.B1(n_580),
.B2(n_573),
.Y(n_747)
);

OAI31xp33_ASAP7_75t_SL g748 ( 
.A1(n_743),
.A2(n_733),
.A3(n_638),
.B(n_681),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_744),
.A2(n_638),
.B1(n_663),
.B2(n_630),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_630),
.B1(n_656),
.B2(n_651),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_746),
.A2(n_565),
.B1(n_651),
.B2(n_660),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_741),
.B(n_636),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_753),
.A2(n_747),
.B(n_660),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_752),
.Y(n_756)
);

XOR2xp5_ASAP7_75t_L g757 ( 
.A(n_754),
.B(n_749),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_756),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_756),
.Y(n_759)
);

NOR2x1_ASAP7_75t_L g760 ( 
.A(n_759),
.B(n_748),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_760),
.B(n_758),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_761),
.B(n_757),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_762),
.A2(n_755),
.B1(n_750),
.B2(n_636),
.Y(n_763)
);


endmodule