module real_jpeg_14656_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g103 ( 
.A(n_0),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_72),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_119),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_5),
.A2(n_62),
.B(n_65),
.C(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_87),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_45),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_5),
.A2(n_45),
.B(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_30),
.C(n_35),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_172),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_5),
.A2(n_106),
.B1(n_107),
.B2(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_48),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_10),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_175),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_175),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_164),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_164),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_14),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_121)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_91),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_77),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_20),
.A2(n_73),
.B1(n_308),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_20),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_58),
.B2(n_59),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_73),
.C(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_23),
.A2(n_24),
.B1(n_78),
.B2(n_79),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_40),
.C(n_58),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_33),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_25),
.A2(n_37),
.B(n_138),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_25),
.A2(n_127),
.B(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_26),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_26),
.B(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_26),
.A2(n_114),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_26),
.A2(n_113),
.B1(n_219),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_26),
.A2(n_113),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_26),
.A2(n_113),
.B1(n_240),
.B2(n_250),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_29),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_SL g225 ( 
.A(n_28),
.B(n_46),
.C(n_50),
.Y(n_225)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_29),
.A2(n_51),
.B(n_223),
.C(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_29),
.B(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_33),
.A2(n_112),
.B(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_33),
.B(n_172),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_34),
.B(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_35),
.B(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_38),
.B(n_113),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_54),
.B(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_48),
.B(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_44),
.A2(n_54),
.B(n_82),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_45),
.A2(n_63),
.B(n_172),
.Y(n_191)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_48),
.A2(n_53),
.B1(n_81),
.B2(n_125),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_49),
.A2(n_52),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_49),
.A2(n_54),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_49),
.A2(n_54),
.B1(n_178),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_49),
.A2(n_54),
.B1(n_198),
.B2(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_69),
.B2(n_71),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_71),
.B(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_60),
.A2(n_86),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_61),
.B1(n_118),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_60),
.A2(n_61),
.B1(n_163),
.B2(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_69),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_73),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_73),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_75),
.A2(n_87),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_77),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_83),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.CI(n_88),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_302),
.B(n_316),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_165),
.B(n_301),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_145),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_94),
.B(n_145),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_122),
.B2(n_144),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_95),
.B(n_123),
.C(n_131),
.Y(n_314)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_115),
.C(n_117),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_98),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_99),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_290)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_102),
.A2(n_106),
.B(n_255),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_103),
.A2(n_155),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_103),
.A2(n_105),
.B(n_188),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_103),
.A2(n_187),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_104),
.A2(n_157),
.B(n_187),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_107),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_106),
.A2(n_107),
.B1(n_253),
.B2(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_107),
.B(n_172),
.Y(n_259)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_129),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_117),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_131),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B(n_130),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_130),
.B(n_305),
.C(n_309),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_130),
.B(n_305),
.CI(n_309),
.CON(n_315),
.SN(n_315)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_132),
.A2(n_133),
.B(n_141),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_140),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_151),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.C(n_161),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_152),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_158),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_292)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_295),
.B(n_300),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_208),
.B(n_286),
.C(n_294),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_199),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_168),
.B(n_199),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_183),
.C(n_192),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_180),
.C(n_182),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_184),
.B1(n_192),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_200),
.B(n_206),
.C(n_207),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_284),
.B(n_285),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_228),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_214),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_220),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_241),
.B(n_283),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_239),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_277),
.B(n_282),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_267),
.B(n_276),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_256),
.B(n_266),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_248),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_265),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_313),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_315),
.Y(n_320)
);


endmodule