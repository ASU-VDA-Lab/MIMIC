module real_jpeg_4512_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_1),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_132),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_132),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_49),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_49),
.B1(n_169),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_2),
.A2(n_49),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_2),
.A2(n_263),
.B(n_266),
.C(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_2),
.B(n_199),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_55),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_303),
.C(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_2),
.B(n_119),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_2),
.B(n_300),
.C(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_2),
.B(n_28),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_3),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_4),
.A2(n_24),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_24),
.B1(n_34),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_4),
.A2(n_24),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_81),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_6),
.A2(n_81),
.B1(n_191),
.B2(n_194),
.Y(n_190)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_8),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_11),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_408),
.B(n_410),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_154),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_152),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_18),
.B(n_133),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_84),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_20),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_20),
.A2(n_135),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_20),
.B(n_161),
.C(n_202),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_20),
.B(n_244),
.C(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_20),
.A2(n_135),
.B1(n_244),
.B2(n_347),
.Y(n_370)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_140)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_23),
.Y(n_130)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_46),
.B1(n_51),
.B2(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_27),
.A2(n_46),
.B(n_51),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_31),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_33),
.Y(n_267)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_49),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_52),
.A2(n_84),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_52),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_52),
.B(n_140),
.C(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_52),
.A2(n_139),
.B1(n_142),
.B2(n_397),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_78),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_53),
.B(n_171),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_54),
.A2(n_65),
.B1(n_164),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_55),
.A2(n_209),
.B(n_213),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_55),
.B(n_165),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_55),
.A2(n_66),
.B1(n_78),
.B2(n_209),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_57),
.Y(n_305)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_66),
.B(n_171),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_70),
.Y(n_301)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B1(n_119),
.B2(n_120),
.Y(n_84)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_93),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_109),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_94),
.A2(n_109),
.B1(n_146),
.B2(n_203),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_94),
.A2(n_109),
.B1(n_146),
.B2(n_203),
.Y(n_244)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_103),
.Y(n_268)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_105),
.Y(n_331)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_127),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_145),
.Y(n_232)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.C(n_141),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_134),
.A2(n_140),
.B1(n_256),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_134),
.Y(n_392)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_221),
.C(n_232),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_140),
.A2(n_232),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_140),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_140),
.A2(n_256),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_140),
.B(n_202),
.C(n_357),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_140),
.A2(n_256),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_141),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_142),
.Y(n_397)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_388),
.B(n_405),
.Y(n_155)
);

OAI211xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_277),
.B(n_382),
.C(n_387),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_249),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_158),
.A2(n_249),
.B(n_383),
.C(n_386),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_233),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_159),
.B(n_233),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_206),
.C(n_220),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_160),
.B(n_206),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_200),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_162),
.A2(n_163),
.B1(n_173),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_162),
.A2(n_163),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_162),
.A2(n_163),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_163),
.B(n_271),
.C(n_314),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_163),
.B(n_339),
.C(n_341),
.Y(n_352)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_181),
.B1(n_189),
.B2(n_196),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_197),
.B(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_178),
.Y(n_307)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_181),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_182),
.A2(n_226),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_182),
.A2(n_226),
.B1(n_272),
.B2(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_201),
.A2(n_202),
.B1(n_230),
.B2(n_298),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_201),
.B(n_298),
.C(n_321),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_201),
.A2(n_202),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_215),
.B2(n_219),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_219),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_215),
.A2(n_239),
.B(n_240),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_216),
.B(n_226),
.Y(n_332)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_223),
.A2(n_230),
.B1(n_298),
.B2(n_373),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_223),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_230),
.A2(n_298),
.B1(n_299),
.B2(n_308),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_247),
.B2(n_248),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_241),
.B1(n_242),
.B2(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_241),
.B(n_246),
.C(n_248),
.Y(n_404)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_244),
.A2(n_343),
.B1(n_344),
.B2(n_347),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_244),
.Y(n_347)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_245),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_245),
.A2(n_394),
.B1(n_398),
.B2(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_250),
.B(n_252),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.C(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_258),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_260),
.B(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_261),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_262),
.A2(n_270),
.B1(n_271),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_262),
.Y(n_364)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_270),
.A2(n_271),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_274),
.Y(n_286)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_366),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_351),
.B(n_365),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_336),
.B(n_350),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_318),
.B(n_335),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_310),
.B(n_317),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_295),
.B(n_309),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_292),
.B(n_294),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_296),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_345),
.C(n_347),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_308),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_320),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_334),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_332),
.B2(n_333),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_333),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_349),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_349),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_341),
.B1(n_342),
.B2(n_348),
.Y(n_337)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_353),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_361),
.C(n_362),
.Y(n_375)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_376),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_375),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_375),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_374),
.C(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_384),
.B(n_385),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_379),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_400),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_393),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.C(n_399),
.Y(n_393)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_399),
.B(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_404),
.Y(n_406)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx13_ASAP7_75t_L g412 ( 
.A(n_409),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);


endmodule