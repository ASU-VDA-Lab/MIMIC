module fake_aes_12521_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
AND2x2_ASAP7_75t_SL g11 ( .A(n_2), .B(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_10), .B(n_0), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_9), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_16) );
BUFx6f_ASAP7_75t_SL g17 ( .A(n_11), .Y(n_17) );
OA21x2_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_13), .B(n_9), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND4xp75_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .C(n_19), .D(n_17), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_17), .B1(n_14), .B2(n_18), .Y(n_22) );
AOI211xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_18), .B(n_3), .C(n_4), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_18), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
OR2x6_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
endmodule