module fake_jpeg_1197_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_40),
.Y(n_41)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_34),
.B1(n_36),
.B2(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_63),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_42),
.C(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_47),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_46),
.B(n_29),
.C(n_44),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_29),
.B(n_15),
.C(n_26),
.D(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_17),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_44),
.B1(n_34),
.B2(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_2),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_14),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_13),
.A3(n_20),
.B1(n_19),
.B2(n_18),
.C1(n_9),
.C2(n_11),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_5),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_12),
.C(n_16),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_79),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_88),
.B(n_86),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_73),
.C(n_24),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_86),
.C(n_85),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_8),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_7),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_94),
.Y(n_95)
);


endmodule