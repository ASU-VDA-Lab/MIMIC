module real_aes_308_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_666;
wire n_320;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_691;
wire n_481;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_0), .A2(n_236), .B1(n_335), .B2(n_339), .Y(n_334) );
INVx1_ASAP7_75t_L g406 ( .A(n_1), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_2), .A2(n_204), .B1(n_460), .B2(n_497), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_3), .A2(n_87), .B1(n_363), .B2(n_570), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_4), .A2(n_129), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g508 ( .A1(n_5), .A2(n_79), .B1(n_237), .B2(n_260), .C1(n_276), .C2(n_290), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_6), .A2(n_62), .B1(n_280), .B2(n_285), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_7), .A2(n_151), .B1(n_313), .B2(n_314), .Y(n_503) );
AO22x2_ASAP7_75t_L g274 ( .A1(n_8), .A2(n_182), .B1(n_263), .B2(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g661 ( .A(n_8), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_9), .A2(n_155), .B1(n_361), .B2(n_363), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_10), .A2(n_57), .B1(n_403), .B2(n_533), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_11), .A2(n_73), .B1(n_380), .B2(n_484), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_12), .A2(n_28), .B1(n_396), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_13), .A2(n_15), .B1(n_545), .B2(n_685), .Y(n_684) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_14), .B(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_16), .A2(n_103), .B1(n_305), .B2(n_307), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_17), .A2(n_184), .B1(n_294), .B2(n_295), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_18), .A2(n_89), .B1(n_313), .B2(n_314), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_19), .A2(n_166), .B1(n_322), .B2(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_20), .A2(n_101), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_21), .A2(n_37), .B1(n_280), .B2(n_285), .Y(n_279) );
AO22x2_ASAP7_75t_L g271 ( .A1(n_22), .A2(n_60), .B1(n_263), .B2(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_22), .B(n_660), .Y(n_659) );
OA22x2_ASAP7_75t_L g620 ( .A1(n_23), .A2(n_621), .B1(n_633), .B2(n_634), .Y(n_620) );
INVx1_ASAP7_75t_L g633 ( .A(n_23), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_24), .A2(n_142), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_25), .A2(n_38), .B1(n_681), .B2(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_26), .A2(n_123), .B1(n_280), .B2(n_285), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_27), .A2(n_189), .B1(n_382), .B2(n_480), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_29), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_30), .A2(n_39), .B1(n_302), .B2(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_31), .A2(n_139), .B1(n_387), .B2(n_477), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_32), .A2(n_176), .B1(n_345), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_33), .A2(n_216), .B1(n_324), .B2(n_484), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_34), .A2(n_229), .B1(n_350), .B2(n_352), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_35), .A2(n_100), .B1(n_347), .B2(n_380), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_36), .A2(n_213), .B1(n_260), .B2(n_276), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_40), .A2(n_214), .B1(n_294), .B2(n_295), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_41), .A2(n_197), .B1(n_350), .B2(n_572), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_42), .A2(n_45), .B1(n_363), .B2(n_404), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_43), .A2(n_226), .B1(n_355), .B2(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_44), .A2(n_232), .B1(n_313), .B2(n_314), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_46), .A2(n_163), .B1(n_392), .B2(n_640), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_47), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_48), .A2(n_199), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_49), .A2(n_160), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_50), .A2(n_196), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_51), .A2(n_145), .B1(n_439), .B2(n_440), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_52), .A2(n_96), .B1(n_363), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_53), .A2(n_67), .B1(n_403), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_54), .A2(n_90), .B1(n_310), .B2(n_311), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_55), .A2(n_107), .B1(n_350), .B2(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_56), .A2(n_201), .B1(n_545), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_58), .A2(n_61), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_59), .A2(n_135), .B1(n_448), .B2(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_63), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_64), .A2(n_218), .B1(n_544), .B2(n_546), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_65), .A2(n_190), .B1(n_345), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_66), .A2(n_191), .B1(n_439), .B2(n_440), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_68), .A2(n_141), .B1(n_206), .B2(n_363), .C1(n_404), .C2(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_69), .A2(n_174), .B1(n_305), .B2(n_307), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_70), .A2(n_130), .B1(n_397), .B2(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g263 ( .A(n_71), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_72), .B(n_527), .Y(n_608) );
XNOR2x2_ASAP7_75t_L g602 ( .A(n_74), .B(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_75), .A2(n_210), .B1(n_294), .B2(n_295), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_76), .A2(n_140), .B1(n_310), .B2(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g409 ( .A(n_77), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_78), .A2(n_113), .B1(n_450), .B2(n_451), .Y(n_449) );
AO22x2_ASAP7_75t_L g521 ( .A1(n_80), .A2(n_522), .B1(n_523), .B2(n_551), .Y(n_521) );
INVx1_ASAP7_75t_L g551 ( .A(n_80), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_81), .B(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_82), .A2(n_168), .B1(n_450), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_83), .A2(n_109), .B1(n_460), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_84), .A2(n_211), .B1(n_387), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_85), .A2(n_114), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx1_ASAP7_75t_SL g268 ( .A(n_86), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_86), .B(n_112), .Y(n_662) );
INVx2_ASAP7_75t_L g249 ( .A(n_88), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_91), .A2(n_149), .B1(n_311), .B2(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_92), .A2(n_148), .B1(n_339), .B2(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_93), .B(n_567), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_94), .A2(n_133), .B1(n_350), .B2(n_437), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_95), .A2(n_106), .B1(n_460), .B2(n_531), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_97), .A2(n_147), .B1(n_392), .B2(n_542), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_98), .A2(n_212), .B1(n_326), .B2(n_477), .Y(n_476) );
OA22x2_ASAP7_75t_L g374 ( .A1(n_99), .A2(n_375), .B1(n_376), .B2(n_410), .Y(n_374) );
INVx1_ASAP7_75t_L g410 ( .A(n_99), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_102), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_104), .A2(n_209), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_105), .A2(n_183), .B1(n_280), .B2(n_285), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_108), .A2(n_208), .B1(n_426), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_110), .A2(n_198), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_111), .A2(n_152), .B1(n_340), .B2(n_383), .Y(n_629) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_112), .A2(n_192), .B1(n_263), .B2(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_115), .B(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_116), .A2(n_185), .B1(n_331), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_117), .A2(n_227), .B1(n_361), .B2(n_363), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_118), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_119), .A2(n_173), .B1(n_363), .B2(n_404), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_120), .A2(n_179), .B1(n_310), .B2(n_311), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_121), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_122), .A2(n_164), .B1(n_387), .B2(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_124), .Y(n_414) );
OA22x2_ASAP7_75t_L g690 ( .A1(n_125), .A2(n_665), .B1(n_666), .B2(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_125), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_126), .A2(n_162), .B1(n_380), .B2(n_484), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_127), .A2(n_207), .B1(n_350), .B2(n_572), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_128), .A2(n_138), .B1(n_326), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_131), .A2(n_171), .B1(n_342), .B2(n_345), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_132), .A2(n_231), .B1(n_450), .B2(n_451), .Y(n_595) );
INVx1_ASAP7_75t_L g269 ( .A(n_134), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_136), .A2(n_165), .B1(n_355), .B2(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_137), .B(n_367), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_143), .A2(n_158), .B1(n_307), .B2(n_389), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_144), .B(n_290), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_146), .A2(n_154), .B1(n_301), .B2(n_302), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_150), .A2(n_170), .B1(n_322), .B2(n_325), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_153), .A2(n_665), .B1(n_666), .B2(n_686), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_153), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_156), .A2(n_222), .B1(n_301), .B2(n_302), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_157), .A2(n_234), .B1(n_310), .B2(n_311), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_159), .A2(n_194), .B1(n_426), .B2(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_161), .A2(n_195), .B1(n_450), .B2(n_451), .Y(n_638) );
INVx1_ASAP7_75t_L g555 ( .A(n_167), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_169), .A2(n_175), .B1(n_355), .B2(n_357), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_172), .A2(n_233), .B1(n_328), .B2(n_331), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_177), .A2(n_186), .B1(n_355), .B2(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_178), .B(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_180), .A2(n_193), .B1(n_383), .B2(n_419), .Y(n_418) );
XNOR2x1_ASAP7_75t_L g318 ( .A(n_181), .B(n_319), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_187), .A2(n_238), .B1(n_352), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_188), .A2(n_202), .B1(n_389), .B2(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_200), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g657 ( .A(n_200), .Y(n_657) );
INVx1_ASAP7_75t_L g245 ( .A(n_203), .Y(n_245) );
AND2x2_ASAP7_75t_R g688 ( .A(n_203), .B(n_657), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g239 ( .A1(n_205), .A2(n_240), .B(n_250), .C(n_663), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_215), .A2(n_221), .B1(n_436), .B2(n_437), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_217), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_220), .Y(n_432) );
INVx1_ASAP7_75t_L g405 ( .A(n_223), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_224), .B(n_363), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_225), .A2(n_235), .B1(n_345), .B2(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_228), .B(n_526), .Y(n_525) );
AO22x1_ASAP7_75t_L g583 ( .A1(n_230), .A2(n_584), .B1(n_598), .B2(n_599), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_230), .Y(n_598) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_SL g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g695 ( .A(n_244), .B(n_246), .Y(n_695) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_245), .B(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_515), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_250) );
INVx1_ASAP7_75t_L g653 ( .A(n_251), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_468), .B1(n_513), .B2(n_514), .Y(n_251) );
INVx1_ASAP7_75t_L g514 ( .A(n_252), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_372), .B1(n_466), .B2(n_467), .Y(n_252) );
INVx1_ASAP7_75t_L g467 ( .A(n_253), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B1(n_316), .B2(n_370), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
XOR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_315), .Y(n_255) );
NAND2x1_ASAP7_75t_SL g256 ( .A(n_257), .B(n_298), .Y(n_256) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_258), .B(n_288), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_279), .Y(n_258) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_270), .Y(n_260) );
AND2x2_ASAP7_75t_L g301 ( .A(n_261), .B(n_281), .Y(n_301) );
AND2x6_ASAP7_75t_L g310 ( .A(n_261), .B(n_291), .Y(n_310) );
AND2x2_ASAP7_75t_L g330 ( .A(n_261), .B(n_291), .Y(n_330) );
AND2x2_ASAP7_75t_L g338 ( .A(n_261), .B(n_281), .Y(n_338) );
AND2x4_ASAP7_75t_L g356 ( .A(n_261), .B(n_270), .Y(n_356) );
AND2x2_ASAP7_75t_L g439 ( .A(n_261), .B(n_270), .Y(n_439) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_261), .B(n_281), .Y(n_505) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
AND2x2_ASAP7_75t_L g278 ( .A(n_262), .B(n_266), .Y(n_278) );
INVx2_ASAP7_75t_L g284 ( .A(n_262), .Y(n_284) );
BUFx2_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx1_ASAP7_75t_L g264 ( .A(n_263), .Y(n_264) );
OAI22x1_ASAP7_75t_L g266 ( .A1(n_263), .A2(n_267), .B1(n_268), .B2(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_263), .Y(n_267) );
INVx2_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
INVx1_ASAP7_75t_L g275 ( .A(n_263), .Y(n_275) );
AND2x4_ASAP7_75t_L g306 ( .A(n_265), .B(n_284), .Y(n_306) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g283 ( .A(n_266), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
AND2x4_ASAP7_75t_L g294 ( .A(n_270), .B(n_283), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_270), .B(n_306), .Y(n_307) );
AND2x4_ASAP7_75t_L g326 ( .A(n_270), .B(n_306), .Y(n_326) );
AND2x2_ASAP7_75t_L g362 ( .A(n_270), .B(n_283), .Y(n_362) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
INVx1_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
AND2x2_ASAP7_75t_L g297 ( .A(n_271), .B(n_274), .Y(n_297) );
INVxp67_ASAP7_75t_L g277 ( .A(n_273), .Y(n_277) );
AND2x4_ASAP7_75t_L g291 ( .A(n_273), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_274), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x4_ASAP7_75t_L g359 ( .A(n_277), .B(n_278), .Y(n_359) );
AND2x2_ASAP7_75t_L g440 ( .A(n_277), .B(n_278), .Y(n_440) );
AND2x2_ASAP7_75t_L g285 ( .A(n_278), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g290 ( .A(n_278), .B(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g353 ( .A(n_278), .B(n_286), .Y(n_353) );
AND2x2_ASAP7_75t_L g369 ( .A(n_278), .B(n_291), .Y(n_369) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AND2x6_ASAP7_75t_L g311 ( .A(n_281), .B(n_306), .Y(n_311) );
AND2x4_ASAP7_75t_L g333 ( .A(n_281), .B(n_306), .Y(n_333) );
AND2x2_ASAP7_75t_L g351 ( .A(n_281), .B(n_283), .Y(n_351) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_282), .Y(n_287) );
AND2x2_ASAP7_75t_L g313 ( .A(n_283), .B(n_291), .Y(n_313) );
AND2x4_ASAP7_75t_L g324 ( .A(n_283), .B(n_291), .Y(n_324) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_293), .Y(n_288) );
INVx2_ASAP7_75t_SL g431 ( .A(n_290), .Y(n_431) );
BUFx2_ASAP7_75t_L g648 ( .A(n_290), .Y(n_648) );
AND2x2_ASAP7_75t_L g305 ( .A(n_291), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g344 ( .A(n_291), .B(n_306), .Y(n_344) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g364 ( .A(n_296), .B(n_297), .Y(n_364) );
AND2x4_ASAP7_75t_L g302 ( .A(n_297), .B(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g314 ( .A(n_297), .B(n_306), .Y(n_314) );
AND2x4_ASAP7_75t_L g340 ( .A(n_297), .B(n_303), .Y(n_340) );
AND2x4_ASAP7_75t_L g347 ( .A(n_297), .B(n_306), .Y(n_347) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_299), .B(n_308), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_304), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVx1_ASAP7_75t_L g422 ( .A(n_310), .Y(n_422) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_318), .Y(n_371) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_348), .Y(n_319) );
NAND4xp25_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .C(n_334), .D(n_341), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g447 ( .A(n_323), .Y(n_447) );
INVx1_ASAP7_75t_SL g549 ( .A(n_323), .Y(n_549) );
INVx3_ASAP7_75t_L g594 ( .A(n_323), .Y(n_594) );
INVx6_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_326), .Y(n_392) );
INVx2_ASAP7_75t_L g428 ( .A(n_326), .Y(n_428) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_326), .Y(n_561) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_326), .Y(n_597) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
INVx2_ASAP7_75t_L g477 ( .A(n_329), .Y(n_477) );
INVx2_ASAP7_75t_SL g577 ( .A(n_329), .Y(n_577) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g445 ( .A(n_330), .Y(n_445) );
BUFx2_ASAP7_75t_L g545 ( .A(n_330), .Y(n_545) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g387 ( .A(n_332), .Y(n_387) );
INVx2_ASAP7_75t_SL g486 ( .A(n_332), .Y(n_486) );
INVx2_ASAP7_75t_L g546 ( .A(n_332), .Y(n_546) );
INVx2_ASAP7_75t_L g631 ( .A(n_332), .Y(n_631) );
INVx8_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
INVx1_ASAP7_75t_L g479 ( .A(n_337), .Y(n_479) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_338), .Y(n_450) );
BUFx3_ASAP7_75t_L g682 ( .A(n_338), .Y(n_682) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g419 ( .A(n_340), .Y(n_419) );
BUFx3_ASAP7_75t_L g451 ( .A(n_340), .Y(n_451) );
INVx5_ASAP7_75t_SL g481 ( .A(n_340), .Y(n_481) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx4_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
INVx3_ASAP7_75t_L g426 ( .A(n_343), .Y(n_426) );
INVx2_ASAP7_75t_SL g453 ( .A(n_343), .Y(n_453) );
INVx2_ASAP7_75t_L g542 ( .A(n_343), .Y(n_542) );
INVx3_ASAP7_75t_SL g640 ( .A(n_343), .Y(n_640) );
INVx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g448 ( .A(n_346), .Y(n_448) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g484 ( .A(n_347), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g348 ( .A(n_349), .B(n_354), .C(n_360), .D(n_365), .Y(n_348) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_351), .Y(n_436) );
INVx3_ASAP7_75t_L g458 ( .A(n_351), .Y(n_458) );
BUFx4f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g400 ( .A(n_353), .Y(n_400) );
BUFx6f_ASAP7_75t_SL g437 ( .A(n_353), .Y(n_437) );
BUFx3_ASAP7_75t_L g572 ( .A(n_353), .Y(n_572) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g460 ( .A(n_356), .Y(n_460) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx2_ASAP7_75t_L g497 ( .A(n_358), .Y(n_497) );
INVx2_ASAP7_75t_L g531 ( .A(n_358), .Y(n_531) );
INVx2_ASAP7_75t_L g588 ( .A(n_358), .Y(n_588) );
INVx2_ASAP7_75t_SL g671 ( .A(n_358), .Y(n_671) );
INVx6_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx5_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
INVx2_ASAP7_75t_L g492 ( .A(n_362), .Y(n_492) );
INVx2_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g535 ( .A(n_364), .Y(n_535) );
INVx3_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx3_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g463 ( .A(n_368), .Y(n_463) );
INVx4_ASAP7_75t_SL g527 ( .A(n_368), .Y(n_527) );
INVx4_ASAP7_75t_SL g567 ( .A(n_368), .Y(n_567) );
INVx6_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g466 ( .A(n_372), .Y(n_466) );
AOI22x1_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_411), .B2(n_412), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_393), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_384), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_380), .Y(n_677) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_389), .Y(n_575) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_401), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .Y(n_394) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g539 ( .A(n_400), .Y(n_539) );
OAI222xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_406), .B2(n_407), .C1(n_408), .C2(n_409), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OA22x2_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_441), .B1(n_464), .B2(n_465), .Y(n_412) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_413), .Y(n_465) );
XNOR2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_416), .B(n_429), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_423), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_432), .B(n_433), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_431), .A2(n_489), .B(n_490), .C(n_493), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
BUFx6f_ASAP7_75t_SL g537 ( .A(n_436), .Y(n_537) );
BUFx2_ASAP7_75t_SL g674 ( .A(n_437), .Y(n_674) );
INVx1_ASAP7_75t_L g464 ( .A(n_441), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_443), .B(n_455), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .C(n_449), .D(n_452), .Y(n_443) );
BUFx2_ASAP7_75t_L g679 ( .A(n_453), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .C(n_461), .D(n_462), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_463), .Y(n_669) );
INVx1_ASAP7_75t_L g513 ( .A(n_468), .Y(n_513) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OA22x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_499), .B2(n_512), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
XOR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_498), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_487), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g563 ( .A(n_481), .Y(n_563) );
INVx2_ASAP7_75t_L g683 ( .A(n_481), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g570 ( .A(n_492), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g512 ( .A(n_499), .Y(n_512) );
XNOR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .C(n_504), .D(n_506), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g652 ( .A(n_515), .Y(n_652) );
AOI22xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_517), .B1(n_617), .B2(n_618), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_580), .B2(n_581), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_552), .B2(n_579), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_540), .Y(n_523) );
NAND4xp25_ASAP7_75t_SL g524 ( .A(n_525), .B(n_528), .C(n_532), .D(n_536), .Y(n_524) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .C(n_547), .D(n_548), .Y(n_540) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g579 ( .A(n_552), .Y(n_579) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_564), .B2(n_578), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_557), .B(n_565), .C(n_573), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_561), .Y(n_685) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_573), .Y(n_564) );
NAND4xp25_ASAP7_75t_SL g565 ( .A(n_566), .B(n_568), .C(n_569), .D(n_571), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_600), .B1(n_614), .B2(n_615), .Y(n_581) );
INVx1_ASAP7_75t_L g614 ( .A(n_582), .Y(n_614) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g599 ( .A(n_584), .Y(n_599) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_591), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_589), .D(n_590), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .C(n_595), .D(n_596), .Y(n_591) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g616 ( .A(n_602), .Y(n_616) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_609), .Y(n_603) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .C(n_607), .D(n_608), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .C(n_612), .D(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AO22x1_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_635), .B1(n_650), .B2(n_651), .Y(n_619) );
INVx1_ASAP7_75t_L g650 ( .A(n_620), .Y(n_650) );
INVx1_ASAP7_75t_L g634 ( .A(n_621), .Y(n_634) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_627), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .C(n_625), .D(n_626), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .C(n_630), .D(n_632), .Y(n_627) );
INVx1_ASAP7_75t_SL g651 ( .A(n_635), .Y(n_651) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_649), .Y(n_635) );
NAND4xp75_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .C(n_644), .D(n_647), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_656), .B(n_659), .Y(n_694) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OAI222xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_687), .B1(n_689), .B2(n_691), .C1(n_692), .C2(n_695), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_675), .Y(n_666) );
NAND4xp25_ASAP7_75t_SL g667 ( .A(n_668), .B(n_670), .C(n_672), .D(n_673), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .C(n_680), .D(n_684), .Y(n_675) );
BUFx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_693), .Y(n_692) );
CKINVDCx6p67_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
endmodule