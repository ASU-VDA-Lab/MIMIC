module fake_jpeg_14849_n_346 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_71),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_36),
.B(n_27),
.C(n_22),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_22),
.B(n_27),
.C(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_34),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_66),
.B1(n_33),
.B2(n_16),
.Y(n_111)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_33),
.B1(n_20),
.B2(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_20),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_86),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_95),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_84),
.Y(n_135)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_110),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_18),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_39),
.C(n_62),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_26),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_23),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_16),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_119)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_18),
.B1(n_49),
.B2(n_38),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_43),
.B1(n_29),
.B2(n_31),
.Y(n_122)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_74),
.B1(n_72),
.B2(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_58),
.B(n_24),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_22),
.C(n_35),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_114),
.B1(n_96),
.B2(n_89),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_39),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_75),
.B(n_99),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_127),
.B1(n_134),
.B2(n_136),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_43),
.B1(n_29),
.B2(n_38),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_39),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_139),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_62),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_40),
.B1(n_38),
.B2(n_56),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_40),
.B1(n_39),
.B2(n_19),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_35),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_39),
.C(n_62),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_40),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_106),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_143),
.A2(n_170),
.B1(n_172),
.B2(n_175),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_106),
.B1(n_88),
.B2(n_77),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_145),
.A2(n_148),
.B1(n_167),
.B2(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_79),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_120),
.B1(n_142),
.B2(n_116),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_150),
.B(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_157),
.B(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_158),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_106),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_105),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_173),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_101),
.B1(n_85),
.B2(n_104),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_166),
.B1(n_129),
.B2(n_135),
.Y(n_182)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_90),
.B1(n_91),
.B2(n_102),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_81),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_84),
.B1(n_19),
.B2(n_109),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_123),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_17),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_62),
.B1(n_19),
.B2(n_32),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_197),
.B1(n_203),
.B2(n_208),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_188),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_139),
.C(n_132),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_149),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_136),
.C(n_135),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_174),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_113),
.B1(n_114),
.B2(n_121),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_201),
.B(n_171),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_30),
.B(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_17),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_186),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_32),
.B1(n_10),
.B2(n_14),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_158),
.B(n_14),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_173),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_28),
.B1(n_76),
.B2(n_17),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_168),
.B1(n_163),
.B2(n_13),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_214),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_167),
.B1(n_159),
.B2(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_215),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_149),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_191),
.B(n_179),
.C(n_196),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_209),
.B1(n_203),
.B2(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_149),
.C(n_162),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_226),
.C(n_230),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_176),
.C(n_151),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_150),
.C(n_146),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_195),
.C(n_179),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_233),
.C(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_155),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_166),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_76),
.C(n_28),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_239),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_200),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_254),
.C(n_233),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_246),
.A2(n_249),
.B1(n_261),
.B2(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_177),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_260),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_200),
.B1(n_183),
.B2(n_192),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_225),
.Y(n_254)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_184),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_208),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_240),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_184),
.B1(n_187),
.B2(n_2),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_268),
.Y(n_285)
);

FAx1_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_215),
.CI(n_229),
.CON(n_265),
.SN(n_265)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_242),
.A2(n_222),
.B(n_212),
.C(n_238),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_244),
.B(n_255),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_231),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_239),
.B1(n_237),
.B2(n_212),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_230),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_272),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_236),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_279),
.C(n_251),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_21),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_281),
.Y(n_290)
);

XOR2x1_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_211),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_21),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_21),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_256),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_0),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

AO221x1_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_301)
);

BUFx12f_ASAP7_75t_SL g286 ( 
.A(n_276),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_295),
.B(n_267),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_291),
.C(n_264),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_256),
.C(n_254),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_243),
.B1(n_248),
.B2(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_297),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_273),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_246),
.B1(n_250),
.B2(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_280),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_265),
.A2(n_3),
.B(n_4),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_267),
.B(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_314),
.B(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_310),
.B1(n_315),
.B2(n_297),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_267),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_287),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_285),
.C(n_304),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_3),
.B(n_5),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_295),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_299),
.A2(n_6),
.B(n_7),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_320),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_321),
.B(n_308),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_291),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_289),
.C(n_296),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_326),
.B(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_313),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_288),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_330),
.B(n_332),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_302),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_331),
.B(n_334),
.Y(n_339)
);

OA21x2_ASAP7_75t_SL g337 ( 
.A1(n_329),
.A2(n_326),
.B(n_321),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_338),
.B(n_315),
.Y(n_341)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_318),
.B(n_324),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_330),
.C(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_339),
.B(n_335),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_7),
.B(n_8),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_9),
.Y(n_346)
);


endmodule