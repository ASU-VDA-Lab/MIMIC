module fake_jpeg_13849_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_36),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_31),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_54),
.B(n_57),
.Y(n_80)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_64),
.B1(n_66),
.B2(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_43),
.B1(n_40),
.B2(n_31),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_24),
.B1(n_20),
.B2(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_16),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_45),
.B1(n_37),
.B2(n_39),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_28),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_62),
.C(n_65),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_82),
.C(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_30),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_22),
.B(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_50),
.Y(n_109)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_57),
.C(n_54),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_34),
.Y(n_96)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_51),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_50),
.B1(n_74),
.B2(n_73),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_79),
.C(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_118),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_122),
.B(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_86),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_128),
.B(n_106),
.C(n_97),
.D(n_93),
.Y(n_134)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_124),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_72),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_70),
.C(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_85),
.B1(n_45),
.B2(n_91),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_93),
.B1(n_99),
.B2(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_94),
.B1(n_106),
.B2(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_135),
.B1(n_124),
.B2(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

NOR4xp25_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_117),
.C(n_116),
.D(n_125),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_99),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_141),
.B(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_119),
.C(n_131),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_144),
.C(n_146),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_122),
.C(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_122),
.B1(n_111),
.B2(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_102),
.C(n_74),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_130),
.B(n_140),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_89),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_51),
.C(n_87),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_135),
.B1(n_134),
.B2(n_141),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_144),
.C(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_1),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_156),
.C(n_155),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_21),
.B(n_30),
.C(n_7),
.D(n_11),
.Y(n_158)
);

AOI31xp33_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_148),
.A3(n_12),
.B(n_14),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_50),
.B(n_58),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_143),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_162),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_165),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_154),
.B1(n_8),
.B2(n_9),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_4),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_161),
.A3(n_8),
.B1(n_12),
.B2(n_14),
.C1(n_2),
.C2(n_4),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_1),
.C(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_170),
.Y(n_176)
);


endmodule