module fake_jpeg_11563_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_0),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_55),
.B1(n_78),
.B2(n_64),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_77),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_64),
.B1(n_78),
.B2(n_55),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_106),
.B1(n_57),
.B2(n_68),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_66),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_74),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_59),
.B1(n_65),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_65),
.B1(n_53),
.B2(n_57),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_71),
.B1(n_76),
.B2(n_73),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_102),
.B1(n_98),
.B2(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_115),
.B1(n_117),
.B2(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_124),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_7),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_81),
.B1(n_62),
.B2(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_68),
.B1(n_75),
.B2(n_82),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_63),
.C(n_58),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_12),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_56),
.B(n_2),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_118),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_148),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_151),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_7),
.B(n_8),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_35),
.C(n_51),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_158),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_34),
.B1(n_49),
.B2(n_47),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_167),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_9),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_150),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_10),
.B(n_11),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_131),
.B(n_142),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_163),
.A2(n_133),
.B1(n_142),
.B2(n_151),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_13),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_177),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_144),
.B(n_27),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_155),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_52),
.B1(n_29),
.B2(n_33),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_179),
.B1(n_170),
.B2(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_164),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_186),
.B(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_171),
.B(n_164),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_185),
.B1(n_172),
.B2(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_187),
.B(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_183),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_153),
.B(n_186),
.C(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_167),
.C(n_38),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_24),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_39),
.Y(n_199)
);


endmodule