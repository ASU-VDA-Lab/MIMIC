module fake_netlist_1_5044_n_525 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_525);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_525;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g76 ( .A(n_41), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_53), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_57), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_47), .Y(n_79) );
INVxp33_ASAP7_75t_L g80 ( .A(n_7), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_56), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_44), .Y(n_82) );
BUFx10_ASAP7_75t_L g83 ( .A(n_65), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_55), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_46), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_24), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_37), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_50), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_66), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_60), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_3), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_75), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_40), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_32), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_64), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_49), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_28), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_48), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_25), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_11), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_86), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_86), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_106), .Y(n_122) );
OR2x6_ASAP7_75t_L g123 ( .A(n_94), .B(n_29), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_94), .B(n_0), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_108), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_108), .B(n_1), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_109), .B(n_1), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx2_ASAP7_75t_SL g137 ( .A(n_113), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_128), .B(n_91), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_121), .B(n_109), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_113), .B(n_96), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_114), .B(n_100), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_121), .B(n_102), .Y(n_143) );
INVx1_ASAP7_75t_SL g144 ( .A(n_121), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_121), .B(n_111), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_124), .B(n_101), .Y(n_146) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_114), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_115), .B(n_104), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_124), .B(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_124), .B(n_83), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_124), .B(n_93), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_130), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_117), .B(n_80), .Y(n_161) );
INVx8_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_161), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_160), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_161), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_161), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g168 ( .A1(n_147), .A2(n_128), .B(n_132), .C(n_133), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_147), .A2(n_132), .B1(n_128), .B2(n_125), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_160), .B(n_117), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_149), .B(n_128), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_137), .B(n_125), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_138), .B(n_126), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_156), .B(n_126), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_146), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_138), .A2(n_132), .B1(n_127), .B2(n_123), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_149), .B(n_132), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_138), .B(n_127), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_146), .B(n_123), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_149), .B(n_85), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_146), .B(n_123), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_149), .B(n_123), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_141), .B(n_151), .C(n_142), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_188), .B(n_143), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_187), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_163), .B(n_154), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_138), .B1(n_146), .B2(n_145), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_175), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_175), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_187), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_187), .A2(n_145), .B1(n_143), .B2(n_144), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_183), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_165), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_187), .B(n_144), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_169), .A2(n_123), .B1(n_142), .B2(n_141), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_169), .A2(n_151), .B1(n_131), .B2(n_133), .Y(n_216) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_188), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_167), .B(n_143), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_173), .B(n_158), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_188), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_187), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_183), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_173), .B(n_191), .Y(n_225) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_191), .B(n_79), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_196), .A2(n_174), .B(n_180), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_197), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_191), .B1(n_178), .B2(n_190), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_215), .A2(n_179), .B1(n_191), .B2(n_192), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g231 ( .A1(n_226), .A2(n_112), .B1(n_95), .B2(n_158), .Y(n_231) );
OAI221xp5_ASAP7_75t_L g232 ( .A1(n_218), .A2(n_179), .B1(n_177), .B2(n_190), .C(n_192), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_205), .A2(n_185), .B1(n_193), .B2(n_158), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_196), .A2(n_171), .B(n_172), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_226), .A2(n_81), .B1(n_92), .B2(n_97), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_196), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_185), .B1(n_181), .B2(n_176), .Y(n_237) );
NOR2xp67_ASAP7_75t_SL g238 ( .A(n_207), .B(n_208), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_222), .B(n_204), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_212), .A2(n_193), .B1(n_177), .B2(n_176), .Y(n_240) );
NOR2xp67_ASAP7_75t_SL g241 ( .A(n_207), .B(n_166), .Y(n_241) );
OAI22xp5_ASAP7_75t_SL g242 ( .A1(n_199), .A2(n_88), .B1(n_105), .B2(n_85), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_223), .A2(n_193), .B1(n_143), .B2(n_145), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_225), .B(n_145), .Y(n_246) );
CKINVDCx11_ASAP7_75t_R g247 ( .A(n_198), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_201), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_216), .A2(n_135), .B1(n_134), .B2(n_168), .C(n_133), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_219), .A2(n_88), .B1(n_186), .B2(n_166), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_202), .A2(n_181), .B1(n_172), .B2(n_186), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_202), .B(n_186), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_222), .B(n_186), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_243), .B(n_248), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_219), .B1(n_225), .B2(n_223), .Y(n_255) );
OAI211xp5_ASAP7_75t_L g256 ( .A1(n_228), .A2(n_135), .B(n_134), .C(n_194), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_216), .B1(n_210), .B2(n_224), .C(n_131), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_209), .B1(n_200), .B2(n_222), .Y(n_258) );
AOI211xp5_ASAP7_75t_L g259 ( .A1(n_235), .A2(n_103), .B(n_209), .C(n_213), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_195), .B1(n_210), .B2(n_224), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_243), .B(n_195), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_248), .B(n_198), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_246), .B(n_195), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_246), .A2(n_220), .B1(n_217), .B2(n_195), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_252), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_240), .B(n_198), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_245), .A2(n_220), .B1(n_217), .B2(n_120), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_239), .Y(n_271) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_232), .A2(n_206), .B1(n_211), .B2(n_204), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_242), .A2(n_198), .B1(n_189), .B2(n_211), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_227), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
OAI211xp5_ASAP7_75t_L g276 ( .A1(n_249), .A2(n_131), .B(n_116), .C(n_84), .Y(n_276) );
OAI33xp33_ASAP7_75t_L g277 ( .A1(n_258), .A2(n_99), .A3(n_116), .B1(n_105), .B2(n_107), .B3(n_89), .Y(n_277) );
BUFx12f_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_264), .B(n_244), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g281 ( .A(n_259), .B(n_118), .C(n_122), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_254), .B(n_244), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_247), .B1(n_229), .B2(n_239), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_258), .A2(n_233), .B1(n_250), .B2(n_239), .Y(n_284) );
BUFx4f_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_259), .A2(n_251), .B1(n_234), .B2(n_206), .Y(n_286) );
AOI33xp33_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_116), .A3(n_136), .B1(n_159), .B2(n_155), .B3(n_139), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_256), .A2(n_267), .B1(n_268), .B2(n_276), .C(n_257), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_269), .A2(n_247), .B1(n_253), .B2(n_120), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_271), .A2(n_253), .B1(n_120), .B2(n_130), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_263), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_267), .B(n_130), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g293 ( .A1(n_273), .A2(n_130), .B1(n_89), .B2(n_107), .C(n_221), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_130), .B1(n_122), .B2(n_118), .C(n_129), .Y(n_294) );
INVx11_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
OAI31xp33_ASAP7_75t_SL g297 ( .A1(n_266), .A2(n_253), .A3(n_238), .B(n_5), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_298), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_284), .A2(n_270), .B1(n_265), .B2(n_272), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_298), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_279), .B(n_275), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
OAI31xp33_ASAP7_75t_L g305 ( .A1(n_284), .A2(n_270), .A3(n_274), .B(n_275), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_277), .A2(n_118), .B1(n_122), .B2(n_119), .C(n_129), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_280), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_278), .B(n_275), .Y(n_309) );
NAND4xp25_ASAP7_75t_SL g310 ( .A(n_289), .B(n_2), .C(n_4), .D(n_5), .Y(n_310) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_155), .A3(n_159), .B1(n_136), .B2(n_7), .B3(n_8), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_278), .A2(n_238), .B1(n_241), .B2(n_204), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_296), .B(n_118), .Y(n_314) );
BUFx2_ASAP7_75t_SL g315 ( .A(n_282), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_282), .B(n_118), .Y(n_317) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_281), .B(n_118), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_285), .B(n_129), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_292), .B(n_129), .Y(n_320) );
AOI33xp33_ASAP7_75t_L g321 ( .A1(n_283), .A2(n_139), .A3(n_148), .B1(n_152), .B2(n_157), .B3(n_9), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_129), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_157), .B(n_139), .Y(n_323) );
O2A1O1Ixp5_ASAP7_75t_L g324 ( .A1(n_285), .A2(n_241), .B(n_148), .C(n_152), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_288), .B(n_122), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_289), .A2(n_211), .B1(n_206), .B2(n_122), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_308), .B(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_308), .B(n_297), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_328), .B(n_2), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_328), .B(n_4), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_305), .B(n_290), .C(n_294), .D(n_293), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_312), .B(n_287), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_129), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_328), .B(n_6), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_299), .B(n_129), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_301), .B(n_122), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_326), .B(n_150), .C(n_153), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_315), .B(n_6), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_302), .B(n_8), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_315), .B(n_9), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_328), .B(n_10), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_11), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_316), .B(n_12), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_305), .B(n_14), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_309), .B(n_14), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_300), .B(n_15), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_320), .B(n_15), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_300), .B(n_16), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_320), .B(n_16), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_325), .B(n_17), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_325), .B(n_214), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_325), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_321), .B(n_17), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_323), .B(n_18), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_323), .B(n_18), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_349), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_363), .B(n_310), .Y(n_375) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_348), .B(n_318), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_354), .B(n_322), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_332), .B(n_318), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_359), .B(n_322), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_330), .B(n_319), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_348), .B(n_313), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_332), .B(n_319), .Y(n_383) );
NAND2x1_ASAP7_75t_L g384 ( .A(n_350), .B(n_313), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_330), .B(n_327), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_346), .B(n_327), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_340), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_306), .Y(n_388) );
NOR2x1_ASAP7_75t_SL g389 ( .A(n_350), .B(n_311), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_331), .B(n_157), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_363), .B(n_19), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_331), .B(n_152), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_329), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_360), .B(n_21), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_355), .B(n_148), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_339), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_358), .B(n_22), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_372), .B(n_324), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_349), .B(n_153), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_150), .B1(n_153), .B2(n_221), .C(n_203), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_361), .B(n_23), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_342), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_343), .Y(n_404) );
OAI21xp33_ASAP7_75t_SL g405 ( .A1(n_371), .A2(n_26), .B(n_27), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_355), .B(n_153), .Y(n_406) );
NAND2x1_ASAP7_75t_SL g407 ( .A(n_333), .B(n_31), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_356), .B(n_153), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_345), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_352), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g411 ( .A(n_367), .B(n_214), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_366), .B(n_371), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_368), .B(n_153), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_352), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_369), .B(n_33), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_362), .Y(n_417) );
AOI211x1_ASAP7_75t_L g418 ( .A1(n_365), .A2(n_34), .B(n_35), .C(n_36), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_362), .B(n_38), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_337), .B(n_42), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_344), .B(n_43), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_417), .B(n_364), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_375), .A2(n_341), .B1(n_334), .B2(n_351), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_376), .B(n_364), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_410), .B(n_414), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
INVx3_ASAP7_75t_SL g430 ( .A(n_378), .Y(n_430) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_380), .B(n_357), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_373), .B(n_372), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_375), .B(n_357), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_412), .B(n_344), .Y(n_434) );
INVxp33_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
XNOR2xp5_ASAP7_75t_L g437 ( .A(n_377), .B(n_353), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_383), .B(n_347), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_387), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_382), .B(n_336), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_403), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g443 ( .A(n_379), .B(n_45), .Y(n_443) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_412), .B(n_214), .Y(n_444) );
OAI32xp33_ASAP7_75t_L g445 ( .A1(n_405), .A2(n_51), .A3(n_54), .B1(n_58), .B2(n_59), .Y(n_445) );
XOR2xp5_ASAP7_75t_L g446 ( .A(n_385), .B(n_61), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_382), .B(n_214), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_396), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g450 ( .A1(n_391), .A2(n_170), .B(n_184), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_399), .B(n_214), .C(n_208), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_397), .B(n_62), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_409), .B(n_63), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_386), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_399), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_390), .Y(n_457) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_391), .A2(n_221), .B(n_203), .C(n_70), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_409), .B(n_68), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_392), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_407), .A2(n_214), .B(n_208), .C(n_207), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_388), .B(n_69), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_398), .B(n_71), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_415), .B(n_72), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_419), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_378), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_408), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_401), .B(n_208), .C(n_207), .Y(n_470) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_418), .B(n_203), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_388), .Y(n_472) );
XNOR2x1_ASAP7_75t_L g473 ( .A(n_411), .B(n_221), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_413), .Y(n_474) );
AOI211xp5_ASAP7_75t_L g475 ( .A1(n_398), .A2(n_182), .B(n_208), .C(n_394), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_421), .Y(n_476) );
XNOR2x1_ASAP7_75t_L g477 ( .A(n_402), .B(n_208), .Y(n_477) );
AOI311xp33_ASAP7_75t_L g478 ( .A1(n_394), .A2(n_375), .A3(n_414), .B(n_410), .C(n_108), .Y(n_478) );
AOI211xp5_ASAP7_75t_SL g479 ( .A1(n_400), .A2(n_375), .B(n_325), .C(n_334), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_416), .B(n_410), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_373), .A2(n_375), .B1(n_350), .B2(n_348), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_381), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_378), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_436), .A2(n_440), .B(n_479), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_436), .A2(n_440), .B(n_435), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_423), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_433), .A2(n_481), .B1(n_456), .B2(n_454), .C(n_435), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_479), .B(n_424), .C(n_478), .D(n_433), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_481), .A2(n_424), .B1(n_456), .B2(n_472), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_426), .B(n_482), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_482), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_449), .B(n_431), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_458), .A2(n_448), .B(n_451), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_425), .A2(n_430), .B1(n_468), .B2(n_466), .C(n_437), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_448), .A2(n_444), .B(n_461), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_475), .B(n_464), .C(n_458), .D(n_468), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_444), .A2(n_443), .B(n_425), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_427), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_428), .A2(n_432), .B(n_439), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_476), .B1(n_457), .B2(n_483), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_441), .B(n_442), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_488), .A2(n_445), .B(n_471), .C(n_470), .Y(n_502) );
NOR3x1_ASAP7_75t_L g503 ( .A(n_484), .B(n_480), .C(n_438), .Y(n_503) );
NAND4xp75_ASAP7_75t_L g504 ( .A(n_497), .B(n_462), .C(n_422), .D(n_453), .Y(n_504) );
NOR2x1p5_ASAP7_75t_L g505 ( .A(n_496), .B(n_483), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_491), .Y(n_506) );
OAI21xp33_ASAP7_75t_SL g507 ( .A1(n_487), .A2(n_477), .B(n_447), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_489), .B(n_434), .Y(n_508) );
NOR2x1p5_ASAP7_75t_L g509 ( .A(n_492), .B(n_467), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_485), .A2(n_465), .B(n_460), .C(n_452), .Y(n_510) );
OAI211xp5_ASAP7_75t_SL g511 ( .A1(n_494), .A2(n_450), .B(n_474), .C(n_463), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_506), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_507), .A2(n_511), .B1(n_506), .B2(n_502), .C(n_510), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_505), .A2(n_500), .B1(n_495), .B2(n_491), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g515 ( .A(n_508), .B(n_493), .C(n_446), .Y(n_515) );
OAI222xp33_ASAP7_75t_L g516 ( .A1(n_503), .A2(n_490), .B1(n_501), .B2(n_486), .C1(n_498), .C2(n_447), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_512), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_514), .Y(n_518) );
OR3x2_ASAP7_75t_L g519 ( .A(n_515), .B(n_509), .C(n_504), .Y(n_519) );
XNOR2xp5_ASAP7_75t_L g520 ( .A(n_518), .B(n_513), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_518), .A2(n_499), .B1(n_516), .B2(n_469), .C(n_473), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_520), .A2(n_519), .B1(n_517), .B2(n_465), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_522), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_523), .A2(n_521), .B1(n_459), .B2(n_455), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_524), .B(n_429), .Y(n_525) );
endmodule