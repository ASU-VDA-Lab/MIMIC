module fake_jpeg_9854_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_4),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_5),
.Y(n_88)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_4),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_55),
.B1(n_46),
.B2(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_63),
.B1(n_62),
.B2(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_58),
.B1(n_50),
.B2(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_59),
.B1(n_57),
.B2(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_48),
.B1(n_25),
.B2(n_26),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_27),
.B1(n_11),
.B2(n_14),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_8),
.B1(n_15),
.B2(n_16),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_93),
.B1(n_86),
.B2(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_44),
.B1(n_20),
.B2(n_21),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_107),
.C(n_112),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_110),
.B1(n_101),
.B2(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_108),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_102),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_93),
.B1(n_113),
.B2(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_109),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_111),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_110),
.B(n_34),
.C(n_35),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_30),
.C(n_39),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);


endmodule