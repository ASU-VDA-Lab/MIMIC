module fake_jpeg_88_n_615 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_65),
.Y(n_170)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_95),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_93),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_10),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_10),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_24),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_104),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_28),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_29),
.B(n_10),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_50),
.B1(n_30),
.B2(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_151),
.B1(n_158),
.B2(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_37),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_22),
.B1(n_46),
.B2(n_47),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_37),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_38),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_154),
.B(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_77),
.B(n_28),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_89),
.A2(n_54),
.B1(n_22),
.B2(n_46),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_35),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_161),
.B(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_25),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_35),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_31),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_62),
.A2(n_50),
.B1(n_30),
.B2(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_58),
.B(n_31),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_76),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_179),
.Y(n_265)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_180),
.B(n_183),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_109),
.B1(n_107),
.B2(n_69),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_181),
.A2(n_209),
.B1(n_223),
.B2(n_233),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_118),
.A2(n_26),
.B1(n_50),
.B2(n_23),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_182),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_185),
.Y(n_295)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_193),
.Y(n_283)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_194),
.Y(n_278)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_120),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_196),
.B(n_201),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_23),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_200),
.B(n_220),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_114),
.B(n_54),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_203),
.B(n_169),
.C(n_48),
.Y(n_284)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_205),
.Y(n_280)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_206),
.Y(n_282)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_112),
.B1(n_102),
.B2(n_100),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_212),
.Y(n_257)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_134),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_216),
.Y(n_242)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_221),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_225),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_27),
.B1(n_41),
.B2(n_94),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_239),
.B1(n_47),
.B2(n_61),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_137),
.B(n_47),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_224),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_132),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_124),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_127),
.Y(n_261)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_230),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_130),
.B(n_64),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_229),
.B(n_48),
.Y(n_296)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_234),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_138),
.A2(n_97),
.B1(n_96),
.B2(n_88),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_240),
.Y(n_243)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_142),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_140),
.A2(n_26),
.B1(n_44),
.B2(n_48),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_136),
.B1(n_140),
.B2(n_26),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_141),
.A2(n_82),
.B1(n_80),
.B2(n_79),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_146),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_128),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_247),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_246),
.A2(n_270),
.B1(n_194),
.B2(n_188),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_147),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_250),
.A2(n_187),
.B1(n_231),
.B2(n_197),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_178),
.A2(n_74),
.B1(n_71),
.B2(n_57),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_260),
.A2(n_266),
.B1(n_267),
.B2(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_261),
.B(n_222),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_153),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_153),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_203),
.A2(n_78),
.B1(n_59),
.B2(n_139),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_209),
.A2(n_139),
.B1(n_127),
.B2(n_162),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_202),
.A2(n_146),
.B1(n_134),
.B2(n_164),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_200),
.A2(n_191),
.B1(n_228),
.B2(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_192),
.A2(n_162),
.B1(n_123),
.B2(n_46),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_275),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_284),
.B(n_266),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_184),
.B(n_206),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_293),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_189),
.B(n_164),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_199),
.B(n_169),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_232),
.C(n_225),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

OAI22x1_ASAP7_75t_L g300 ( 
.A1(n_263),
.A2(n_240),
.B1(n_198),
.B2(n_211),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_300),
.B(n_285),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_301),
.B(n_326),
.Y(n_362)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_263),
.A2(n_195),
.B1(n_204),
.B2(n_190),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_303),
.A2(n_308),
.B1(n_321),
.B2(n_327),
.Y(n_364)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_305),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_247),
.A2(n_213),
.A3(n_224),
.B1(n_235),
.B2(n_193),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_306),
.B(n_324),
.Y(n_359)
);

XOR2x2_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_240),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_SL g354 ( 
.A(n_307),
.B(n_273),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_245),
.A2(n_221),
.B1(n_216),
.B2(n_217),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_227),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_310),
.B(n_323),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_325),
.B(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_328),
.Y(n_351)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_318),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_317),
.A2(n_320),
.B1(n_330),
.B2(n_331),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_264),
.A2(n_215),
.B1(n_207),
.B2(n_233),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_260),
.A2(n_262),
.B1(n_279),
.B2(n_267),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_244),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_279),
.A2(n_250),
.B1(n_253),
.B2(n_275),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_218),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_248),
.A2(n_236),
.B1(n_230),
.B2(n_44),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_334),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_218),
.B1(n_54),
.B2(n_186),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_257),
.A2(n_54),
.B1(n_41),
.B2(n_27),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_12),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_344),
.B(n_346),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_253),
.A2(n_65),
.B1(n_36),
.B2(n_43),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_65),
.B1(n_55),
.B2(n_43),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_335),
.A2(n_339),
.B1(n_341),
.B2(n_278),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_343),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_249),
.A2(n_55),
.B(n_43),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_337),
.A2(n_335),
.B(n_339),
.Y(n_384)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_342),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_243),
.A2(n_55),
.B1(n_43),
.B2(n_2),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_248),
.B(n_55),
.C(n_1),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_273),
.C(n_285),
.Y(n_360)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_11),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_293),
.A2(n_243),
.B1(n_287),
.B2(n_281),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_297),
.B1(n_280),
.B2(n_273),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_243),
.B(n_0),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g386 ( 
.A1(n_348),
.A2(n_259),
.B(n_290),
.C(n_3),
.D(n_4),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_328),
.A2(n_272),
.B1(n_292),
.B2(n_254),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_350),
.A2(n_341),
.B1(n_302),
.B2(n_299),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_354),
.B(n_366),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_304),
.A2(n_258),
.B1(n_269),
.B2(n_254),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_367),
.B1(n_369),
.B2(n_377),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_386),
.C(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_365),
.B(n_373),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_287),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_304),
.A2(n_258),
.B1(n_292),
.B2(n_272),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_289),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_371),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_280),
.C(n_295),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_372),
.A2(n_381),
.B(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_285),
.C(n_286),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_242),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_319),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_291),
.B1(n_286),
.B2(n_242),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_346),
.A2(n_291),
.B1(n_242),
.B2(n_259),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_378),
.A2(n_385),
.B1(n_393),
.B2(n_308),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_259),
.B1(n_277),
.B2(n_283),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_379),
.A2(n_388),
.B1(n_392),
.B2(n_364),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_319),
.A2(n_278),
.B(n_252),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_310),
.B(n_277),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_344),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_301),
.A2(n_252),
.B1(n_283),
.B2(n_291),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_346),
.A2(n_290),
.B1(n_1),
.B2(n_3),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_0),
.C(n_1),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_298),
.B(n_0),
.C(n_1),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_4),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_298),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_394),
.B(n_396),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_347),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_404),
.Y(n_452)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_359),
.A2(n_337),
.B(n_330),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_399),
.A2(n_402),
.B(n_429),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_351),
.B(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_400),
.B(n_418),
.Y(n_463)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_359),
.A2(n_326),
.B(n_348),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_382),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_405),
.B(n_410),
.Y(n_461)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_406),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_407),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_438)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_409),
.B(n_416),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_387),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_417),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_364),
.A2(n_300),
.B1(n_320),
.B2(n_303),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_365),
.A2(n_300),
.B1(n_324),
.B2(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_334),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_356),
.B(n_327),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_367),
.A2(n_309),
.B1(n_312),
.B2(n_329),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_422),
.B1(n_424),
.B2(n_426),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_387),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_427),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_342),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_421),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_388),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_357),
.A2(n_338),
.B1(n_315),
.B2(n_313),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_380),
.A2(n_361),
.B1(n_378),
.B2(n_381),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_362),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_379),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_428),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_372),
.A2(n_305),
.B(n_331),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_358),
.A2(n_322),
.B1(n_340),
.B2(n_4),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_430),
.A2(n_376),
.B1(n_391),
.B2(n_386),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_432),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_352),
.C(n_368),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_440),
.C(n_444),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_352),
.C(n_371),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_407),
.A2(n_426),
.B1(n_401),
.B2(n_398),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_442),
.A2(n_445),
.B1(n_429),
.B2(n_414),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_354),
.C(n_373),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_362),
.B1(n_384),
.B2(n_353),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_360),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_453),
.C(n_458),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_390),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_411),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_400),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_395),
.A2(n_355),
.B(n_375),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_455),
.A2(n_468),
.B(n_397),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_355),
.C(n_375),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_389),
.C(n_376),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_460),
.C(n_464),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_389),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_462),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_402),
.B(n_393),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_399),
.B(n_322),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_469),
.C(n_431),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_395),
.B(n_12),
.CI(n_18),
.CON(n_466),
.SN(n_466)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_412),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_405),
.A2(n_13),
.B(n_18),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_19),
.Y(n_469)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_438),
.A2(n_428),
.B1(n_403),
.B2(n_413),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_471),
.A2(n_478),
.B1(n_496),
.B2(n_498),
.Y(n_508)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_480),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_477),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_441),
.A2(n_403),
.B1(n_415),
.B2(n_422),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_444),
.B(n_412),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_479),
.B(n_447),
.Y(n_506)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_437),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_483),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_437),
.B(n_410),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_453),
.Y(n_503)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_486),
.Y(n_526)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_488),
.Y(n_509)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_490),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_446),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_491),
.B(n_492),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_468),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_442),
.A2(n_421),
.B1(n_419),
.B2(n_430),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_452),
.A2(n_420),
.B1(n_424),
.B2(n_418),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_443),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_497),
.A2(n_14),
.B(n_8),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_432),
.B1(n_416),
.B2(n_406),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_499),
.A2(n_500),
.B1(n_501),
.B2(n_436),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_408),
.B1(n_6),
.B2(n_8),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_515),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_445),
.B(n_465),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_504),
.A2(n_525),
.B1(n_474),
.B2(n_486),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_506),
.B(n_516),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_SL g507 ( 
.A(n_472),
.B(n_448),
.C(n_434),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_507),
.B(n_482),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_440),
.C(n_458),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_513),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_511),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_473),
.B(n_459),
.C(n_460),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_472),
.B(n_455),
.C(n_464),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_514),
.B(n_520),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_457),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_479),
.B(n_467),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_452),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_18),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_439),
.C(n_463),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_480),
.C(n_498),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_527),
.C(n_497),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_462),
.B1(n_408),
.B2(n_469),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_483),
.B(n_466),
.C(n_5),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_471),
.A2(n_466),
.B1(n_6),
.B2(n_8),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g545 ( 
.A(n_528),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_529),
.A2(n_500),
.B(n_499),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_487),
.B(n_9),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_488),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_532),
.B(n_537),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_534),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_513),
.B(n_478),
.C(n_485),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_546),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_539),
.B(n_520),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_474),
.C(n_493),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_543),
.C(n_548),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_514),
.B(n_494),
.C(n_501),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_549),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_502),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_547),
.B(n_526),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_495),
.C(n_477),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_529),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_508),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_551),
.A2(n_525),
.B1(n_505),
.B2(n_523),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_523),
.B(n_526),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_553),
.A2(n_562),
.B(n_532),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_556),
.B(n_564),
.Y(n_576)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_524),
.C(n_515),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_563),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_545),
.A2(n_519),
.B1(n_522),
.B2(n_534),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_560),
.A2(n_549),
.B1(n_542),
.B2(n_535),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_540),
.A2(n_519),
.B(n_521),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_538),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_531),
.B(n_506),
.C(n_516),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_567),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_548),
.B(n_530),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_551),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_569),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_543),
.B(n_527),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_570),
.B(n_16),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_536),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_573),
.Y(n_593)
);

XOR2x2_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_578),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_535),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_553),
.A2(n_547),
.B(n_542),
.Y(n_574)
);

OAI21x1_ASAP7_75t_SL g591 ( 
.A1(n_574),
.A2(n_583),
.B(n_570),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_577),
.A2(n_578),
.B1(n_556),
.B2(n_561),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_560),
.A2(n_563),
.B1(n_557),
.B2(n_555),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_5),
.C(n_16),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_581),
.B(n_582),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_566),
.B(n_555),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_558),
.B(n_17),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_561),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_564),
.B(n_17),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_585),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_590),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_554),
.B(n_569),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_589),
.A2(n_572),
.B(n_580),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_559),
.C(n_554),
.Y(n_590)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_591),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_567),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_585),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_594),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_568),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_595),
.B(n_596),
.Y(n_598)
);

MAJx2_ASAP7_75t_L g606 ( 
.A(n_600),
.B(n_603),
.C(n_565),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_593),
.A2(n_586),
.B1(n_577),
.B2(n_574),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_602),
.B(n_597),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_599),
.B(n_596),
.C(n_592),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_606),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_604),
.B(n_588),
.Y(n_607)
);

AO21x1_ASAP7_75t_L g609 ( 
.A1(n_607),
.A2(n_608),
.B(n_598),
.Y(n_609)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_609),
.Y(n_612)
);

OAI21x1_ASAP7_75t_SL g611 ( 
.A1(n_610),
.A2(n_598),
.B(n_601),
.Y(n_611)
);

AO21x1_ASAP7_75t_L g613 ( 
.A1(n_611),
.A2(n_597),
.B(n_581),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_612),
.C(n_17),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_17),
.Y(n_615)
);


endmodule