module fake_netlist_5_1403_n_71 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_71);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_71;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_53;
wire n_42;
wire n_64;
wire n_45;
wire n_46;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_70;
wire n_38;
wire n_61;
wire n_68;
wire n_35;
wire n_41;
wire n_32;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_57;
wire n_37;
wire n_59;
wire n_30;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_39;

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_3),
.B(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_10),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_42),
.B1(n_34),
.B2(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_45),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_14),
.Y(n_55)
);

AOI221xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_38),
.B1(n_37),
.B2(n_43),
.C(n_31),
.Y(n_56)
);

OAI221xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_36),
.B1(n_43),
.B2(n_40),
.C(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B(n_55),
.C(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_48),
.B1(n_54),
.B2(n_47),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_R g63 ( 
.A(n_59),
.B(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_58),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_65),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule