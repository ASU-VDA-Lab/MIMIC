module fake_jpeg_29536_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_29),
.B1(n_18),
.B2(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_22),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_30),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_28),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_75),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_67),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_77),
.B1(n_40),
.B2(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_70),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_35),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_80),
.C(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_24),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_33),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_74),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_32),
.B(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_39),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_40),
.B1(n_39),
.B2(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_31),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_16),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_65),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_79),
.B1(n_81),
.B2(n_59),
.Y(n_110)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_39),
.A3(n_8),
.B1(n_9),
.B2(n_14),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_13),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_5),
.Y(n_119)
);

AO21x1_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_5),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_120),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_82),
.B1(n_68),
.B2(n_63),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_118),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_59),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_121),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_72),
.B1(n_73),
.B2(n_69),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_5),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_91),
.B(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_96),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_100),
.B(n_88),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_118),
.C(n_120),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_144),
.C(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_86),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_118),
.C(n_113),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_110),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_136),
.B1(n_124),
.B2(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_126),
.B1(n_90),
.B2(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_154),
.B1(n_146),
.B2(n_140),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_127),
.B(n_135),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_153),
.A2(n_146),
.B(n_144),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_135),
.B1(n_123),
.B2(n_129),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_125),
.C(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_87),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_154),
.B(n_150),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_155),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_140),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.C(n_101),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

AOI31xp33_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_149),
.A3(n_153),
.B(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_123),
.C(n_101),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OA21x2_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_159),
.B(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_172),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_165),
.B(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_166),
.B(n_92),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_85),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_10),
.Y(n_178)
);


endmodule