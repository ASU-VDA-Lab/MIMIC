module fake_netlist_6_3840_n_1788 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1788);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1788;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVxp67_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_163),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_137),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_199),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_55),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_107),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_162),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_136),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_218),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_5),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_158),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_11),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_147),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_239),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_134),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_70),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_159),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_165),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_120),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_250),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_53),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_54),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_41),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_175),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_205),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_252),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_60),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_123),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_21),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_31),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_73),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_45),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_81),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_224),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_232),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_20),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_90),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_124),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_53),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_13),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_254),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_135),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_108),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_60),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_154),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_105),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_131),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_87),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_231),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_212),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_1),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_174),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_96),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_23),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_183),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_167),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_256),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_216),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_153),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_213),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_66),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_128),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_16),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_33),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_146),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_177),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_141),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_81),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_191),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_161),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_244),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_80),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_253),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_46),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_233),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_104),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_197),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_198),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_55),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_58),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_74),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_32),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_14),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_43),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_226),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_119),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_229),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_164),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_246),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_21),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_51),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_188),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_85),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_75),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_223),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_91),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_50),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_248),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_68),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_132),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_222),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_12),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_150),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_85),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_129),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_20),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_12),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_145),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_25),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_127),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_74),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_186),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_24),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_214),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_217),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_166),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_83),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_103),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_138),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_187),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_33),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_207),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_89),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_148),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_225),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_37),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_171),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_94),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_114),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_241),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_251),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_79),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_113),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_83),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_118),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_240),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_40),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_219),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_92),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_38),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_220),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_180),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_176),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_204),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_9),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_7),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_71),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_63),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_84),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_235),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_47),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_42),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_31),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_6),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_77),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_190),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_238),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_116),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_39),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_196),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_290),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_276),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_295),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_284),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_266),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_276),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_398),
.B(n_0),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_306),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_266),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_284),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_307),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_311),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_316),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_282),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_258),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_309),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_353),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_319),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_309),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_322),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_329),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_343),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_346),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_420),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_329),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_355),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_357),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_284),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_380),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_380),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_286),
.B(n_0),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_286),
.B(n_1),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_336),
.B(n_2),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_265),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_260),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_293),
.Y(n_494)
);

BUFx2_ASAP7_75t_SL g495 ( 
.A(n_399),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_336),
.B(n_3),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_299),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_362),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_261),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_303),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_269),
.B(n_3),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_263),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_348),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_364),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_368),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_305),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_317),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_367),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_399),
.B(n_4),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_332),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_264),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_289),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_374),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_292),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_333),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_368),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_296),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_275),
.B(n_4),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_368),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_377),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_381),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_265),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_388),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_395),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_347),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_366),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_257),
.B(n_6),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_375),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_378),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_352),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_297),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_383),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_298),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_531),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_438),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_531),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_469),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_348),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_472),
.B(n_275),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_531),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_492),
.B(n_312),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_454),
.A2(n_302),
.B1(n_397),
.B2(n_274),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_270),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_496),
.B(n_312),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_495),
.B(n_270),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_492),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_500),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_495),
.B(n_271),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_503),
.B(n_271),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_511),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_519),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_496),
.B(n_272),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_526),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_460),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_466),
.B(n_272),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_530),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_534),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_344),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_489),
.B(n_273),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_493),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_501),
.B(n_273),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_490),
.B(n_352),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_450),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_480),
.B(n_344),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_457),
.A2(n_354),
.B(n_268),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_455),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_459),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_280),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_465),
.B(n_328),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_463),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_354),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_473),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_269),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_451),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_554),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_582),
.B(n_352),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_473),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_557),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_554),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_556),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_582),
.B(n_352),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_419),
.B1(n_391),
.B2(n_393),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_582),
.B(n_429),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_583),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_557),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_552),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_547),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_566),
.B(n_265),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_580),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_566),
.B(n_265),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_580),
.B(n_476),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_586),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_429),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_566),
.B(n_265),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_536),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_536),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_582),
.B(n_476),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_536),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_582),
.B(n_429),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_566),
.B(n_429),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_536),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_566),
.B(n_265),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_587),
.B(n_478),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_552),
.A2(n_419),
.B1(n_433),
.B2(n_390),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_589),
.B(n_478),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_545),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_549),
.A2(n_302),
.B1(n_397),
.B2(n_274),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_547),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_547),
.B(n_265),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_545),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_479),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_539),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_545),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_552),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_541),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_552),
.B(n_591),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_579),
.B(n_590),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_589),
.B(n_479),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_539),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_587),
.B(n_482),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_579),
.B(n_482),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_545),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_552),
.B(n_259),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_545),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_628),
.B(n_567),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_607),
.B(n_589),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_628),
.B(n_567),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_607),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_648),
.B(n_604),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_581),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_664),
.B(n_590),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_607),
.Y(n_679)
);

OAI221xp5_ASAP7_75t_L g680 ( 
.A1(n_618),
.A2(n_551),
.B1(n_581),
.B2(n_549),
.C(n_574),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_624),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_625),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_662),
.B(n_551),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_650),
.B(n_568),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_662),
.B(n_664),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_664),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_624),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_629),
.A2(n_552),
.B1(n_590),
.B2(n_591),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_659),
.B(n_604),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_659),
.B(n_604),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_616),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_553),
.Y(n_694)
);

AOI221x1_ASAP7_75t_L g695 ( 
.A1(n_627),
.A2(n_602),
.B1(n_598),
.B2(n_605),
.C(n_593),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_610),
.A2(n_605),
.B1(n_602),
.B2(n_598),
.Y(n_696)
);

INVx8_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_663),
.B(n_552),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_666),
.B(n_553),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_616),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_616),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_562),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_650),
.A2(n_552),
.B1(n_590),
.B2(n_591),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_667),
.B(n_562),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_653),
.B(n_481),
.C(n_598),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_632),
.B(n_590),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_667),
.B(n_598),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_632),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_SL g709 ( 
.A(n_618),
.B(n_589),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_663),
.A2(n_599),
.B(n_602),
.C(n_603),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_624),
.B(n_573),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_650),
.B(n_589),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_651),
.B(n_602),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_608),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_650),
.B(n_589),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_612),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_642),
.A2(n_589),
.B1(n_593),
.B2(n_592),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_592),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_658),
.B(n_592),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_654),
.B(n_592),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_658),
.B(n_592),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_633),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_608),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_654),
.B(n_592),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_654),
.B(n_592),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_613),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_654),
.B(n_593),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_651),
.A2(n_593),
.B1(n_597),
.B2(n_595),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_654),
.B(n_593),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_615),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_624),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_608),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_609),
.B(n_593),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_658),
.B(n_593),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_668),
.B(n_595),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_614),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_609),
.B(n_595),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_633),
.B(n_570),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_665),
.B(n_568),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_668),
.B(n_595),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_627),
.A2(n_599),
.B(n_603),
.C(n_596),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_617),
.B(n_595),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_617),
.B(n_595),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_655),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_668),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_614),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_665),
.B(n_568),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_621),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_619),
.B(n_595),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_631),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_655),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_649),
.B(n_597),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_670),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_676),
.A2(n_661),
.B(n_670),
.C(n_636),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_702),
.B(n_452),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_697),
.B(n_753),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_743),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_707),
.B(n_597),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_SL g764 ( 
.A(n_675),
.B(n_653),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_704),
.B(n_597),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_672),
.B(n_597),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_688),
.Y(n_767)
);

AOI21x1_ASAP7_75t_L g768 ( 
.A1(n_736),
.A2(n_644),
.B(n_619),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_674),
.B(n_597),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_712),
.A2(n_644),
.B(n_620),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_683),
.B(n_597),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_679),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_682),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_750),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_682),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_749),
.A2(n_756),
.B(n_710),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_715),
.A2(n_620),
.B(n_631),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_568),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_684),
.Y(n_779)
);

CKINVDCx10_ASAP7_75t_R g780 ( 
.A(n_705),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_706),
.B(n_599),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_724),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_684),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_706),
.B(n_636),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_694),
.B(n_647),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_680),
.A2(n_574),
.B(n_645),
.C(n_563),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_708),
.B(n_550),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_719),
.A2(n_620),
.B(n_647),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_699),
.B(n_563),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_708),
.B(n_678),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_688),
.B(n_594),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_722),
.A2(n_728),
.B(n_727),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_687),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_678),
.B(n_649),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_603),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_456),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_690),
.A2(n_468),
.B1(n_477),
.B2(n_474),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_697),
.B(n_485),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_730),
.A2(n_620),
.B(n_645),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_749),
.A2(n_626),
.B(n_622),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_681),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_732),
.A2(n_620),
.B(n_661),
.Y(n_802)
);

AOI21x1_ASAP7_75t_L g803 ( 
.A1(n_742),
.A2(n_623),
.B(n_622),
.Y(n_803)
);

AOI21xp33_ASAP7_75t_L g804 ( 
.A1(n_744),
.A2(n_600),
.B(n_537),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_687),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_721),
.B(n_601),
.C(n_517),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_691),
.B(n_623),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_698),
.B(n_695),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_755),
.A2(n_661),
.B(n_611),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_673),
.B(n_486),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_693),
.Y(n_811)
);

AO21x1_ASAP7_75t_L g812 ( 
.A1(n_709),
.A2(n_278),
.B(n_277),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_755),
.A2(n_686),
.B(n_703),
.Y(n_813)
);

AND2x6_ASAP7_75t_L g814 ( 
.A(n_681),
.B(n_661),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_696),
.A2(n_412),
.B1(n_596),
.B2(n_588),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_743),
.B(n_499),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_723),
.B(n_502),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_692),
.B(n_746),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_698),
.A2(n_611),
.B(n_623),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_752),
.A2(n_600),
.B(n_586),
.C(n_588),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_681),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_737),
.B(n_512),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_695),
.A2(n_626),
.B(n_622),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_758),
.A2(n_552),
.B1(n_635),
.B2(n_570),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_611),
.B(n_622),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_681),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_SL g827 ( 
.A(n_739),
.B(n_515),
.C(n_513),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_748),
.A2(n_611),
.B(n_626),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_693),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_745),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_681),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_758),
.B(n_626),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_731),
.B(n_630),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_689),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_697),
.B(n_718),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_700),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_754),
.A2(n_611),
.B(n_630),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_697),
.B(n_518),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_716),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_757),
.A2(n_611),
.B(n_630),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_734),
.B(n_630),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_711),
.A2(n_611),
.B(n_634),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_734),
.A2(n_412),
.B1(n_436),
.B2(n_434),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_689),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_711),
.B(n_634),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_711),
.A2(n_611),
.B(n_634),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_709),
.A2(n_634),
.B(n_641),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_689),
.A2(n_646),
.B(n_641),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_689),
.B(n_541),
.Y(n_849)
);

AO21x1_ASAP7_75t_L g850 ( 
.A1(n_716),
.A2(n_294),
.B(n_291),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_685),
.B(n_532),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_689),
.A2(n_646),
.B(n_641),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_685),
.A2(n_646),
.B(n_641),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_714),
.A2(n_614),
.B(n_637),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_720),
.B(n_606),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_720),
.A2(n_646),
.B(n_641),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_726),
.A2(n_646),
.B(n_641),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_726),
.A2(n_646),
.B(n_641),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_811),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_776),
.A2(n_813),
.B(n_786),
.C(n_785),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_784),
.A2(n_646),
.B(n_641),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_760),
.B(n_535),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_764),
.B(n_483),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_789),
.B(n_729),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_827),
.B(n_483),
.Y(n_865)
);

CKINVDCx10_ASAP7_75t_R g866 ( 
.A(n_761),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_829),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_820),
.A2(n_584),
.B(n_541),
.C(n_729),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_781),
.B(n_733),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_762),
.B(n_606),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_778),
.A2(n_584),
.B(n_738),
.C(n_733),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_765),
.B(n_738),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_771),
.A2(n_803),
.B(n_788),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_815),
.A2(n_359),
.B(n_279),
.C(n_301),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_774),
.B(n_606),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_836),
.Y(n_876)
);

OAI21xp33_ASAP7_75t_L g877 ( 
.A1(n_816),
.A2(n_504),
.B(n_498),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_793),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_792),
.A2(n_652),
.B(n_646),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_782),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_773),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_804),
.B(n_700),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_SL g883 ( 
.A(n_806),
.B(n_504),
.C(n_498),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_796),
.B(n_509),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_766),
.A2(n_769),
.B(n_853),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_772),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_821),
.Y(n_888)
);

CKINVDCx11_ASAP7_75t_R g889 ( 
.A(n_761),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_821),
.B(n_701),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_835),
.A2(n_652),
.B(n_701),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_851),
.B(n_573),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_810),
.A2(n_514),
.B(n_509),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_790),
.B(n_514),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_805),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_855),
.B(n_521),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_826),
.B(n_714),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_826),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_826),
.B(n_717),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_834),
.B(n_717),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_817),
.A2(n_522),
.B1(n_524),
.B2(n_521),
.Y(n_902)
);

CKINVDCx14_ASAP7_75t_R g903 ( 
.A(n_797),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_761),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_779),
.Y(n_905)
);

AO22x1_ASAP7_75t_L g906 ( 
.A1(n_822),
.A2(n_522),
.B1(n_525),
.B2(n_524),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_783),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_815),
.A2(n_304),
.B(n_310),
.C(n_300),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_767),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_795),
.B(n_725),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_777),
.A2(n_652),
.B(n_725),
.Y(n_911)
);

O2A1O1Ixp5_ASAP7_75t_L g912 ( 
.A1(n_763),
.A2(n_751),
.B(n_740),
.C(n_741),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_834),
.B(n_844),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_797),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_834),
.B(n_735),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_839),
.B(n_735),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_844),
.B(n_740),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_844),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_814),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_776),
.A2(n_751),
.B1(n_741),
.B2(n_585),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_768),
.A2(n_638),
.B(n_637),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_801),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_794),
.A2(n_585),
.B1(n_267),
.B2(n_400),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_832),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_830),
.B(n_525),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_849),
.A2(n_652),
.B(n_638),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_791),
.B(n_506),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_838),
.A2(n_484),
.B(n_351),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_770),
.A2(n_652),
.B(n_638),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_799),
.A2(n_652),
.B(n_638),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_801),
.B(n_652),
.Y(n_931)
);

AND2x4_ASAP7_75t_SL g932 ( 
.A(n_831),
.B(n_578),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_818),
.B(n_573),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_759),
.A2(n_831),
.B1(n_808),
.B2(n_824),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_845),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_833),
.A2(n_639),
.B(n_637),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_807),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_798),
.B(n_652),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_842),
.A2(n_846),
.B(n_809),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_814),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_848),
.A2(n_639),
.B(n_637),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_814),
.B(n_578),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_843),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_843),
.A2(n_446),
.B1(n_288),
.B2(n_427),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_800),
.B(n_808),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_800),
.A2(n_585),
.B1(n_287),
.B2(n_315),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_787),
.B(n_841),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_814),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_802),
.B(n_578),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_812),
.A2(n_314),
.B(n_324),
.C(n_320),
.Y(n_950)
);

AOI221xp5_ASAP7_75t_L g951 ( 
.A1(n_850),
.A2(n_440),
.B1(n_441),
.B2(n_439),
.C(n_438),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_819),
.B(n_640),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_780),
.B(n_520),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_854),
.B(n_640),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_878),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_896),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_874),
.A2(n_847),
.B(n_840),
.C(n_825),
.Y(n_957)
);

AOI221x1_ASAP7_75t_L g958 ( 
.A1(n_860),
.A2(n_934),
.B1(n_886),
.B2(n_939),
.C(n_885),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_864),
.A2(n_857),
.B1(n_858),
.B2(n_856),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_925),
.B(n_828),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_879),
.A2(n_837),
.B(n_823),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_889),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_862),
.B(n_280),
.Y(n_964)
);

NOR2x1_ASAP7_75t_R g965 ( 
.A(n_922),
.B(n_281),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_881),
.Y(n_966)
);

AO31x2_ASAP7_75t_L g967 ( 
.A1(n_860),
.A2(n_852),
.A3(n_823),
.B(n_325),
.Y(n_967)
);

AO31x2_ASAP7_75t_L g968 ( 
.A1(n_920),
.A2(n_326),
.A3(n_335),
.B(n_334),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_875),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_880),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_SL g971 ( 
.A1(n_938),
.A2(n_854),
.B(n_341),
.C(n_342),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_909),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_945),
.A2(n_635),
.B(n_639),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_SL g974 ( 
.A1(n_938),
.A2(n_345),
.B(n_360),
.C(n_338),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_SL g975 ( 
.A(n_885),
.B(n_862),
.C(n_863),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_872),
.A2(n_643),
.B(n_639),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_919),
.B(n_328),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_933),
.A2(n_656),
.B(n_643),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_863),
.A2(n_392),
.B(n_396),
.C(n_384),
.Y(n_979)
);

BUFx12f_ASAP7_75t_L g980 ( 
.A(n_870),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_914),
.A2(n_373),
.B1(n_328),
.B2(n_327),
.Y(n_981)
);

AOI221xp5_ASAP7_75t_SL g982 ( 
.A1(n_908),
.A2(n_564),
.B1(n_571),
.B2(n_555),
.C(n_575),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_919),
.A2(n_882),
.B(n_869),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_903),
.A2(n_313),
.B1(n_318),
.B2(n_308),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_904),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_948),
.B(n_555),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_897),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_948),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_927),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_943),
.A2(n_373),
.B1(n_262),
.B2(n_403),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_945),
.A2(n_656),
.B(n_643),
.Y(n_991)
);

AO31x2_ASAP7_75t_L g992 ( 
.A1(n_946),
.A2(n_404),
.A3(n_411),
.B(n_410),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_924),
.B(n_937),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_SL g994 ( 
.A(n_877),
.B(n_440),
.C(n_439),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_935),
.B(n_947),
.Y(n_995)
);

O2A1O1Ixp5_ASAP7_75t_SL g996 ( 
.A1(n_882),
.A2(n_561),
.B(n_564),
.C(n_560),
.Y(n_996)
);

CKINVDCx8_ASAP7_75t_R g997 ( 
.A(n_866),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_947),
.B(n_635),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_905),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_888),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_911),
.A2(n_656),
.B(n_643),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_895),
.B(n_560),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_888),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_883),
.B(n_561),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_918),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_895),
.B(n_281),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_927),
.B(n_571),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_918),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_940),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_893),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_923),
.A2(n_575),
.B(n_425),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_893),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_921),
.A2(n_657),
.B(n_656),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_907),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_929),
.A2(n_660),
.B(n_657),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_930),
.A2(n_418),
.A3(n_437),
.B(n_428),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_926),
.A2(n_660),
.B(n_657),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_949),
.A2(n_660),
.B(n_657),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_894),
.A2(n_285),
.B(n_423),
.C(n_283),
.Y(n_1020)
);

NAND3xp33_ASAP7_75t_SL g1021 ( 
.A(n_865),
.B(n_442),
.C(n_441),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_861),
.A2(n_671),
.B(n_660),
.Y(n_1022)
);

AO31x2_ASAP7_75t_L g1023 ( 
.A1(n_891),
.A2(n_952),
.A3(n_941),
.B(n_954),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_910),
.A2(n_671),
.A3(n_540),
.B(n_546),
.Y(n_1024)
);

OA21x2_ASAP7_75t_L g1025 ( 
.A1(n_936),
.A2(n_671),
.B(n_540),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_865),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_902),
.B(n_373),
.Y(n_1028)
);

AOI221x1_ASAP7_75t_L g1029 ( 
.A1(n_928),
.A2(n_544),
.B1(n_546),
.B2(n_542),
.C(n_558),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_906),
.B(n_867),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_SL g1031 ( 
.A1(n_871),
.A2(n_671),
.B(n_585),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_873),
.A2(n_542),
.B(n_544),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_876),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_892),
.B(n_283),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_912),
.A2(n_890),
.B(n_898),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_SL g1036 ( 
.A(n_940),
.B(n_442),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_953),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_868),
.A2(n_635),
.B(n_640),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_951),
.A2(n_953),
.B1(n_944),
.B2(n_942),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_548),
.A3(n_538),
.B(n_558),
.Y(n_1040)
);

AOI31xp67_ASAP7_75t_L g1041 ( 
.A1(n_931),
.A2(n_542),
.A3(n_548),
.B(n_538),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_944),
.B(n_285),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_890),
.A2(n_669),
.B(n_640),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_913),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_899),
.B(n_635),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_899),
.B(n_423),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_913),
.A2(n_559),
.B(n_558),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_932),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_931),
.A2(n_900),
.B(n_898),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_900),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_901),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_901),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_915),
.B(n_635),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_915),
.B(n_640),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_917),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_917),
.A2(n_669),
.B(n_548),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_950),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_875),
.B(n_446),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_889),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_887),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_860),
.A2(n_635),
.B(n_669),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_864),
.A2(n_405),
.B1(n_421),
.B2(n_401),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_864),
.B(n_635),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_886),
.A2(n_669),
.B(n_545),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_955),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_985),
.B(n_559),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1006),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1065),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1006),
.Y(n_1070)
);

OAI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_975),
.A2(n_430),
.B1(n_431),
.B2(n_426),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1007),
.A2(n_446),
.B1(n_430),
.B2(n_431),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_997),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_956),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_970),
.Y(n_1075)
);

INVx6_ASAP7_75t_L g1076 ( 
.A(n_1009),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1060),
.Y(n_1077)
);

OAI22x1_ASAP7_75t_SL g1078 ( 
.A1(n_1026),
.A2(n_426),
.B1(n_323),
.B2(n_330),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_972),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_964),
.A2(n_635),
.B1(n_542),
.B2(n_331),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_966),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_988),
.B(n_1006),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_999),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_988),
.B(n_669),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_977),
.A2(n_337),
.B1(n_339),
.B2(n_321),
.Y(n_1085)
);

INVx6_ASAP7_75t_L g1086 ( 
.A(n_963),
.Y(n_1086)
);

BUFx2_ASAP7_75t_SL g1087 ( 
.A(n_963),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_983),
.A2(n_635),
.B(n_565),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_980),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1028),
.A2(n_542),
.B1(n_340),
.B2(n_407),
.Y(n_1090)
);

BUFx2_ASAP7_75t_SL g1091 ( 
.A(n_963),
.Y(n_1091)
);

BUFx2_ASAP7_75t_SL g1092 ( 
.A(n_1001),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1000),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1011),
.B(n_559),
.Y(n_1094)
);

BUFx2_ASAP7_75t_SL g1095 ( 
.A(n_962),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_994),
.A2(n_408),
.B1(n_350),
.B2(n_356),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_989),
.A2(n_409),
.B1(n_358),
.B2(n_361),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1015),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1013),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1039),
.A2(n_414),
.B1(n_369),
.B2(n_370),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1027),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1003),
.B(n_565),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1033),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1021),
.A2(n_415),
.B1(n_371),
.B2(n_372),
.Y(n_1104)
);

INVx6_ASAP7_75t_L g1105 ( 
.A(n_1059),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1004),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_993),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1042),
.A2(n_1012),
.B1(n_990),
.B2(n_981),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_977),
.A2(n_416),
.B1(n_376),
.B2(n_379),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_1030),
.Y(n_1110)
);

BUFx4f_ASAP7_75t_L g1111 ( 
.A(n_986),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1013),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_993),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1044),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_SL g1115 ( 
.A1(n_1008),
.A2(n_417),
.B1(n_382),
.B2(n_385),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1012),
.A2(n_444),
.B1(n_387),
.B2(n_389),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1050),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_969),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_987),
.A2(n_445),
.B1(n_394),
.B2(n_402),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_SL g1120 ( 
.A1(n_984),
.A2(n_572),
.B(n_565),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1055),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_1058),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_1048),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1037),
.A2(n_422),
.B1(n_406),
.B2(n_447),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_995),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1062),
.A2(n_443),
.B1(n_413),
.B2(n_349),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_986),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1051),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_995),
.B(n_572),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1046),
.B(n_572),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1047),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1005),
.A2(n_577),
.B1(n_576),
.B2(n_569),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1020),
.B(n_577),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_960),
.A2(n_577),
.B1(n_576),
.B2(n_569),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1062),
.B(n_569),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1034),
.A2(n_576),
.B1(n_569),
.B2(n_538),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1036),
.B(n_543),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1024),
.Y(n_1140)
);

CKINVDCx6p67_ASAP7_75t_R g1141 ( 
.A(n_998),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_998),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1057),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1045),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1057),
.A2(n_1063),
.B1(n_1038),
.B2(n_1049),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_979),
.A2(n_7),
.B(n_8),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1010),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1049),
.B(n_569),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1024),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1024),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1045),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1063),
.A2(n_1038),
.B1(n_1061),
.B2(n_959),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_982),
.A2(n_576),
.B1(n_569),
.B2(n_543),
.Y(n_1153)
);

INVx5_ASAP7_75t_L g1154 ( 
.A(n_982),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_959),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_958),
.A2(n_576),
.B1(n_569),
.B2(n_543),
.Y(n_1156)
);

BUFx2_ASAP7_75t_SL g1157 ( 
.A(n_991),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1054),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1140),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1146),
.A2(n_957),
.B(n_1061),
.C(n_961),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1149),
.B(n_967),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1150),
.A2(n_1064),
.B(n_1032),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1125),
.B(n_967),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1148),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1114),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1148),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1148),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1128),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1128),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1158),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1155),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1157),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1066),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1145),
.A2(n_1035),
.B(n_1064),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1131),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1152),
.B(n_967),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1074),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1143),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1132),
.B(n_1023),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1108),
.A2(n_576),
.B1(n_973),
.B2(n_976),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1083),
.Y(n_1181)
);

INVxp67_ASAP7_75t_SL g1182 ( 
.A(n_1147),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1142),
.B(n_968),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1141),
.B(n_968),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1093),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1073),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1101),
.B(n_968),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1153),
.A2(n_1031),
.B(n_973),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1154),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1099),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1107),
.B(n_992),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1158),
.B(n_1041),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1100),
.A2(n_996),
.B(n_1029),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1158),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1113),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1098),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1099),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1154),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1154),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1103),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1144),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1069),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1081),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1129),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1146),
.A2(n_1053),
.B1(n_1054),
.B2(n_991),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1088),
.A2(n_1002),
.B(n_1016),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1112),
.B(n_992),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1136),
.A2(n_1022),
.B(n_1014),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1102),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1153),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1137),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1110),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1134),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1130),
.A2(n_1032),
.B(n_1025),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1112),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1110),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1151),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1087),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1121),
.B(n_1017),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1156),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1117),
.B(n_1017),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_978),
.A3(n_1019),
.B(n_1053),
.Y(n_1222)
);

INVxp33_ASAP7_75t_L g1223 ( 
.A(n_1094),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1077),
.B(n_974),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1190),
.B(n_1077),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1217),
.A2(n_1100),
.B1(n_1122),
.B2(n_1071),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1176),
.B(n_1017),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1190),
.B(n_1197),
.Y(n_1228)
);

AO32x2_ASAP7_75t_L g1229 ( 
.A1(n_1205),
.A2(n_1212),
.A3(n_1194),
.B1(n_1106),
.B2(n_1182),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_SL g1230 ( 
.A(n_1199),
.B(n_1095),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1176),
.B(n_1117),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1212),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1186),
.B(n_1111),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1224),
.A2(n_1126),
.B(n_1115),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1165),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1167),
.B(n_1091),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1176),
.B(n_992),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1174),
.A2(n_1120),
.B(n_1018),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1171),
.A2(n_1122),
.B1(n_1118),
.B2(n_1072),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1217),
.B(n_1078),
.Y(n_1241)
);

CKINVDCx8_ASAP7_75t_R g1242 ( 
.A(n_1218),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1161),
.B(n_1040),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1171),
.A2(n_1079),
.B(n_1075),
.C(n_1120),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_1056),
.B(n_1043),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1177),
.B(n_1040),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1177),
.B(n_1040),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1177),
.B(n_1023),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1197),
.B(n_1079),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1215),
.B(n_1067),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1224),
.A2(n_1090),
.B(n_1085),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1161),
.B(n_1207),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1177),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1215),
.B(n_1067),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1165),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1181),
.B(n_1023),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1181),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1217),
.B(n_1089),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1160),
.A2(n_1109),
.B(n_1111),
.C(n_1096),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1165),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1162),
.A2(n_971),
.B(n_1133),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1216),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1164),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1209),
.B(n_1094),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1161),
.B(n_1025),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1165),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1164),
.B(n_1068),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1164),
.B(n_1068),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1181),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_R g1272 ( 
.A(n_1218),
.B(n_1105),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1217),
.A2(n_1116),
.B1(n_1086),
.B2(n_1104),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1181),
.B(n_1082),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1169),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1162),
.A2(n_1139),
.B(n_1138),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1268),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1228),
.B(n_1221),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1268),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1271),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1271),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1253),
.B(n_1207),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1225),
.B(n_1221),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1250),
.B(n_1221),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1236),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1236),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1232),
.B(n_1179),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1256),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1232),
.B(n_1179),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1233),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1256),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1261),
.B(n_1179),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1264),
.B(n_1219),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1253),
.B(n_1163),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1262),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1262),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1274),
.B(n_1219),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1241),
.B(n_1216),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1261),
.B(n_1265),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1238),
.B(n_1179),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1237),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1265),
.B(n_1164),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1254),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1254),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_1163),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1258),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1258),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1274),
.B(n_1219),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1275),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1233),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1275),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1227),
.B(n_1179),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1227),
.B(n_1179),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1275),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1244),
.B(n_1159),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1229),
.B(n_1164),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1235),
.A2(n_1183),
.B1(n_1184),
.B2(n_1178),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1247),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1252),
.A2(n_1183),
.B1(n_1184),
.B2(n_1178),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1244),
.B(n_1159),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1267),
.B(n_1159),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1229),
.B(n_1166),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1247),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1229),
.B(n_1166),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1259),
.B(n_1212),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1249),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1237),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1249),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1257),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1248),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1248),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1226),
.A2(n_1183),
.B1(n_1184),
.B2(n_1178),
.Y(n_1332)
);

OR2x2_ASAP7_75t_SL g1333 ( 
.A(n_1301),
.B(n_1105),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1277),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1316),
.B(n_1229),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1316),
.B(n_1229),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1285),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1277),
.Y(n_1338)
);

AND2x4_ASAP7_75t_SL g1339 ( 
.A(n_1301),
.B(n_1237),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1299),
.Y(n_1340)
);

AND2x2_ASAP7_75t_SL g1341 ( 
.A(n_1301),
.B(n_1234),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1317),
.B(n_1260),
.C(n_1319),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1280),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1280),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1281),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1301),
.A2(n_1160),
.B(n_1188),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1303),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1281),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1279),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1285),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1286),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1322),
.B(n_1231),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1322),
.B(n_1231),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1295),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1303),
.A2(n_1199),
.B(n_1191),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1282),
.B(n_1294),
.Y(n_1356)
);

OAI211xp5_ASAP7_75t_L g1357 ( 
.A1(n_1332),
.A2(n_1240),
.B(n_1245),
.C(n_1242),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1282),
.B(n_1257),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1324),
.B(n_1300),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1240),
.B1(n_1273),
.B2(n_1178),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1304),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1295),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1286),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1324),
.B(n_1231),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1338),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1335),
.B(n_1299),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1334),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1338),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1356),
.B(n_1278),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1361),
.B(n_1325),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1335),
.B(n_1299),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1337),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1361),
.B(n_1283),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1356),
.B(n_1294),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1334),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1336),
.B(n_1327),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1337),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1341),
.B(n_1301),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1336),
.B(n_1327),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1359),
.B(n_1300),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1334),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1359),
.B(n_1312),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1360),
.B(n_1305),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1345),
.Y(n_1385)
);

NAND4xp25_ASAP7_75t_SL g1386 ( 
.A(n_1342),
.B(n_1186),
.C(n_1272),
.D(n_1242),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1352),
.B(n_1312),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1345),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1360),
.B(n_1326),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1345),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1341),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1339),
.B(n_1352),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1353),
.B(n_1365),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1343),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1343),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1351),
.Y(n_1396)
);

NOR2x1_ASAP7_75t_L g1397 ( 
.A(n_1355),
.B(n_1344),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1371),
.Y(n_1398)
);

AOI322xp5_ASAP7_75t_L g1399 ( 
.A1(n_1374),
.A2(n_1341),
.A3(n_1342),
.B1(n_1357),
.B2(n_1284),
.C1(n_1358),
.C2(n_1293),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1391),
.B(n_1340),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1368),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1371),
.B(n_1086),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1374),
.B(n_1347),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1368),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1391),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1392),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1392),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1392),
.B(n_1339),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1392),
.B(n_1340),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1392),
.B(n_1353),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1366),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1366),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1381),
.B(n_1365),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1384),
.B(n_1358),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1384),
.B(n_1362),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1369),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1370),
.B(n_1375),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1381),
.B(n_1339),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1368),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1396),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1370),
.B(n_1349),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1379),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1369),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1379),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1349),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1373),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1394),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1381),
.B(n_1351),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1394),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1395),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1344),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

OAI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1398),
.A2(n_1357),
.B1(n_1346),
.B2(n_1386),
.C(n_1397),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1408),
.B(n_1418),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1401),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1408),
.B(n_1383),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1424),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1408),
.B(n_1418),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1405),
.B(n_1395),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1399),
.B(n_1383),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1378),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1407),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1408),
.B(n_1383),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1411),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1403),
.B(n_1399),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1422),
.B(n_1387),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1401),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1411),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1404),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1412),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1404),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1406),
.B(n_1393),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1407),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1403),
.B(n_1378),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1417),
.B(n_1373),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_SL g1457 ( 
.A(n_1400),
.B(n_1346),
.C(n_1386),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1407),
.B(n_1377),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1412),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1406),
.B(n_1393),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1416),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1457),
.A2(n_1400),
.B1(n_1409),
.B2(n_1406),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1434),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1434),
.B(n_1410),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1445),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1461),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1437),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1446),
.A2(n_1402),
.B(n_1426),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.B(n_1410),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1446),
.A2(n_1427),
.B1(n_1429),
.B2(n_1423),
.C(n_1416),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1445),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1438),
.B(n_1413),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1442),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1440),
.B(n_1413),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1436),
.B(n_1409),
.Y(n_1477)
);

AO21x1_ASAP7_75t_L g1478 ( 
.A1(n_1458),
.A2(n_1419),
.B(n_1404),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1433),
.A2(n_1406),
.B1(n_1124),
.B2(n_1397),
.C(n_1425),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1442),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1419),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1436),
.A2(n_1414),
.B(n_1428),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1449),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1443),
.B(n_1453),
.Y(n_1484)
);

AOI222xp33_ASAP7_75t_L g1485 ( 
.A1(n_1455),
.A2(n_1124),
.B1(n_1425),
.B2(n_1380),
.C1(n_1377),
.C2(n_1421),
.Y(n_1485)
);

OAI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1447),
.A2(n_1414),
.B(n_1423),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1449),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1455),
.B(n_1135),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1443),
.A2(n_1431),
.B(n_1428),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1441),
.A2(n_1456),
.B(n_1454),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1451),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1454),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1456),
.A2(n_1430),
.B(n_1429),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1451),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1468),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1479),
.A2(n_1462),
.B1(n_1463),
.B2(n_1459),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1465),
.B(n_1462),
.Y(n_1498)
);

AOI322xp5_ASAP7_75t_L g1499 ( 
.A1(n_1469),
.A2(n_1380),
.A3(n_1377),
.B1(n_1459),
.B2(n_1463),
.C1(n_1419),
.C2(n_1448),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1471),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1476),
.B(n_1474),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1484),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1488),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1460),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1479),
.A2(n_1444),
.B1(n_1460),
.B2(n_1439),
.Y(n_1505)
);

NAND5xp2_ASAP7_75t_L g1506 ( 
.A(n_1485),
.B(n_1464),
.C(n_1470),
.D(n_1490),
.E(n_1472),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1467),
.Y(n_1507)
);

OA21x2_ASAP7_75t_SL g1508 ( 
.A1(n_1475),
.A2(n_1302),
.B(n_1333),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1477),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1472),
.A2(n_1439),
.B1(n_1448),
.B2(n_1435),
.C(n_1432),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1482),
.A2(n_1333),
.B(n_1380),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1492),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1493),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1432),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1481),
.A2(n_1435),
.B(n_1432),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1473),
.Y(n_1518)
);

AOI211xp5_ASAP7_75t_L g1519 ( 
.A1(n_1478),
.A2(n_1435),
.B(n_1450),
.C(n_1448),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1486),
.A2(n_1494),
.B1(n_1491),
.B2(n_1487),
.C(n_1483),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1494),
.A2(n_1452),
.B(n_1450),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

OAI21xp33_ASAP7_75t_L g1523 ( 
.A1(n_1493),
.A2(n_1452),
.B(n_1450),
.Y(n_1523)
);

NAND4xp25_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1452),
.C(n_1255),
.D(n_1251),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1470),
.A2(n_1430),
.B(n_1420),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1470),
.B(n_1420),
.C(n_1123),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1479),
.A2(n_1237),
.B1(n_1243),
.B2(n_1213),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1465),
.B(n_1393),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1529)
);

AOI322xp5_ASAP7_75t_L g1530 ( 
.A1(n_1472),
.A2(n_1367),
.A3(n_1372),
.B1(n_1390),
.B2(n_1388),
.C1(n_1382),
.C2(n_1385),
.Y(n_1530)
);

AND2x6_ASAP7_75t_L g1531 ( 
.A(n_1475),
.B(n_1135),
.Y(n_1531)
);

OAI211xp5_ASAP7_75t_L g1532 ( 
.A1(n_1470),
.A2(n_1420),
.B(n_1119),
.C(n_1382),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1468),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1468),
.Y(n_1534)
);

OAI211xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1485),
.A2(n_1396),
.B(n_1382),
.C(n_1385),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1479),
.A2(n_1230),
.B(n_1070),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1465),
.B(n_1367),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1505),
.A2(n_1076),
.B1(n_1355),
.B2(n_1092),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1534),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1506),
.A2(n_1376),
.B(n_1388),
.C(n_1385),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1531),
.Y(n_1543)
);

XNOR2xp5_ASAP7_75t_L g1544 ( 
.A(n_1526),
.B(n_1223),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1497),
.A2(n_1290),
.B1(n_1310),
.B2(n_1367),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1496),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1535),
.A2(n_1243),
.B1(n_1213),
.B2(n_1269),
.Y(n_1547)
);

XNOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1501),
.B(n_8),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1509),
.A2(n_1076),
.B1(n_1355),
.B2(n_1123),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1533),
.B(n_1372),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1531),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1531),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1515),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1513),
.B(n_1387),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1504),
.A2(n_1388),
.B(n_1376),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1498),
.B(n_1372),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1507),
.Y(n_1559)
);

AOI21xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1520),
.A2(n_1503),
.B(n_1525),
.Y(n_1560)
);

XOR2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1537),
.Y(n_1561)
);

AOI222xp33_ASAP7_75t_L g1562 ( 
.A1(n_1517),
.A2(n_1193),
.B1(n_1230),
.B2(n_1211),
.C1(n_1220),
.C2(n_1180),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1536),
.A2(n_1390),
.B1(n_1376),
.B2(n_1396),
.C(n_1350),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1530),
.B(n_1499),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1518),
.B(n_1387),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1522),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1529),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1508),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1523),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1512),
.B(n_1396),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1527),
.A2(n_1310),
.B1(n_1290),
.B2(n_1396),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1523),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1521),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1519),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

XNOR2xp5_ASAP7_75t_L g1577 ( 
.A(n_1511),
.B(n_1223),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1530),
.A2(n_1390),
.B(n_1355),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

XNOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1501),
.B(n_9),
.Y(n_1580)
);

XNOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1501),
.B(n_10),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1534),
.Y(n_1582)
);

AOI211xp5_ASAP7_75t_L g1583 ( 
.A1(n_1506),
.A2(n_1193),
.B(n_13),
.C(n_10),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1579),
.Y(n_1584)
);

NOR4xp25_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1350),
.C(n_1363),
.D(n_1354),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1351),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1583),
.B(n_1070),
.C(n_1068),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

NAND4xp75_ASAP7_75t_L g1589 ( 
.A(n_1564),
.B(n_1204),
.C(n_15),
.D(n_11),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1551),
.B(n_1364),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1583),
.A2(n_1191),
.B(n_1364),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1557),
.B(n_1364),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1539),
.B(n_1354),
.Y(n_1593)
);

NAND4xp25_ASAP7_75t_L g1594 ( 
.A(n_1568),
.B(n_1266),
.C(n_1204),
.D(n_1269),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1538),
.A2(n_1348),
.B(n_1363),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1348),
.Y(n_1596)
);

NAND4xp25_ASAP7_75t_L g1597 ( 
.A(n_1560),
.B(n_1269),
.C(n_1270),
.D(n_1194),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1548),
.Y(n_1598)
);

NOR2x1p5_ASAP7_75t_SL g1599 ( 
.A(n_1570),
.B(n_1304),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1582),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1569),
.A2(n_1270),
.B1(n_1302),
.B2(n_1243),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1543),
.B(n_1070),
.Y(n_1602)
);

CKINVDCx14_ASAP7_75t_R g1603 ( 
.A(n_1543),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1567),
.B(n_1576),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1538),
.B(n_1270),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1542),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1573),
.B(n_1313),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1574),
.A2(n_1198),
.B(n_1189),
.C(n_16),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1580),
.B(n_1313),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1581),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1549),
.A2(n_1189),
.B1(n_1198),
.B2(n_1302),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1554),
.B(n_1287),
.Y(n_1612)
);

NAND4xp25_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1194),
.C(n_1196),
.D(n_1209),
.Y(n_1613)
);

NOR3x1_ASAP7_75t_L g1614 ( 
.A(n_1553),
.B(n_1308),
.C(n_1297),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1577),
.A2(n_1182),
.B(n_1196),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1549),
.B(n_1194),
.C(n_1209),
.D(n_1200),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1559),
.B(n_14),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1558),
.B(n_1287),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1566),
.B(n_15),
.Y(n_1620)
);

NAND4xp25_ASAP7_75t_SL g1621 ( 
.A(n_1562),
.B(n_1292),
.C(n_1289),
.D(n_1306),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1565),
.B(n_1289),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1544),
.B(n_1307),
.Y(n_1623)
);

NAND4xp75_ASAP7_75t_L g1624 ( 
.A(n_1571),
.B(n_19),
.C(n_17),
.D(n_18),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1562),
.A2(n_1080),
.B(n_1180),
.Y(n_1625)
);

OAI21xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1578),
.A2(n_1292),
.B(n_1173),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_L g1627 ( 
.A(n_1545),
.B(n_1194),
.C(n_1170),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1545),
.B(n_1318),
.Y(n_1628)
);

NOR3x1_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1330),
.C(n_1318),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1541),
.Y(n_1630)
);

OAI211xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1563),
.A2(n_1209),
.B(n_1200),
.C(n_1211),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1555),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1547),
.Y(n_1633)
);

NOR3x1_ASAP7_75t_L g1634 ( 
.A(n_1569),
.B(n_1331),
.C(n_1330),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1564),
.A2(n_1173),
.B(n_1185),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1564),
.A2(n_1166),
.B1(n_1187),
.B2(n_1189),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1579),
.B(n_1331),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1598),
.B(n_1323),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1610),
.A2(n_17),
.B(n_18),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1630),
.A2(n_1170),
.B1(n_1187),
.B2(n_1166),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1618),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1608),
.A2(n_1198),
.B(n_1189),
.C(n_1185),
.Y(n_1642)
);

NAND4xp25_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1170),
.C(n_1187),
.D(n_1205),
.Y(n_1643)
);

XOR2x2_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1644)
);

NOR4xp25_ASAP7_75t_L g1645 ( 
.A(n_1584),
.B(n_19),
.C(n_22),
.D(n_23),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1588),
.A2(n_22),
.B(n_24),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1603),
.A2(n_1170),
.B1(n_1309),
.B2(n_1311),
.Y(n_1647)
);

OAI211xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1636),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1600),
.Y(n_1649)
);

AOI221x1_ASAP7_75t_L g1650 ( 
.A1(n_1606),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.C(n_29),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_R g1651 ( 
.A(n_1632),
.B(n_28),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1601),
.A2(n_1198),
.B1(n_1170),
.B2(n_1175),
.C(n_1195),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1634),
.B(n_1326),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1624),
.B(n_29),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1626),
.B(n_1201),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1635),
.A2(n_1175),
.B1(n_1288),
.B2(n_1296),
.C(n_1195),
.Y(n_1657)
);

NAND4xp25_ASAP7_75t_L g1658 ( 
.A(n_1597),
.B(n_1633),
.C(n_1586),
.D(n_1607),
.Y(n_1658)
);

OAI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1585),
.A2(n_30),
.B(n_32),
.C(n_34),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1593),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1615),
.A2(n_1595),
.B1(n_1621),
.B2(n_1637),
.C(n_1594),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1620),
.A2(n_30),
.B(n_34),
.C(n_35),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_35),
.C(n_36),
.Y(n_1663)
);

AOI222xp33_ASAP7_75t_L g1664 ( 
.A1(n_1599),
.A2(n_1220),
.B1(n_1210),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1625),
.A2(n_1082),
.B(n_1202),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1605),
.A2(n_1296),
.B1(n_1314),
.B2(n_1329),
.Y(n_1666)
);

NAND4xp25_ASAP7_75t_L g1667 ( 
.A(n_1592),
.B(n_36),
.C(n_37),
.D(n_41),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1609),
.B(n_1328),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1587),
.B(n_1590),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1596),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1617),
.A2(n_1168),
.B1(n_1210),
.B2(n_44),
.C(n_45),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_SL g1672 ( 
.A(n_1625),
.B(n_1139),
.C(n_42),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1611),
.A2(n_1168),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_1673)
);

OAI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1627),
.A2(n_43),
.B(n_48),
.C(n_49),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

XNOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1611),
.B(n_49),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1591),
.A2(n_50),
.B(n_52),
.C(n_54),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1613),
.A2(n_1172),
.B1(n_1321),
.B2(n_1201),
.C(n_1166),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1641),
.Y(n_1679)
);

AO22x2_ASAP7_75t_L g1680 ( 
.A1(n_1650),
.A2(n_1628),
.B1(n_1622),
.B2(n_1619),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1677),
.B(n_1631),
.C(n_1612),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1654),
.B(n_1614),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1675),
.B(n_1638),
.Y(n_1683)
);

AND3x2_ASAP7_75t_L g1684 ( 
.A(n_1645),
.B(n_52),
.C(n_56),
.Y(n_1684)
);

AOI322xp5_ASAP7_75t_L g1685 ( 
.A1(n_1672),
.A2(n_1329),
.A3(n_1328),
.B1(n_1314),
.B2(n_1291),
.C1(n_1172),
.C2(n_1201),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1661),
.A2(n_1172),
.B1(n_1203),
.B2(n_1202),
.C(n_1201),
.Y(n_1686)
);

XOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1676),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1659),
.A2(n_1669),
.B(n_1642),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_R g1689 ( 
.A(n_1649),
.B(n_56),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1667),
.B(n_57),
.Y(n_1690)
);

OAI31xp33_ASAP7_75t_L g1691 ( 
.A1(n_1648),
.A2(n_57),
.A3(n_58),
.B(n_59),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1677),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_1692)
);

OAI21xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1653),
.A2(n_1321),
.B(n_1291),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1674),
.A2(n_61),
.B(n_62),
.C(n_64),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1658),
.A2(n_1172),
.B1(n_1202),
.B2(n_1203),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1667),
.A2(n_1320),
.B1(n_1315),
.B2(n_1169),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1663),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.C(n_67),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1646),
.Y(n_1698)
);

AOI31xp33_ASAP7_75t_L g1699 ( 
.A1(n_1655),
.A2(n_1084),
.A3(n_67),
.B(n_68),
.Y(n_1699)
);

OAI21xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1656),
.A2(n_1320),
.B(n_1315),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1662),
.A2(n_65),
.B(n_69),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1646),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_69),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1639),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C(n_73),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1673),
.A2(n_72),
.B(n_75),
.C(n_76),
.Y(n_1705)
);

OAI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1640),
.A2(n_1203),
.B1(n_1202),
.B2(n_78),
.C(n_79),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1671),
.A2(n_76),
.B(n_77),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_78),
.Y(n_1708)
);

AOI211x1_ASAP7_75t_SL g1709 ( 
.A1(n_1665),
.A2(n_80),
.B(n_82),
.C(n_84),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1678),
.A2(n_1169),
.B1(n_1203),
.B2(n_1192),
.Y(n_1710)
);

AOI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1651),
.A2(n_82),
.B(n_86),
.C(n_576),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1643),
.A2(n_86),
.B1(n_1169),
.B2(n_1188),
.C(n_1276),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1664),
.A2(n_1192),
.B1(n_1159),
.B2(n_1188),
.C(n_1222),
.Y(n_1713)
);

AOI211xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1652),
.A2(n_93),
.B(n_95),
.C(n_97),
.Y(n_1714)
);

NAND4xp25_ASAP7_75t_L g1715 ( 
.A(n_1668),
.B(n_98),
.C(n_99),
.D(n_100),
.Y(n_1715)
);

AOI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1657),
.A2(n_1188),
.B1(n_1276),
.B2(n_1263),
.C(n_111),
.Y(n_1716)
);

OAI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1647),
.A2(n_1239),
.B(n_1214),
.C(n_1162),
.Y(n_1717)
);

AOI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1666),
.A2(n_1174),
.B(n_102),
.C(n_110),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1645),
.A2(n_1188),
.B1(n_1276),
.B2(n_1263),
.C(n_117),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1640),
.A2(n_1192),
.B1(n_1239),
.B2(n_1214),
.Y(n_1720)
);

XNOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1687),
.B(n_101),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1682),
.A2(n_1192),
.B1(n_1263),
.B2(n_1239),
.Y(n_1722)
);

NAND4xp75_ASAP7_75t_L g1723 ( 
.A(n_1708),
.B(n_1683),
.C(n_1690),
.D(n_1702),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1698),
.A2(n_1239),
.B1(n_1246),
.B2(n_122),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1679),
.B(n_1222),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1684),
.B(n_1222),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1698),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1222),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1703),
.Y(n_1731)
);

NAND4xp75_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_112),
.C(n_115),
.D(n_125),
.Y(n_1732)
);

XNOR2xp5_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_126),
.Y(n_1733)
);

OAI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1701),
.A2(n_1192),
.B1(n_1214),
.B2(n_1246),
.C(n_140),
.Y(n_1734)
);

XNOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_1694),
.B(n_130),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1681),
.B(n_1705),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1689),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1691),
.B(n_1222),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_SL g1739 ( 
.A(n_1715),
.B(n_1192),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1707),
.B(n_1222),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_L g1741 ( 
.A(n_1692),
.B(n_543),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1686),
.A2(n_1192),
.B1(n_1246),
.B2(n_1208),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1730),
.C(n_1728),
.D(n_1727),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1723),
.Y(n_1744)
);

OR3x2_ASAP7_75t_L g1745 ( 
.A(n_1731),
.B(n_1711),
.C(n_1699),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1737),
.A2(n_1697),
.B1(n_1704),
.B2(n_1696),
.C(n_1706),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1740),
.B(n_1695),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_1714),
.B(n_1713),
.C(n_1719),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1735),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1733),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1721),
.Y(n_1751)
);

NOR2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1732),
.B(n_1685),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1729),
.A2(n_1712),
.B1(n_1693),
.B2(n_1710),
.C(n_1700),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1744),
.A2(n_1739),
.B1(n_1738),
.B2(n_1734),
.Y(n_1754)
);

AOI222xp33_ASAP7_75t_L g1755 ( 
.A1(n_1750),
.A2(n_1726),
.B1(n_1716),
.B2(n_1720),
.C1(n_1725),
.C2(n_1717),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1745),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1752),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1746),
.A2(n_1724),
.B(n_1718),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1743),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1751),
.B(n_1742),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1749),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1759),
.A2(n_1747),
.B1(n_1753),
.B2(n_1722),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1757),
.Y(n_1763)
);

AO22x2_ASAP7_75t_L g1764 ( 
.A1(n_1761),
.A2(n_1748),
.B1(n_1725),
.B2(n_142),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1756),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1754),
.A2(n_1246),
.B1(n_1208),
.B2(n_1206),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1763),
.B(n_1765),
.Y(n_1767)
);

INVxp33_ASAP7_75t_L g1768 ( 
.A(n_1764),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1762),
.A2(n_1760),
.B1(n_1758),
.B2(n_1755),
.Y(n_1769)
);

AOI22x1_ASAP7_75t_L g1770 ( 
.A1(n_1766),
.A2(n_133),
.B1(n_139),
.B2(n_143),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1765),
.A2(n_1208),
.B1(n_1206),
.B2(n_151),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1767),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1769),
.A2(n_144),
.B1(n_149),
.B2(n_152),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

AO22x2_ASAP7_75t_L g1775 ( 
.A1(n_1770),
.A2(n_155),
.B1(n_160),
.B2(n_168),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1773),
.B(n_1775),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1772),
.Y(n_1777)
);

AO21x2_ASAP7_75t_L g1778 ( 
.A1(n_1772),
.A2(n_1771),
.B(n_170),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1772),
.A2(n_1206),
.B(n_172),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1777),
.A2(n_169),
.B1(n_178),
.B2(n_179),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1777),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1776),
.B(n_193),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1779),
.B(n_1778),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1780),
.B(n_195),
.C(n_200),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1784),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_1783),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_R g1787 ( 
.A1(n_1786),
.A2(n_1781),
.B1(n_203),
.B2(n_206),
.C(n_209),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1785),
.B(n_210),
.C(n_211),
.Y(n_1788)
);


endmodule