module fake_netlist_5_421_n_2635 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2635);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2635;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1587;
wire n_1473;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_809;
wire n_931;
wire n_870;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1400;
wire n_1214;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2332;
wire n_1235;
wire n_703;
wire n_1115;
wire n_980;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_1367;
wire n_928;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_2599;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

INVx2_ASAP7_75t_L g619 ( 
.A(n_596),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_102),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_23),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_73),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_209),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_612),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_377),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_565),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_368),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_124),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_210),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_618),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_137),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_205),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_469),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_326),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_377),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_255),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_508),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_85),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_47),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_561),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_581),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_552),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_564),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_33),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_357),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_583),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_338),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_474),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_549),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_181),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_148),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_137),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_288),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_343),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_93),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_421),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_318),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_322),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_138),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_132),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_111),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_297),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_231),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_492),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_412),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_455),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_502),
.Y(n_668)
);

CKINVDCx16_ASAP7_75t_R g669 ( 
.A(n_82),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_186),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_310),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_73),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_75),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_580),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_533),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_100),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_530),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_107),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_205),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_551),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_491),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_97),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_591),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_128),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_134),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_65),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_485),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_494),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_100),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_576),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_355),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_570),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_454),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_43),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_614),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_281),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_435),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_586),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_239),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_141),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_589),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_396),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_470),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_510),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_300),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_319),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_595),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_29),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_557),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_402),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_127),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_388),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_86),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_256),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_493),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_435),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_507),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_38),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_160),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_555),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_375),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_518),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_346),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_97),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_352),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_19),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_8),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_508),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_215),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_509),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_578),
.Y(n_733)
);

CKINVDCx14_ASAP7_75t_R g734 ( 
.A(n_214),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_340),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_224),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_357),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_471),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_30),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_553),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_75),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_9),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_329),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_143),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_224),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_539),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_247),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_388),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_528),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_538),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_87),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_500),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_517),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_156),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_490),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_484),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_271),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_415),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_414),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_220),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_350),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_498),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_366),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_13),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_365),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_615),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_605),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_515),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_16),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_194),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_534),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_33),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_492),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_443),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_185),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_157),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_32),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_588),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_107),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_126),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_247),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_376),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_475),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_145),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_393),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_474),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_328),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_617),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_353),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_183),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_451),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_468),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_129),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_290),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_206),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_44),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_276),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_503),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_87),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_80),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_426),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_141),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_246),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_285),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_213),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_556),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_287),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_418),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_113),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_63),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_385),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_221),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_82),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_21),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_336),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_558),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_569),
.Y(n_817)
);

BUFx2_ASAP7_75t_SL g818 ( 
.A(n_594),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_603),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_370),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_216),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_270),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_412),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_489),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_68),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_264),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_613),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_45),
.Y(n_828)
);

BUFx10_ASAP7_75t_L g829 ( 
.A(n_15),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_396),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_272),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_577),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_306),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_359),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_191),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_294),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_426),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_347),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_369),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_590),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_352),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_532),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_79),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_81),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_182),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_456),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_434),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_12),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_57),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_58),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_49),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_587),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_122),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_503),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_328),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_450),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_246),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_61),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_488),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_518),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_118),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_842),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_763),
.Y(n_863)
);

INVxp33_ASAP7_75t_L g864 ( 
.A(n_747),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_861),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_763),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_669),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_763),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_763),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_763),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_778),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_763),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_797),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_797),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_797),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_684),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_626),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_684),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_851),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_851),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_851),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_851),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_851),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_851),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_624),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_851),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_649),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_740),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_628),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_628),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_717),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_628),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_631),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_628),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_663),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_675),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_674),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_677),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_663),
.Y(n_900)
);

INVxp33_ASAP7_75t_L g901 ( 
.A(n_625),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_663),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_663),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_717),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_676),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_676),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_693),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_676),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_638),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_676),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_860),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_619),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_635),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_635),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_649),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_637),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_637),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_696),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_699),
.Y(n_919)
);

INVxp33_ASAP7_75t_L g920 ( 
.A(n_629),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_658),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_658),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_659),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_764),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_659),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_717),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_710),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_710),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_721),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_721),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_719),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_722),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_759),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_674),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_638),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_759),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_799),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_733),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_749),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_639),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_799),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_702),
.Y(n_942)
);

INVxp67_ASAP7_75t_SL g943 ( 
.A(n_719),
.Y(n_943)
);

CKINVDCx16_ASAP7_75t_R g944 ( 
.A(n_816),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_809),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_809),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_828),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_829),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_828),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_860),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_750),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_720),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_630),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_720),
.Y(n_954)
);

INVxp33_ASAP7_75t_L g955 ( 
.A(n_633),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_839),
.Y(n_956)
);

INVxp33_ASAP7_75t_L g957 ( 
.A(n_636),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_734),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_839),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_854),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_868),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_890),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_908),
.B(n_619),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_869),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_865),
.A2(n_653),
.B1(n_654),
.B2(n_620),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_874),
.B(n_644),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_890),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_875),
.B(n_644),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_869),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_915),
.B(n_931),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_891),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_912),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_891),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_870),
.A2(n_873),
.B(n_866),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_870),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_895),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_878),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_895),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_873),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_896),
.Y(n_980)
);

NOR2x1_ASAP7_75t_L g981 ( 
.A(n_896),
.B(n_818),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_877),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_912),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_864),
.A2(n_653),
.B1(n_654),
.B2(n_620),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_900),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_894),
.B(n_819),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_912),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_863),
.A2(n_806),
.B(n_788),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_876),
.B(n_641),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_912),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_863),
.A2(n_806),
.B(n_788),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_892),
.A2(n_672),
.B1(n_712),
.B2(n_666),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_912),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_900),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_866),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_897),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_867),
.A2(n_651),
.B(n_645),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_899),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_867),
.Y(n_999)
);

OAI22x1_ASAP7_75t_R g1000 ( 
.A1(n_898),
.A2(n_672),
.B1(n_728),
.B2(n_712),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_907),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_924),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_958),
.B(n_702),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_902),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_871),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_902),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_893),
.B(n_641),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_877),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_903),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_940),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_903),
.B(n_852),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_893),
.B(n_852),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_871),
.A2(n_664),
.B(n_652),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_880),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_SL g1015 ( 
.A(n_879),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_L g1016 ( 
.A(n_905),
.B(n_679),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_880),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_879),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_910),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_881),
.B(n_681),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_910),
.B(n_691),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_881),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_905),
.B(n_642),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_882),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_882),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_972),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_977),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_996),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_964),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_964),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_972),
.Y(n_1031)
);

CKINVDCx8_ASAP7_75t_R g1032 ( 
.A(n_998),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_1001),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_1001),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_1000),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_966),
.B(n_958),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_1000),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_972),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_970),
.B(n_944),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_1003),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_965),
.Y(n_1041)
);

CKINVDCx8_ASAP7_75t_R g1042 ( 
.A(n_961),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_1001),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_964),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_995),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_1024),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_969),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_1001),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_995),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_965),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_986),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_1015),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_989),
.B(n_862),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_1015),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_961),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_984),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_982),
.B(n_911),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_1015),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_982),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_972),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_982),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1008),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1008),
.Y(n_1064)
);

BUFx8_ASAP7_75t_L g1065 ( 
.A(n_970),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_1008),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_995),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_984),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_969),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1019),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1018),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1018),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_989),
.B(n_886),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_972),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_1010),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1019),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1019),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_992),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1012),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_972),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_1020),
.B(n_918),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_992),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1012),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1021),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_1002),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_969),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_983),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1021),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_966),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_966),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_966),
.B(n_889),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_983),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_968),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1021),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_968),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_968),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_968),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_975),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1007),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_999),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1007),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1023),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_983),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_1016),
.B(n_703),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_983),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_1023),
.B(n_919),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_963),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1079),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1073),
.B(n_932),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1056),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_1046),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1058),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1104),
.A2(n_1013),
.B1(n_997),
.B2(n_730),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_1058),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1029),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1027),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1089),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1083),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_1028),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1061),
.Y(n_1120)
);

CKINVDCx6p67_ASAP7_75t_R g1121 ( 
.A(n_1035),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1032),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1029),
.Y(n_1123)
);

INVx6_ASAP7_75t_L g1124 ( 
.A(n_1065),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1102),
.B(n_938),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1099),
.B(n_1101),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1030),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1051),
.Y(n_1128)
);

CKINVDCx16_ASAP7_75t_R g1129 ( 
.A(n_1082),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1039),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1075),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1104),
.A2(n_1013),
.B1(n_997),
.B2(n_730),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1046),
.Y(n_1133)
);

NOR2x1p5_ASAP7_75t_L g1134 ( 
.A(n_1052),
.B(n_872),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1030),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1072),
.B(n_963),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1044),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1044),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1090),
.B(n_1093),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1084),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1047),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1061),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1095),
.B(n_939),
.Y(n_1143)
);

INVx8_ASAP7_75t_L g1144 ( 
.A(n_1060),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_1036),
.B(n_904),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1088),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_1061),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1036),
.B(n_926),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1104),
.A2(n_997),
.B1(n_1013),
.B2(n_657),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_SL g1150 ( 
.A(n_1042),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1091),
.B(n_948),
.Y(n_1151)
);

NOR2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1054),
.B(n_943),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1096),
.B(n_951),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1047),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1069),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1097),
.B(n_1024),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1069),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1107),
.B(n_1024),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1104),
.A2(n_997),
.B1(n_1013),
.B2(n_657),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1094),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1104),
.A2(n_997),
.B1(n_1013),
.B2(n_1020),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1070),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1076),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1085),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1086),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1086),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_R g1167 ( 
.A(n_1053),
.B(n_909),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1077),
.B(n_963),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1046),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1062),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1081),
.A2(n_991),
.B(n_988),
.Y(n_1171)
);

AND3x2_ASAP7_75t_L g1172 ( 
.A(n_1035),
.B(n_731),
.C(n_673),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1026),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1061),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1045),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1033),
.B(n_1024),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1098),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1049),
.Y(n_1178)
);

CKINVDCx6p67_ASAP7_75t_R g1179 ( 
.A(n_1037),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1098),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1055),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1067),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_L g1183 ( 
.A(n_1104),
.B(n_1020),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1063),
.B(n_935),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1100),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1026),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1034),
.A2(n_1043),
.B1(n_1048),
.B2(n_1064),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1026),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1066),
.B(n_952),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1040),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1080),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1071),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1031),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1031),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1059),
.B(n_959),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1080),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1031),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1038),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1038),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1038),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1074),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1103),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1065),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1103),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1106),
.B(n_1024),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1103),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1040),
.B(n_901),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_R g1210 ( 
.A(n_1057),
.B(n_639),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_R g1211 ( 
.A(n_1057),
.B(n_640),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1105),
.B(n_963),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1105),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1105),
.B(n_1020),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1080),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1080),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1087),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1087),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1065),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1087),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1087),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1092),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1092),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1092),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1092),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1078),
.A2(n_709),
.B1(n_746),
.B2(n_647),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1068),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1078),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1041),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1041),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1050),
.B(n_689),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1050),
.B(n_1020),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1037),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1079),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1029),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1126),
.B(n_934),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1117),
.B(n_1136),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1120),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1109),
.B(n_1189),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1209),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1112),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1110),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1112),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1113),
.B(n_999),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1113),
.B(n_999),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1132),
.B(n_1005),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1132),
.B(n_1005),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1149),
.A2(n_974),
.B(n_988),
.Y(n_1248)
);

INVxp33_ASAP7_75t_L g1249 ( 
.A(n_1231),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1108),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1149),
.B(n_1005),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1189),
.B(n_942),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1126),
.B(n_666),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1159),
.B(n_1014),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1159),
.B(n_1014),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1118),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1125),
.B(n_728),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1234),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1125),
.B(n_729),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1187),
.B(n_981),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1130),
.B(n_981),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_L g1262 ( 
.A(n_1226),
.B(n_888),
.C(n_715),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1140),
.B(n_1020),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1146),
.B(n_1020),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1151),
.B(n_888),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1160),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1162),
.Y(n_1267)
);

NOR2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1122),
.B(n_640),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1184),
.B(n_729),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_741),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1136),
.B(n_642),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1151),
.B(n_920),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1163),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1115),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1151),
.B(n_955),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1232),
.A2(n_1020),
.B1(n_711),
.B2(n_767),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1231),
.B(n_741),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1185),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1195),
.B(n_745),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_L g1280 ( 
.A(n_1161),
.B(n_1016),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1123),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_SL g1282 ( 
.A(n_1119),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1195),
.B(n_745),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1114),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1136),
.B(n_1014),
.Y(n_1285)
);

NOR3xp33_ASAP7_75t_L g1286 ( 
.A(n_1129),
.B(n_708),
.C(n_954),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1128),
.B(n_754),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1123),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1128),
.B(n_754),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1127),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1170),
.B(n_643),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1131),
.B(n_761),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_SL g1293 ( 
.A(n_1119),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1175),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1212),
.A2(n_991),
.B(n_974),
.C(n_832),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1192),
.B(n_643),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1164),
.B(n_954),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1168),
.B(n_1017),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1178),
.Y(n_1299)
);

INVxp33_ASAP7_75t_L g1300 ( 
.A(n_1228),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1135),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1212),
.B(n_1181),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1182),
.B(n_1017),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1117),
.B(n_650),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_956),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1143),
.B(n_761),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1135),
.B(n_1022),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1156),
.B(n_1022),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1156),
.B(n_1022),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1137),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1137),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1158),
.B(n_1176),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1138),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1120),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1167),
.B(n_622),
.C(n_621),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_SL g1316 ( 
.A(n_1119),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1138),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1139),
.B(n_650),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1120),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1141),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1227),
.A2(n_957),
.B1(n_834),
.B2(n_836),
.C(n_648),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1158),
.B(n_1025),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1230),
.B(n_956),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_1025),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1207),
.B(n_1025),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1228),
.Y(n_1326)
);

AO221x1_ASAP7_75t_L g1327 ( 
.A1(n_1173),
.A2(n_670),
.B1(n_705),
.B2(n_697),
.C(n_678),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1141),
.Y(n_1328)
);

AO221x1_ASAP7_75t_L g1329 ( 
.A1(n_1173),
.A2(n_707),
.B1(n_739),
.B2(n_735),
.C(n_724),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1139),
.B(n_766),
.Y(n_1330)
);

NOR3xp33_ASAP7_75t_L g1331 ( 
.A(n_1229),
.B(n_960),
.C(n_627),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1152),
.B(n_953),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1207),
.B(n_987),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1154),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1143),
.B(n_822),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1228),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1155),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1186),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1116),
.B(n_960),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1155),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1235),
.B(n_987),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1186),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1157),
.B(n_987),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1157),
.B(n_987),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1235),
.B(n_993),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1165),
.B(n_993),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1166),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1177),
.B(n_993),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1230),
.A2(n_834),
.B1(n_836),
.B2(n_648),
.C(n_646),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1116),
.B(n_771),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1153),
.B(n_817),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1177),
.B(n_993),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1180),
.B(n_990),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1180),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1188),
.B(n_990),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1193),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1153),
.B(n_822),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1188),
.B(n_1204),
.Y(n_1358)
);

NAND2xp33_ASAP7_75t_L g1359 ( 
.A(n_1161),
.B(n_827),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1204),
.B(n_990),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1197),
.B(n_990),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1198),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1144),
.Y(n_1363)
);

NAND2xp33_ASAP7_75t_L g1364 ( 
.A(n_1120),
.B(n_840),
.Y(n_1364)
);

INVxp33_ASAP7_75t_L g1365 ( 
.A(n_1134),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1191),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1198),
.Y(n_1367)
);

AND2x6_ASAP7_75t_SL g1368 ( 
.A(n_1145),
.B(n_742),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1199),
.B(n_975),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1200),
.B(n_962),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1200),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1145),
.B(n_854),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1111),
.B(n_983),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_962),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1215),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1203),
.B(n_967),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1208),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1208),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1145),
.B(n_835),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1148),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1194),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1201),
.B(n_975),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1202),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1148),
.B(n_835),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1206),
.B(n_979),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1191),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1213),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1215),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1144),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1111),
.B(n_1133),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_L g1391 ( 
.A(n_1191),
.B(n_1011),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1217),
.B(n_979),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1111),
.B(n_983),
.Y(n_1393)
);

NOR3xp33_ASAP7_75t_L g1394 ( 
.A(n_1233),
.B(n_632),
.C(n_623),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1144),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1148),
.A2(n_1011),
.B1(n_884),
.B2(n_885),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1218),
.B(n_883),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1218),
.B(n_883),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1220),
.Y(n_1399)
);

INVxp67_ASAP7_75t_L g1400 ( 
.A(n_1210),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1221),
.B(n_885),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1221),
.B(n_1223),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1223),
.B(n_887),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1224),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1191),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1224),
.B(n_887),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1205),
.B(n_829),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1124),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1225),
.B(n_967),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1133),
.B(n_971),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1216),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1222),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1196),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1196),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1150),
.B(n_634),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1133),
.B(n_973),
.Y(n_1416)
);

BUFx2_ASAP7_75t_R g1417 ( 
.A(n_1121),
.Y(n_1417)
);

AO22x2_ASAP7_75t_L g1418 ( 
.A1(n_1380),
.A2(n_1252),
.B1(n_1239),
.B2(n_1400),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1237),
.B(n_1219),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1250),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1422)
);

NAND2x1p5_ASAP7_75t_L g1423 ( 
.A(n_1389),
.B(n_1169),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1256),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1395),
.B(n_1124),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1242),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1279),
.B(n_1124),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1282),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1336),
.B(n_1326),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1283),
.B(n_1179),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1408),
.B(n_1174),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1277),
.A2(n_1259),
.B1(n_1257),
.B2(n_1335),
.C(n_1306),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1363),
.B(n_1174),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1258),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1266),
.Y(n_1435)
);

AO22x2_ASAP7_75t_L g1436 ( 
.A1(n_1262),
.A2(n_1211),
.B1(n_1210),
.B2(n_748),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1278),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1409),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1409),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1238),
.B(n_1174),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1238),
.B(n_1196),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1240),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1313),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1323),
.B(n_1172),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1334),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1337),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1302),
.B(n_1214),
.Y(n_1449)
);

AO22x2_ASAP7_75t_L g1450 ( 
.A1(n_1315),
.A2(n_1211),
.B1(n_751),
.B2(n_753),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1340),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1284),
.B(n_1171),
.Y(n_1452)
);

NAND2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1238),
.B(n_1142),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1357),
.A2(n_841),
.B1(n_843),
.B2(n_838),
.C(n_646),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1347),
.Y(n_1455)
);

OAI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1269),
.A2(n_843),
.B1(n_844),
.B2(n_841),
.C(n_838),
.Y(n_1456)
);

AO22x2_ASAP7_75t_L g1457 ( 
.A1(n_1312),
.A2(n_758),
.B1(n_760),
.B2(n_743),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1267),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1339),
.B(n_1142),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1368),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1300),
.B(n_829),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1273),
.B(n_1171),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1274),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1302),
.B(n_1294),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1281),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1288),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1282),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1372),
.A2(n_768),
.B1(n_772),
.B2(n_765),
.Y(n_1468)
);

AO22x2_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_779),
.B1(n_780),
.B2(n_774),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1290),
.Y(n_1470)
);

AO22x2_ASAP7_75t_L g1471 ( 
.A1(n_1331),
.A2(n_784),
.B1(n_786),
.B2(n_783),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1299),
.B(n_973),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1301),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1311),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1317),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1270),
.A2(n_844),
.B1(n_660),
.B2(n_661),
.C(n_656),
.Y(n_1476)
);

AO22x2_ASAP7_75t_L g1477 ( 
.A1(n_1286),
.A2(n_802),
.B1(n_805),
.B2(n_791),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1272),
.B(n_1150),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1253),
.B(n_662),
.C(n_655),
.Y(n_1479)
);

AO22x2_ASAP7_75t_L g1480 ( 
.A1(n_1260),
.A2(n_820),
.B1(n_824),
.B2(n_814),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1292),
.B(n_665),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1320),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1328),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1321),
.A2(n_671),
.B1(n_680),
.B2(n_668),
.C(n_667),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1236),
.A2(n_1183),
.B1(n_978),
.B2(n_980),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1271),
.A2(n_985),
.B1(n_994),
.B2(n_976),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1303),
.Y(n_1488)
);

OR2x2_ASAP7_75t_SL g1489 ( 
.A(n_1305),
.B(n_845),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1293),
.Y(n_1490)
);

AO22x2_ASAP7_75t_L g1491 ( 
.A1(n_1412),
.A2(n_846),
.B1(n_850),
.B2(n_849),
.Y(n_1491)
);

OR2x2_ASAP7_75t_SL g1492 ( 
.A(n_1287),
.B(n_858),
.Y(n_1492)
);

AO22x2_ASAP7_75t_L g1493 ( 
.A1(n_1379),
.A2(n_837),
.B1(n_945),
.B2(n_941),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1303),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1384),
.A2(n_837),
.B1(n_945),
.B2(n_941),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1397),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1397),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_SL g1498 ( 
.A(n_1332),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1298),
.B(n_985),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1398),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1314),
.B(n_1142),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1275),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1351),
.A2(n_1004),
.B1(n_1006),
.B2(n_994),
.Y(n_1503)
);

AO22x2_ASAP7_75t_L g1504 ( 
.A1(n_1330),
.A2(n_837),
.B1(n_947),
.B2(n_946),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1398),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1265),
.B(n_1142),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1314),
.B(n_1147),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1349),
.A2(n_685),
.B1(n_686),
.B2(n_683),
.C(n_682),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1356),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1401),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1401),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1289),
.B(n_911),
.Y(n_1512)
);

AO22x2_ASAP7_75t_L g1513 ( 
.A1(n_1388),
.A2(n_1399),
.B1(n_1404),
.B2(n_1394),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1403),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1244),
.B(n_1004),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1293),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1350),
.B(n_687),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1403),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1415),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1411),
.Y(n_1521)
);

AO22x2_ASAP7_75t_L g1522 ( 
.A1(n_1244),
.A2(n_914),
.B1(n_916),
.B2(n_913),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1314),
.B(n_1147),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1297),
.B(n_1147),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1245),
.B(n_1006),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1362),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1359),
.A2(n_1009),
.B1(n_690),
.B2(n_692),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1407),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1304),
.A2(n_695),
.B1(n_698),
.B2(n_694),
.C(n_688),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1246),
.B(n_1009),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1291),
.B(n_1296),
.Y(n_1531)
);

BUFx8_ASAP7_75t_L g1532 ( 
.A(n_1316),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1268),
.B(n_949),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1406),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1417),
.Y(n_1535)
);

NAND2x1p5_ASAP7_75t_L g1536 ( 
.A(n_1319),
.B(n_1366),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1406),
.Y(n_1537)
);

AO22x2_ASAP7_75t_L g1538 ( 
.A1(n_1247),
.A2(n_936),
.B1(n_937),
.B2(n_933),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1247),
.B(n_1147),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1251),
.B(n_700),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1377),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1261),
.B(n_701),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1365),
.B(n_704),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1319),
.B(n_906),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1367),
.Y(n_1545)
);

AO22x2_ASAP7_75t_L g1546 ( 
.A1(n_1251),
.A2(n_914),
.B1(n_916),
.B2(n_913),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1254),
.B(n_706),
.Y(n_1547)
);

BUFx8_ASAP7_75t_L g1548 ( 
.A(n_1316),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_L g1549 ( 
.A(n_1319),
.B(n_713),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1371),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1381),
.B(n_917),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1254),
.B(n_714),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1378),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1327),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1280),
.A2(n_718),
.B1(n_723),
.B2(n_716),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1396),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1370),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1374),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1376),
.Y(n_1559)
);

AO22x2_ASAP7_75t_L g1560 ( 
.A1(n_1255),
.A2(n_929),
.B1(n_930),
.B2(n_928),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1366),
.B(n_725),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1285),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1387),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_L g1564 ( 
.A(n_1386),
.B(n_726),
.Y(n_1564)
);

AO22x2_ASAP7_75t_L g1565 ( 
.A1(n_1255),
.A2(n_947),
.B1(n_950),
.B2(n_946),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1383),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1382),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1382),
.Y(n_1568)
);

OAI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1276),
.A2(n_736),
.B1(n_737),
.B2(n_732),
.C(n_727),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1385),
.Y(n_1570)
);

AO22x2_ASAP7_75t_L g1571 ( 
.A1(n_1248),
.A2(n_922),
.B1(n_923),
.B2(n_921),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1329),
.A2(n_744),
.B1(n_752),
.B2(n_738),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1386),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1413),
.A2(n_776),
.B1(n_792),
.B2(n_755),
.Y(n_1574)
);

AO22x2_ASAP7_75t_L g1575 ( 
.A1(n_1248),
.A2(n_927),
.B1(n_928),
.B2(n_925),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1308),
.A2(n_762),
.B1(n_769),
.B2(n_757),
.C(n_756),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1385),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1369),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1410),
.B(n_770),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1338),
.B(n_522),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1338),
.B(n_921),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1386),
.Y(n_1582)
);

NOR2xp67_ASAP7_75t_L g1583 ( 
.A(n_1342),
.B(n_523),
.Y(n_1583)
);

AO22x2_ASAP7_75t_L g1584 ( 
.A1(n_1402),
.A2(n_929),
.B1(n_930),
.B2(n_922),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1307),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1402),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1392),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1392),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1342),
.A2(n_794),
.B1(n_807),
.B2(n_777),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1405),
.Y(n_1590)
);

INVx3_ASAP7_75t_R g1591 ( 
.A(n_1364),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1358),
.A2(n_796),
.B1(n_811),
.B2(n_781),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1375),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1405),
.B(n_950),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1375),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1405),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1410),
.A2(n_775),
.B1(n_782),
.B2(n_773),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1416),
.B(n_785),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1420),
.Y(n_1599)
);

O2A1O1Ixp5_ASAP7_75t_L g1600 ( 
.A1(n_1481),
.A2(n_1393),
.B(n_1295),
.C(n_1325),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1432),
.B(n_1502),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1427),
.B(n_1416),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1582),
.Y(n_1603)
);

O2A1O1Ixp5_ASAP7_75t_L g1604 ( 
.A1(n_1561),
.A2(n_1333),
.B(n_1324),
.C(n_1390),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1421),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1479),
.A2(n_1263),
.B(n_1264),
.C(n_1309),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1449),
.A2(n_1322),
.B(n_1355),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1464),
.A2(n_1360),
.B(n_1391),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1424),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1512),
.B(n_1430),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1443),
.B(n_1341),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1438),
.B(n_1353),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1439),
.B(n_1361),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1426),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1421),
.Y(n_1615)
);

OAI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1456),
.A2(n_789),
.B(n_787),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1499),
.A2(n_1373),
.B(n_1414),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1496),
.A2(n_1414),
.B(n_1344),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1557),
.B(n_1558),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1497),
.A2(n_1505),
.B(n_1500),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1559),
.B(n_1343),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1531),
.A2(n_1346),
.B(n_1348),
.C(n_1345),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1434),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1556),
.B(n_1352),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1435),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1454),
.A2(n_793),
.B(n_795),
.C(n_790),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1445),
.B(n_798),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1458),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1441),
.Y(n_1629)
);

AOI33xp33_ASAP7_75t_L g1630 ( 
.A1(n_1572),
.A2(n_804),
.A3(n_801),
.B1(n_808),
.B2(n_803),
.B3(n_800),
.Y(n_1630)
);

BUFx4f_ASAP7_75t_L g1631 ( 
.A(n_1425),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1590),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1510),
.A2(n_525),
.B(n_524),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1476),
.A2(n_812),
.B(n_813),
.C(n_810),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1511),
.A2(n_821),
.B1(n_823),
.B2(n_815),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1488),
.B(n_825),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1514),
.A2(n_1534),
.B(n_1518),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1494),
.B(n_826),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1586),
.B(n_830),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1537),
.A2(n_527),
.B(n_526),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1528),
.B(n_831),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1517),
.A2(n_847),
.B(n_848),
.C(n_833),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1562),
.B(n_853),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1542),
.A2(n_856),
.B(n_857),
.C(n_855),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1532),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1579),
.B(n_1598),
.Y(n_1646)
);

AOI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1515),
.A2(n_531),
.B(n_529),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1429),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1485),
.A2(n_859),
.B(n_2),
.C(n_0),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1444),
.Y(n_1650)
);

CKINVDCx10_ASAP7_75t_R g1651 ( 
.A(n_1498),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1539),
.A2(n_536),
.B(n_535),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1525),
.A2(n_540),
.B(n_537),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1530),
.A2(n_542),
.B(n_541),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1563),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1501),
.A2(n_544),
.B(n_543),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1436),
.B(n_1),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1543),
.B(n_1),
.C(n_2),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1585),
.A2(n_546),
.B(n_545),
.Y(n_1659)
);

AO22x1_ASAP7_75t_L g1660 ( 
.A1(n_1428),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1567),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1540),
.B(n_6),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1568),
.A2(n_548),
.B(n_547),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1576),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1425),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1446),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1447),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1467),
.B(n_7),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1570),
.A2(n_554),
.B(n_550),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1577),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1436),
.B(n_10),
.Y(n_1671)
);

AO21x1_ASAP7_75t_L g1672 ( 
.A1(n_1452),
.A2(n_1462),
.B(n_1547),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1461),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1554),
.A2(n_1450),
.B1(n_1480),
.B2(n_1418),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1429),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1480),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1578),
.A2(n_1588),
.B(n_1587),
.Y(n_1677)
);

AO22x2_ASAP7_75t_L g1678 ( 
.A1(n_1493),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1529),
.A2(n_18),
.B(n_14),
.C(n_17),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1418),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1680)
);

BUFx2_ASAP7_75t_SL g1681 ( 
.A(n_1520),
.Y(n_1681)
);

AO21x1_ASAP7_75t_L g1682 ( 
.A1(n_1452),
.A2(n_22),
.B(n_21),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1508),
.A2(n_20),
.B(n_22),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1486),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1451),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1450),
.B(n_24),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1581),
.B(n_1448),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1573),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1492),
.B(n_25),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1552),
.B(n_26),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1489),
.B(n_27),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1571),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1422),
.A2(n_560),
.B(n_559),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1437),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1581),
.B(n_31),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1459),
.A2(n_563),
.B(n_562),
.Y(n_1696)
);

INVx11_ASAP7_75t_L g1697 ( 
.A(n_1548),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1575),
.A2(n_567),
.B(n_566),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1566),
.B(n_34),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1575),
.A2(n_571),
.B(n_568),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1478),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1580),
.A2(n_573),
.B(n_572),
.Y(n_1702)
);

OA22x2_ASAP7_75t_L g1703 ( 
.A1(n_1555),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1506),
.B(n_37),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1583),
.A2(n_575),
.B(n_574),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1536),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1455),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1472),
.A2(n_1519),
.B(n_1550),
.C(n_1545),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1553),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1506),
.B(n_38),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1468),
.B(n_39),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1419),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1551),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1521),
.B(n_40),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1469),
.B(n_41),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1503),
.A2(n_584),
.B(n_582),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1592),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1524),
.B(n_46),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1522),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1719)
);

CKINVDCx11_ASAP7_75t_R g1720 ( 
.A(n_1460),
.Y(n_1720)
);

AO21x1_ASAP7_75t_L g1721 ( 
.A1(n_1595),
.A2(n_48),
.B(n_50),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1524),
.B(n_50),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1596),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1597),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1442),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1487),
.A2(n_616),
.B(n_592),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1469),
.B(n_51),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1431),
.B(n_1593),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1431),
.B(n_585),
.Y(n_1729)
);

CKINVDCx10_ASAP7_75t_R g1730 ( 
.A(n_1478),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1440),
.A2(n_597),
.B(n_593),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1549),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1513),
.A2(n_599),
.B(n_598),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1504),
.B(n_54),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1513),
.A2(n_601),
.B(n_600),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1589),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1736)
);

O2A1O1Ixp5_ASAP7_75t_L g1737 ( 
.A1(n_1463),
.A2(n_1465),
.B(n_1470),
.C(n_1466),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1473),
.B(n_1474),
.Y(n_1738)
);

AO22x1_ASAP7_75t_L g1739 ( 
.A1(n_1490),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1475),
.B(n_1482),
.Y(n_1740)
);

NOR2xp67_ASAP7_75t_L g1741 ( 
.A(n_1535),
.B(n_604),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1453),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1483),
.B(n_59),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1574),
.B(n_60),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1569),
.B(n_60),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1527),
.A2(n_1484),
.B(n_1526),
.C(n_1509),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1541),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1584),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1433),
.B(n_62),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1584),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1544),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1564),
.B(n_62),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1538),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1591),
.B(n_63),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1457),
.B(n_64),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1457),
.B(n_65),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1468),
.B(n_66),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1471),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1507),
.A2(n_607),
.B(n_606),
.Y(n_1759)
);

BUFx4f_ASAP7_75t_SL g1760 ( 
.A(n_1516),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1546),
.A2(n_609),
.B(n_608),
.Y(n_1761)
);

AO21x1_ASAP7_75t_L g1762 ( 
.A1(n_1594),
.A2(n_67),
.B(n_69),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_SL g1763 ( 
.A(n_1423),
.B(n_1523),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1631),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1610),
.B(n_1495),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1634),
.A2(n_1471),
.B(n_1495),
.C(n_1477),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1602),
.A2(n_1477),
.B1(n_1491),
.B2(n_1533),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1631),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1619),
.B(n_1491),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1608),
.A2(n_1560),
.B(n_1546),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1648),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1607),
.A2(n_1565),
.B(n_1560),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1681),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1624),
.B(n_610),
.Y(n_1774)
);

OAI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1745),
.A2(n_70),
.B(n_71),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_R g1776 ( 
.A(n_1760),
.B(n_611),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1658),
.B(n_70),
.C(n_71),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1646),
.B(n_72),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1675),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1618),
.A2(n_74),
.B(n_76),
.Y(n_1780)
);

BUFx10_ASAP7_75t_L g1781 ( 
.A(n_1665),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1601),
.B(n_74),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1605),
.B(n_76),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1625),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1673),
.B(n_77),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1603),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1605),
.B(n_77),
.Y(n_1787)
);

A2O1A1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1626),
.A2(n_1716),
.B(n_1726),
.C(n_1649),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_SL g1789 ( 
.A(n_1645),
.B(n_78),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1723),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1733),
.A2(n_78),
.B(n_80),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1655),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1620),
.A2(n_521),
.B(n_81),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1611),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1665),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1683),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1796)
);

AO21x1_ASAP7_75t_L g1797 ( 
.A1(n_1680),
.A2(n_83),
.B(n_84),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1735),
.A2(n_86),
.B(n_88),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1639),
.B(n_88),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1665),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1614),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1632),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1636),
.B(n_89),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1695),
.B(n_89),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1637),
.A2(n_90),
.B(n_91),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1603),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1599),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1603),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1612),
.A2(n_90),
.B(n_91),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1662),
.B(n_92),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1690),
.B(n_92),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1613),
.A2(n_521),
.B(n_93),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1651),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1600),
.A2(n_94),
.B(n_95),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1674),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_SL g1816 ( 
.A(n_1716),
.B(n_96),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1730),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1708),
.A2(n_1744),
.B1(n_1713),
.B2(n_1638),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1752),
.B(n_98),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1643),
.A2(n_101),
.B1(n_98),
.B2(n_99),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1687),
.B(n_99),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_1720),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1609),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1725),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1621),
.B(n_103),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1717),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1736),
.A2(n_108),
.B1(n_105),
.B2(n_106),
.Y(n_1827)
);

INVx6_ASAP7_75t_L g1828 ( 
.A(n_1701),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_SL g1829 ( 
.A(n_1668),
.B(n_106),
.C(n_108),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1630),
.B(n_109),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1718),
.B(n_1722),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1689),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_1832)
);

A2O1A1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1726),
.A2(n_113),
.B(n_110),
.C(n_112),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1615),
.B(n_114),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1615),
.B(n_1672),
.Y(n_1835)
);

O2A1O1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1758),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1677),
.B(n_116),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1699),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1714),
.B(n_117),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1704),
.B(n_119),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1617),
.A2(n_520),
.B(n_119),
.Y(n_1841)
);

INVx5_ASAP7_75t_L g1842 ( 
.A(n_1725),
.Y(n_1842)
);

NOR2xp67_ASAP7_75t_SL g1843 ( 
.A(n_1653),
.B(n_120),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1606),
.A2(n_120),
.B(n_121),
.Y(n_1844)
);

NOR3xp33_ASAP7_75t_SL g1845 ( 
.A(n_1680),
.B(n_121),
.C(n_122),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1623),
.B(n_123),
.Y(n_1846)
);

BUFx4f_ASAP7_75t_L g1847 ( 
.A(n_1725),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1753),
.B(n_123),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1628),
.Y(n_1849)
);

INVx6_ASAP7_75t_L g1850 ( 
.A(n_1706),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1653),
.A2(n_124),
.B(n_125),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1622),
.A2(n_520),
.B(n_125),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1747),
.B(n_126),
.Y(n_1853)
);

CKINVDCx10_ASAP7_75t_R g1854 ( 
.A(n_1697),
.Y(n_1854)
);

O2A1O1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1664),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_1855)
);

O2A1O1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1679),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1732),
.A2(n_133),
.B(n_130),
.C(n_131),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1710),
.B(n_133),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1629),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1604),
.A2(n_519),
.B(n_134),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1650),
.B(n_135),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1688),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1627),
.B(n_135),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1641),
.B(n_1616),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1666),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1654),
.A2(n_519),
.B(n_136),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1667),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_SL g1868 ( 
.A(n_1734),
.B(n_136),
.C(n_138),
.Y(n_1868)
);

O2A1O1Ixp5_ASAP7_75t_L g1869 ( 
.A1(n_1698),
.A2(n_142),
.B(n_139),
.C(n_140),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1685),
.B(n_139),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1702),
.A2(n_516),
.B(n_142),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1706),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1707),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1729),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1642),
.A2(n_143),
.B(n_144),
.Y(n_1875)
);

A2O1A1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1724),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1705),
.A2(n_516),
.B(n_146),
.Y(n_1877)
);

OR2x2_ASAP7_75t_SL g1878 ( 
.A(n_1715),
.B(n_147),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1729),
.B(n_147),
.Y(n_1879)
);

NAND2xp33_ASAP7_75t_R g1880 ( 
.A(n_1742),
.B(n_148),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1749),
.B(n_1644),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1742),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1754),
.B(n_149),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1691),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1709),
.B(n_152),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1738),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1740),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1656),
.A2(n_156),
.B(n_157),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1635),
.B(n_158),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1737),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1743),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1746),
.A2(n_158),
.B(n_159),
.Y(n_1892)
);

NAND2xp33_ASAP7_75t_R g1893 ( 
.A(n_1751),
.B(n_159),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_SL g1894 ( 
.A(n_1668),
.B(n_160),
.C(n_161),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1741),
.B(n_161),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1763),
.B(n_162),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1711),
.B(n_162),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1750),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1748),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1728),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_R g1901 ( 
.A(n_1647),
.B(n_166),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1757),
.B(n_166),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1759),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1712),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1652),
.A2(n_515),
.B(n_167),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1703),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1663),
.A2(n_514),
.B(n_168),
.Y(n_1907)
);

CKINVDCx6p67_ASAP7_75t_R g1908 ( 
.A(n_1755),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1727),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1788),
.A2(n_1684),
.B(n_1700),
.Y(n_1910)
);

AO31x2_ASAP7_75t_L g1911 ( 
.A1(n_1772),
.A2(n_1682),
.A3(n_1692),
.B(n_1721),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1794),
.B(n_1686),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1833),
.A2(n_1703),
.B(n_1692),
.Y(n_1913)
);

AO31x2_ASAP7_75t_L g1914 ( 
.A1(n_1770),
.A2(n_1890),
.A3(n_1851),
.B(n_1903),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1771),
.Y(n_1915)
);

OAI21xp33_ASAP7_75t_L g1916 ( 
.A1(n_1816),
.A2(n_1678),
.B(n_1756),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1891),
.B(n_1657),
.Y(n_1917)
);

AOI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1843),
.A2(n_1852),
.B(n_1892),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1779),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1818),
.B(n_1864),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1775),
.A2(n_1676),
.B(n_1719),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1769),
.B(n_1671),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1859),
.Y(n_1923)
);

NOR2xp67_ASAP7_75t_L g1924 ( 
.A(n_1802),
.B(n_1693),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1867),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1844),
.A2(n_1640),
.B(n_1633),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1814),
.A2(n_1669),
.B(n_1659),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1899),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1854),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1806),
.Y(n_1930)
);

OAI22x1_ASAP7_75t_L g1931 ( 
.A1(n_1884),
.A2(n_1660),
.B1(n_1739),
.B2(n_1676),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1874),
.B(n_1761),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1807),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1838),
.B(n_1661),
.Y(n_1934)
);

OA21x2_ASAP7_75t_L g1935 ( 
.A1(n_1869),
.A2(n_1860),
.B(n_1780),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1835),
.A2(n_1731),
.B(n_1696),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1909),
.B(n_1762),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1841),
.A2(n_1670),
.B(n_1694),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1907),
.A2(n_169),
.B(n_170),
.Y(n_1939)
);

AOI211x1_ASAP7_75t_L g1940 ( 
.A1(n_1775),
.A2(n_1826),
.B(n_1819),
.C(n_1827),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1909),
.B(n_514),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1768),
.Y(n_1942)
);

AO31x2_ASAP7_75t_L g1943 ( 
.A1(n_1797),
.A2(n_172),
.A3(n_170),
.B(n_171),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1875),
.A2(n_171),
.B(n_172),
.Y(n_1944)
);

AOI21x1_ASAP7_75t_SL g1945 ( 
.A1(n_1782),
.A2(n_1889),
.B(n_1837),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1823),
.Y(n_1946)
);

AO22x1_ASAP7_75t_L g1947 ( 
.A1(n_1883),
.A2(n_1863),
.B1(n_1858),
.B2(n_1840),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1808),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1888),
.A2(n_173),
.B(n_174),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1849),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1866),
.A2(n_173),
.B(n_174),
.Y(n_1951)
);

NAND3x1_ASAP7_75t_L g1952 ( 
.A(n_1884),
.B(n_175),
.C(n_176),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1905),
.A2(n_1805),
.B(n_1793),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1881),
.B(n_175),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1909),
.B(n_176),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1790),
.Y(n_1956)
);

BUFx2_ASAP7_75t_L g1957 ( 
.A(n_1795),
.Y(n_1957)
);

AO22x2_ASAP7_75t_L g1958 ( 
.A1(n_1815),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1824),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1865),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1801),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_SL g1962 ( 
.A1(n_1857),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_1962)
);

OAI21xp33_ASAP7_75t_L g1963 ( 
.A1(n_1845),
.A2(n_180),
.B(n_181),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1856),
.A2(n_180),
.B(n_182),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1855),
.A2(n_183),
.B(n_184),
.Y(n_1965)
);

AO31x2_ASAP7_75t_L g1966 ( 
.A1(n_1766),
.A2(n_186),
.A3(n_184),
.B(n_185),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1795),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1876),
.A2(n_187),
.B(n_188),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1871),
.A2(n_187),
.B(n_188),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1804),
.B(n_189),
.Y(n_1970)
);

BUFx2_ASAP7_75t_L g1971 ( 
.A(n_1795),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_SL g1972 ( 
.A(n_1832),
.B(n_189),
.C(n_190),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1877),
.A2(n_192),
.B(n_193),
.Y(n_1973)
);

NOR2xp67_ASAP7_75t_L g1974 ( 
.A(n_1764),
.B(n_193),
.Y(n_1974)
);

AO21x2_ASAP7_75t_L g1975 ( 
.A1(n_1901),
.A2(n_194),
.B(n_195),
.Y(n_1975)
);

NOR4xp25_ASAP7_75t_L g1976 ( 
.A(n_1777),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_1976)
);

BUFx12f_ASAP7_75t_L g1977 ( 
.A(n_1813),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1908),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_1978)
);

OAI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1791),
.A2(n_198),
.B(n_199),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1778),
.B(n_513),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1796),
.A2(n_199),
.B(n_200),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1874),
.B(n_200),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1825),
.B(n_513),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1791),
.A2(n_201),
.B(n_202),
.Y(n_1984)
);

OA22x2_ASAP7_75t_L g1985 ( 
.A1(n_1848),
.A2(n_1879),
.B1(n_1765),
.B2(n_1767),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_R g1986 ( 
.A(n_1854),
.B(n_201),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1768),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1798),
.A2(n_203),
.B(n_204),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1784),
.B(n_512),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1773),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1836),
.A2(n_207),
.B(n_208),
.Y(n_1991)
);

NAND2x1_ASAP7_75t_L g1992 ( 
.A(n_1900),
.B(n_208),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1774),
.B(n_209),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1906),
.B(n_210),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1768),
.Y(n_1995)
);

AOI211x1_ASAP7_75t_L g1996 ( 
.A1(n_1829),
.A2(n_1894),
.B(n_1902),
.C(n_1897),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1831),
.B(n_512),
.Y(n_1997)
);

A2O1A1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1809),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1812),
.A2(n_211),
.B(n_212),
.Y(n_1999)
);

BUFx12f_ASAP7_75t_L g2000 ( 
.A(n_1781),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1904),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.C(n_217),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1800),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1895),
.A2(n_217),
.B(n_218),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1792),
.B(n_511),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1873),
.B(n_218),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1928),
.Y(n_2006)
);

OAI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1944),
.A2(n_1820),
.B(n_1811),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1933),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1912),
.B(n_1868),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1946),
.B(n_1848),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1923),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1927),
.A2(n_1830),
.B(n_1803),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1920),
.A2(n_1810),
.B1(n_1887),
.B2(n_1886),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1961),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1925),
.B(n_1878),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1916),
.A2(n_1968),
.B(n_1969),
.C(n_1963),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1950),
.Y(n_2017)
);

OAI22x1_ASAP7_75t_SL g2018 ( 
.A1(n_1929),
.A2(n_1822),
.B1(n_1817),
.B2(n_1893),
.Y(n_2018)
);

OA21x2_ASAP7_75t_L g2019 ( 
.A1(n_1984),
.A2(n_1861),
.B(n_1846),
.Y(n_2019)
);

OAI21x1_ASAP7_75t_SL g2020 ( 
.A1(n_1964),
.A2(n_1898),
.B(n_1885),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1932),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1967),
.Y(n_2022)
);

NAND2x1p5_ASAP7_75t_L g2023 ( 
.A(n_1932),
.B(n_1956),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1960),
.Y(n_2024)
);

NAND2x1_ASAP7_75t_L g2025 ( 
.A(n_1921),
.B(n_1850),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1922),
.B(n_1848),
.Y(n_2026)
);

OAI21x1_ASAP7_75t_L g2027 ( 
.A1(n_1936),
.A2(n_1853),
.B(n_1870),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1926),
.A2(n_1834),
.B(n_1896),
.Y(n_2028)
);

AO21x2_ASAP7_75t_L g2029 ( 
.A1(n_1910),
.A2(n_1839),
.B(n_1799),
.Y(n_2029)
);

OA21x2_ASAP7_75t_L g2030 ( 
.A1(n_1979),
.A2(n_1988),
.B(n_1938),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1914),
.B(n_1821),
.Y(n_2031)
);

AOI332xp33_ASAP7_75t_L g2032 ( 
.A1(n_1978),
.A2(n_1880),
.A3(n_220),
.B1(n_221),
.B2(n_222),
.B3(n_223),
.C1(n_225),
.C2(n_226),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1919),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1977),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1918),
.A2(n_1785),
.B(n_1842),
.Y(n_2035)
);

INVx6_ASAP7_75t_L g2036 ( 
.A(n_1942),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1937),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_SL g2038 ( 
.A(n_1975),
.B(n_1842),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1972),
.A2(n_1789),
.B1(n_1783),
.B2(n_1787),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1935),
.A2(n_1953),
.B(n_1939),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1914),
.Y(n_2041)
);

BUFx12f_ASAP7_75t_L g2042 ( 
.A(n_2000),
.Y(n_2042)
);

NAND2x1p5_ASAP7_75t_L g2043 ( 
.A(n_1953),
.B(n_1842),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1914),
.B(n_1824),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1917),
.B(n_1947),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1990),
.B(n_1828),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1915),
.B(n_1783),
.Y(n_2047)
);

OAI21x1_ASAP7_75t_L g2048 ( 
.A1(n_1935),
.A2(n_1847),
.B(n_1781),
.Y(n_2048)
);

OA21x2_ASAP7_75t_L g2049 ( 
.A1(n_1949),
.A2(n_1862),
.B(n_1786),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1966),
.B(n_1800),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1951),
.A2(n_219),
.B(n_222),
.Y(n_2051)
);

INVx5_ASAP7_75t_L g2052 ( 
.A(n_2002),
.Y(n_2052)
);

INVx2_ASAP7_75t_SL g2053 ( 
.A(n_2002),
.Y(n_2053)
);

AO31x2_ASAP7_75t_L g2054 ( 
.A1(n_1931),
.A2(n_225),
.A3(n_219),
.B(n_223),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1993),
.A2(n_1828),
.B1(n_1847),
.B2(n_1850),
.Y(n_2055)
);

INVx6_ASAP7_75t_L g2056 ( 
.A(n_1942),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1940),
.A2(n_1800),
.B1(n_1882),
.B2(n_1872),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1966),
.Y(n_2058)
);

A2O1A1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_1965),
.A2(n_1776),
.B(n_1872),
.C(n_1824),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1973),
.A2(n_1872),
.B(n_226),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_1948),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1966),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1911),
.B(n_1985),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2006),
.Y(n_2064)
);

OAI21x1_ASAP7_75t_L g2065 ( 
.A1(n_2040),
.A2(n_1999),
.B(n_1945),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_2021),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_2058),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2008),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_2030),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_2050),
.Y(n_2070)
);

OAI22xp33_ASAP7_75t_SL g2071 ( 
.A1(n_2045),
.A2(n_1954),
.B1(n_1934),
.B2(n_1997),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2062),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_2034),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_2021),
.B(n_1957),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_2050),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_2007),
.A2(n_1981),
.B1(n_1958),
.B2(n_2003),
.Y(n_2076)
);

INVx4_ASAP7_75t_L g2077 ( 
.A(n_2052),
.Y(n_2077)
);

AO21x1_ASAP7_75t_L g2078 ( 
.A1(n_2012),
.A2(n_1980),
.B(n_1983),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_2021),
.Y(n_2079)
);

AO21x2_ASAP7_75t_L g2080 ( 
.A1(n_2040),
.A2(n_1913),
.B(n_1991),
.Y(n_2080)
);

BUFx3_ASAP7_75t_L g2081 ( 
.A(n_2023),
.Y(n_2081)
);

AOI21x1_ASAP7_75t_L g2082 ( 
.A1(n_2041),
.A2(n_1924),
.B(n_1941),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2017),
.Y(n_2083)
);

AOI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_2020),
.A2(n_1958),
.B1(n_1955),
.B2(n_1970),
.Y(n_2084)
);

AOI21xp33_ASAP7_75t_L g2085 ( 
.A1(n_2016),
.A2(n_2001),
.B(n_1952),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_2023),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2011),
.B(n_1943),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_2044),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_2034),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2013),
.A2(n_1994),
.B1(n_2005),
.B2(n_1986),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2024),
.Y(n_2091)
);

OAI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2032),
.A2(n_1974),
.B1(n_1976),
.B2(n_1992),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_2081),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2078),
.A2(n_2016),
.B(n_2059),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2064),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_2079),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2076),
.A2(n_2059),
.B1(n_2039),
.B2(n_2025),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2064),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2064),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_L g2100 ( 
.A1(n_2092),
.A2(n_1998),
.B(n_1962),
.C(n_2009),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2085),
.A2(n_2029),
.B1(n_2063),
.B2(n_2019),
.Y(n_2101)
);

BUFx4f_ASAP7_75t_SL g2102 ( 
.A(n_2089),
.Y(n_2102)
);

BUFx4f_ASAP7_75t_SL g2103 ( 
.A(n_2089),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2078),
.B(n_2033),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2085),
.A2(n_2029),
.B1(n_2063),
.B2(n_2019),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2064),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2076),
.A2(n_2029),
.B1(n_2019),
.B2(n_2026),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2068),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2084),
.A2(n_1996),
.B1(n_2055),
.B2(n_2015),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2070),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2068),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_2078),
.A2(n_2026),
.B1(n_2051),
.B2(n_2028),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2092),
.A2(n_2051),
.B1(n_2028),
.B2(n_2037),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_R g2114 ( 
.A(n_2102),
.B(n_2073),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_2104),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2110),
.B(n_2070),
.Y(n_2116)
);

OR2x6_ASAP7_75t_L g2117 ( 
.A(n_2094),
.B(n_2077),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_2103),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2108),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_2109),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_R g2121 ( 
.A(n_2096),
.B(n_2070),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2110),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_2113),
.B(n_2042),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_2093),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2116),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2124),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2119),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2117),
.B(n_2093),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2124),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2117),
.B(n_2093),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2125),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2125),
.B(n_2115),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2128),
.B(n_2130),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2130),
.B(n_2117),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2126),
.B(n_2120),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2129),
.B(n_2117),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2127),
.B(n_2117),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2126),
.A2(n_2123),
.B1(n_2097),
.B2(n_2107),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_2130),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2134),
.B(n_2116),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2132),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2131),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2134),
.B(n_2140),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2136),
.B(n_2015),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2131),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2133),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2140),
.B(n_2139),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2138),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2138),
.B(n_2100),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2137),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_2144),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_2144),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2141),
.B(n_2137),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_2147),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2148),
.A2(n_2135),
.B1(n_2080),
.B2(n_2105),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2141),
.B(n_2135),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2143),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2146),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2145),
.B(n_2122),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2152),
.B(n_2155),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2155),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2153),
.B(n_2151),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_2150),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2162),
.B(n_2153),
.Y(n_2165)
);

NOR4xp25_ASAP7_75t_L g2166 ( 
.A(n_2161),
.B(n_2158),
.C(n_2159),
.D(n_2142),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2164),
.B(n_2157),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2163),
.Y(n_2168)
);

O2A1O1Ixp33_ASAP7_75t_SL g2169 ( 
.A1(n_2167),
.A2(n_2158),
.B(n_2159),
.C(n_2149),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2168),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2165),
.A2(n_2160),
.B1(n_2149),
.B2(n_2121),
.Y(n_2171)
);

OAI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2166),
.A2(n_2160),
.B1(n_2154),
.B2(n_2157),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2168),
.Y(n_2173)
);

INVxp33_ASAP7_75t_L g2174 ( 
.A(n_2167),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_SL g2175 ( 
.A1(n_2174),
.A2(n_2156),
.B(n_2154),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2169),
.Y(n_2176)
);

OAI21xp33_ASAP7_75t_L g2177 ( 
.A1(n_2170),
.A2(n_2118),
.B(n_2114),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2173),
.Y(n_2178)
);

AOI222xp33_ASAP7_75t_L g2179 ( 
.A1(n_2172),
.A2(n_2018),
.B1(n_2090),
.B2(n_2038),
.C1(n_2084),
.C2(n_2101),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2171),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2171),
.A2(n_2118),
.B1(n_2100),
.B2(n_2042),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2169),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2172),
.B(n_2119),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2171),
.A2(n_2046),
.B1(n_2071),
.B2(n_2090),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_L g2185 ( 
.A(n_2176),
.B(n_2004),
.C(n_1989),
.Y(n_2185)
);

AOI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_2183),
.A2(n_2071),
.B(n_2051),
.Y(n_2186)
);

AOI211xp5_ASAP7_75t_SL g2187 ( 
.A1(n_2182),
.A2(n_2057),
.B(n_1982),
.C(n_1959),
.Y(n_2187)
);

NAND3xp33_ASAP7_75t_SL g2188 ( 
.A(n_2181),
.B(n_2177),
.C(n_2175),
.Y(n_2188)
);

OAI22xp33_ASAP7_75t_SL g2189 ( 
.A1(n_2180),
.A2(n_2014),
.B1(n_2061),
.B2(n_2096),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2178),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2184),
.B(n_2014),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2179),
.B(n_2112),
.Y(n_2192)
);

INVx1_ASAP7_75t_SL g2193 ( 
.A(n_2176),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2178),
.Y(n_2194)
);

AOI21xp33_ASAP7_75t_SL g2195 ( 
.A1(n_2176),
.A2(n_227),
.B(n_228),
.Y(n_2195)
);

NAND3xp33_ASAP7_75t_SL g2196 ( 
.A(n_2176),
.B(n_2047),
.C(n_2075),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2178),
.Y(n_2197)
);

INVx1_ASAP7_75t_SL g2198 ( 
.A(n_2193),
.Y(n_2198)
);

NOR3xp33_ASAP7_75t_L g2199 ( 
.A(n_2188),
.B(n_1930),
.C(n_2060),
.Y(n_2199)
);

AOI221xp5_ASAP7_75t_L g2200 ( 
.A1(n_2195),
.A2(n_1982),
.B1(n_2080),
.B2(n_2075),
.C(n_1995),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2190),
.B(n_1942),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2194),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2197),
.B(n_1987),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2196),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2187),
.B(n_1995),
.C(n_1987),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2191),
.B(n_2096),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2189),
.B(n_2083),
.Y(n_2207)
);

INVx1_ASAP7_75t_SL g2208 ( 
.A(n_2192),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2185),
.B(n_2186),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2190),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2190),
.Y(n_2211)
);

BUFx2_ASAP7_75t_L g2212 ( 
.A(n_2190),
.Y(n_2212)
);

OAI322xp33_ASAP7_75t_L g2213 ( 
.A1(n_2198),
.A2(n_2075),
.A3(n_2087),
.B1(n_1995),
.B2(n_1987),
.C1(n_232),
.C2(n_233),
.Y(n_2213)
);

NOR2xp67_ASAP7_75t_L g2214 ( 
.A(n_2204),
.B(n_227),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2209),
.A2(n_2060),
.B(n_2027),
.Y(n_2215)
);

AO22x1_ASAP7_75t_L g2216 ( 
.A1(n_2212),
.A2(n_2002),
.B1(n_2052),
.B2(n_2022),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2199),
.A2(n_2080),
.B1(n_2022),
.B2(n_2056),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2210),
.B(n_228),
.Y(n_2218)
);

A2O1A1Ixp33_ASAP7_75t_L g2219 ( 
.A1(n_2201),
.A2(n_2027),
.B(n_2065),
.C(n_2035),
.Y(n_2219)
);

OAI211xp5_ASAP7_75t_SL g2220 ( 
.A1(n_2202),
.A2(n_232),
.B(n_229),
.C(n_230),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_2211),
.B(n_229),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2205),
.A2(n_2036),
.B1(n_2056),
.B2(n_2077),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2208),
.A2(n_2056),
.B1(n_2036),
.B2(n_2080),
.Y(n_2223)
);

NAND4xp25_ASAP7_75t_L g2224 ( 
.A(n_2203),
.B(n_2010),
.C(n_2077),
.D(n_2081),
.Y(n_2224)
);

AOI221xp5_ASAP7_75t_L g2225 ( 
.A1(n_2206),
.A2(n_2080),
.B1(n_2069),
.B2(n_1971),
.C(n_2087),
.Y(n_2225)
);

AOI211xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2207),
.A2(n_234),
.B(n_230),
.C(n_233),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_R g2227 ( 
.A(n_2221),
.B(n_234),
.Y(n_2227)
);

OAI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2214),
.A2(n_2200),
.B1(n_2077),
.B2(n_2086),
.C(n_2081),
.Y(n_2228)
);

AO22x2_ASAP7_75t_L g2229 ( 
.A1(n_2218),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2226),
.B(n_235),
.C(n_236),
.Y(n_2230)
);

NOR3xp33_ASAP7_75t_L g2231 ( 
.A(n_2220),
.B(n_237),
.C(n_238),
.Y(n_2231)
);

AOI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_2213),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_2232)
);

AOI321xp33_ASAP7_75t_L g2233 ( 
.A1(n_2217),
.A2(n_2010),
.A3(n_242),
.B1(n_244),
.B2(n_240),
.C(n_241),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_2222),
.B(n_1959),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2216),
.B(n_2054),
.Y(n_2235)
);

AOI221x1_ASAP7_75t_L g2236 ( 
.A1(n_2224),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_2236)
);

OAI211xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2225),
.A2(n_248),
.B(n_243),
.C(n_245),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2223),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2215),
.A2(n_248),
.B(n_249),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2219),
.B(n_2069),
.Y(n_2240)
);

OAI221xp5_ASAP7_75t_SL g2241 ( 
.A1(n_2217),
.A2(n_2086),
.B1(n_2081),
.B2(n_2054),
.C(n_2031),
.Y(n_2241)
);

NOR2x1_ASAP7_75t_L g2242 ( 
.A(n_2218),
.B(n_249),
.Y(n_2242)
);

AOI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2214),
.A2(n_2036),
.B1(n_2056),
.B2(n_2086),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_SL g2244 ( 
.A1(n_2226),
.A2(n_250),
.B(n_251),
.Y(n_2244)
);

AOI211xp5_ASAP7_75t_L g2245 ( 
.A1(n_2214),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_2245)
);

OAI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_2214),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2246)
);

OAI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2214),
.A2(n_2077),
.B1(n_2086),
.B2(n_2043),
.C(n_2036),
.Y(n_2247)
);

AOI221xp5_ASAP7_75t_L g2248 ( 
.A1(n_2213),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.C(n_256),
.Y(n_2248)
);

AOI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2228),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.C(n_260),
.Y(n_2249)
);

NAND3xp33_ASAP7_75t_SL g2250 ( 
.A(n_2244),
.B(n_257),
.C(n_258),
.Y(n_2250)
);

OAI21xp33_ASAP7_75t_L g2251 ( 
.A1(n_2231),
.A2(n_2053),
.B(n_2079),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2229),
.B(n_2242),
.Y(n_2252)
);

OAI211xp5_ASAP7_75t_L g2253 ( 
.A1(n_2232),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_2253)
);

OAI211xp5_ASAP7_75t_SL g2254 ( 
.A1(n_2238),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_2254)
);

AOI221xp5_ASAP7_75t_L g2255 ( 
.A1(n_2248),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2243),
.A2(n_2053),
.B1(n_2052),
.B2(n_2066),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_L g2257 ( 
.A1(n_2230),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2257)
);

A2O1A1Ixp33_ASAP7_75t_L g2258 ( 
.A1(n_2246),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_2258)
);

OAI21xp33_ASAP7_75t_SL g2259 ( 
.A1(n_2235),
.A2(n_2240),
.B(n_2234),
.Y(n_2259)
);

AOI211xp5_ASAP7_75t_L g2260 ( 
.A1(n_2237),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_2260)
);

A2O1A1Ixp33_ASAP7_75t_L g2261 ( 
.A1(n_2245),
.A2(n_272),
.B(n_269),
.C(n_271),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_2227),
.A2(n_2088),
.B1(n_2066),
.B2(n_2074),
.Y(n_2262)
);

OAI21xp33_ASAP7_75t_SL g2263 ( 
.A1(n_2247),
.A2(n_2035),
.B(n_2048),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2229),
.Y(n_2264)
);

NAND2x1p5_ASAP7_75t_L g2265 ( 
.A(n_2239),
.B(n_2052),
.Y(n_2265)
);

AOI221xp5_ASAP7_75t_L g2266 ( 
.A1(n_2241),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.C(n_276),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2236),
.B(n_273),
.Y(n_2267)
);

AOI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2233),
.A2(n_2088),
.B1(n_2066),
.B2(n_2074),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2244),
.B(n_274),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2239),
.A2(n_275),
.B(n_277),
.Y(n_2270)
);

AOI222xp33_ASAP7_75t_L g2271 ( 
.A1(n_2232),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.C1(n_280),
.C2(n_281),
.Y(n_2271)
);

AOI322xp5_ASAP7_75t_L g2272 ( 
.A1(n_2231),
.A2(n_2054),
.A3(n_2067),
.B1(n_2072),
.B2(n_2088),
.C1(n_1943),
.C2(n_2111),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2229),
.Y(n_2273)
);

AOI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2228),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.C(n_282),
.Y(n_2274)
);

AOI221xp5_ASAP7_75t_L g2275 ( 
.A1(n_2228),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2275)
);

AOI222xp33_ASAP7_75t_L g2276 ( 
.A1(n_2232),
.A2(n_283),
.B1(n_284),
.B2(n_286),
.C1(n_287),
.C2(n_288),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2243),
.A2(n_2052),
.B1(n_2072),
.B2(n_2067),
.Y(n_2277)
);

AOI211xp5_ASAP7_75t_L g2278 ( 
.A1(n_2244),
.A2(n_290),
.B(n_286),
.C(n_289),
.Y(n_2278)
);

OAI321xp33_ASAP7_75t_L g2279 ( 
.A1(n_2237),
.A2(n_2082),
.A3(n_291),
.B1(n_292),
.B2(n_293),
.C(n_294),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_SL g2280 ( 
.A1(n_2228),
.A2(n_2111),
.B1(n_2108),
.B2(n_2098),
.Y(n_2280)
);

NOR4xp25_ASAP7_75t_L g2281 ( 
.A(n_2244),
.B(n_292),
.C(n_289),
.D(n_291),
.Y(n_2281)
);

OAI21xp5_ASAP7_75t_SL g2282 ( 
.A1(n_2244),
.A2(n_293),
.B(n_295),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2242),
.Y(n_2283)
);

AOI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2228),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2242),
.Y(n_2285)
);

AOI21xp33_ASAP7_75t_L g2286 ( 
.A1(n_2283),
.A2(n_296),
.B(n_298),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2267),
.A2(n_2088),
.B1(n_2074),
.B2(n_2095),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2264),
.B(n_299),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2252),
.Y(n_2289)
);

NAND3xp33_ASAP7_75t_L g2290 ( 
.A(n_2278),
.B(n_299),
.C(n_300),
.Y(n_2290)
);

NAND3xp33_ASAP7_75t_SL g2291 ( 
.A(n_2281),
.B(n_301),
.C(n_302),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2273),
.B(n_301),
.Y(n_2292)
);

NOR3x2_ASAP7_75t_L g2293 ( 
.A(n_2285),
.B(n_302),
.C(n_303),
.Y(n_2293)
);

NAND4xp25_ASAP7_75t_L g2294 ( 
.A(n_2260),
.B(n_305),
.C(n_303),
.D(n_304),
.Y(n_2294)
);

NOR2x1_ASAP7_75t_L g2295 ( 
.A(n_2250),
.B(n_304),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2258),
.B(n_305),
.Y(n_2296)
);

INVxp67_ASAP7_75t_L g2297 ( 
.A(n_2269),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2254),
.B(n_2282),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2270),
.A2(n_2065),
.B(n_2048),
.Y(n_2299)
);

NOR2x1_ASAP7_75t_L g2300 ( 
.A(n_2261),
.B(n_306),
.Y(n_2300)
);

NOR2x1_ASAP7_75t_L g2301 ( 
.A(n_2253),
.B(n_307),
.Y(n_2301)
);

NOR3xp33_ASAP7_75t_L g2302 ( 
.A(n_2255),
.B(n_2274),
.C(n_2249),
.Y(n_2302)
);

OAI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_2251),
.A2(n_2079),
.B(n_2088),
.Y(n_2303)
);

NOR3x2_ASAP7_75t_L g2304 ( 
.A(n_2257),
.B(n_307),
.C(n_308),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2265),
.Y(n_2305)
);

NAND3xp33_ASAP7_75t_L g2306 ( 
.A(n_2271),
.B(n_308),
.C(n_309),
.Y(n_2306)
);

OAI22x1_ASAP7_75t_L g2307 ( 
.A1(n_2265),
.A2(n_2049),
.B1(n_2082),
.B2(n_311),
.Y(n_2307)
);

NOR2x1_ASAP7_75t_L g2308 ( 
.A(n_2256),
.B(n_309),
.Y(n_2308)
);

NAND3xp33_ASAP7_75t_L g2309 ( 
.A(n_2276),
.B(n_310),
.C(n_311),
.Y(n_2309)
);

NOR2xp67_ASAP7_75t_L g2310 ( 
.A(n_2279),
.B(n_312),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_L g2311 ( 
.A(n_2277),
.B(n_312),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2262),
.B(n_2054),
.Y(n_2312)
);

NAND3xp33_ASAP7_75t_SL g2313 ( 
.A(n_2275),
.B(n_2284),
.C(n_2266),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2259),
.Y(n_2314)
);

OAI211xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2263),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_2315)
);

NOR2xp67_ASAP7_75t_L g2316 ( 
.A(n_2268),
.B(n_313),
.Y(n_2316)
);

NOR3xp33_ASAP7_75t_L g2317 ( 
.A(n_2280),
.B(n_314),
.C(n_315),
.Y(n_2317)
);

HB1xp67_ASAP7_75t_L g2318 ( 
.A(n_2272),
.Y(n_2318)
);

NAND4xp25_ASAP7_75t_L g2319 ( 
.A(n_2260),
.B(n_318),
.C(n_316),
.D(n_317),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2252),
.B(n_2074),
.Y(n_2320)
);

NAND3xp33_ASAP7_75t_SL g2321 ( 
.A(n_2278),
.B(n_316),
.C(n_317),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2252),
.B(n_319),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2252),
.Y(n_2323)
);

NAND4xp75_ASAP7_75t_L g2324 ( 
.A(n_2288),
.B(n_322),
.C(n_320),
.D(n_321),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2322),
.B(n_320),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2294),
.B(n_321),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2293),
.Y(n_2327)
);

AND3x4_ASAP7_75t_L g2328 ( 
.A(n_2310),
.B(n_323),
.C(n_324),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2291),
.B(n_323),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2320),
.B(n_2099),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2292),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2289),
.B(n_324),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2323),
.B(n_2099),
.Y(n_2333)
);

NOR2x1_ASAP7_75t_L g2334 ( 
.A(n_2305),
.B(n_325),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2298),
.B(n_2079),
.Y(n_2335)
);

NOR2x1_ASAP7_75t_L g2336 ( 
.A(n_2295),
.B(n_2321),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2300),
.B(n_325),
.Y(n_2337)
);

NOR2x1_ASAP7_75t_L g2338 ( 
.A(n_2314),
.B(n_2290),
.Y(n_2338)
);

A2O1A1Ixp33_ASAP7_75t_L g2339 ( 
.A1(n_2316),
.A2(n_329),
.B(n_326),
.C(n_327),
.Y(n_2339)
);

NAND2x1_ASAP7_75t_SL g2340 ( 
.A(n_2301),
.B(n_327),
.Y(n_2340)
);

NAND2x1p5_ASAP7_75t_SL g2341 ( 
.A(n_2308),
.B(n_330),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2296),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2317),
.B(n_330),
.Y(n_2343)
);

NAND4xp75_ASAP7_75t_L g2344 ( 
.A(n_2311),
.B(n_333),
.C(n_331),
.D(n_332),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2287),
.B(n_331),
.Y(n_2345)
);

NOR2x1_ASAP7_75t_L g2346 ( 
.A(n_2319),
.B(n_332),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_2306),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2313),
.A2(n_333),
.B(n_334),
.Y(n_2348)
);

NOR3x2_ASAP7_75t_L g2349 ( 
.A(n_2304),
.B(n_334),
.C(n_335),
.Y(n_2349)
);

NOR2x1_ASAP7_75t_L g2350 ( 
.A(n_2309),
.B(n_335),
.Y(n_2350)
);

NAND3xp33_ASAP7_75t_SL g2351 ( 
.A(n_2302),
.B(n_336),
.C(n_337),
.Y(n_2351)
);

AND3x4_ASAP7_75t_L g2352 ( 
.A(n_2297),
.B(n_337),
.C(n_338),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2286),
.B(n_339),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2318),
.B(n_339),
.Y(n_2354)
);

OA21x2_ASAP7_75t_L g2355 ( 
.A1(n_2303),
.A2(n_340),
.B(n_341),
.Y(n_2355)
);

OAI21xp33_ASAP7_75t_SL g2356 ( 
.A1(n_2312),
.A2(n_2065),
.B(n_341),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2307),
.B(n_342),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2315),
.A2(n_342),
.B(n_343),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2299),
.Y(n_2359)
);

NOR3xp33_ASAP7_75t_L g2360 ( 
.A(n_2289),
.B(n_344),
.C(n_345),
.Y(n_2360)
);

AOI211x1_ASAP7_75t_L g2361 ( 
.A1(n_2291),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2320),
.B(n_2095),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2293),
.Y(n_2363)
);

NOR2x1p5_ASAP7_75t_L g2364 ( 
.A(n_2291),
.B(n_347),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2289),
.B(n_348),
.C(n_349),
.Y(n_2365)
);

NAND4xp75_ASAP7_75t_L g2366 ( 
.A(n_2288),
.B(n_350),
.C(n_348),
.D(n_349),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2320),
.B(n_351),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2288),
.B(n_351),
.Y(n_2368)
);

AO22x2_ASAP7_75t_L g2369 ( 
.A1(n_2289),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_2289),
.Y(n_2370)
);

NOR3xp33_ASAP7_75t_SL g2371 ( 
.A(n_2291),
.B(n_354),
.C(n_356),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_2289),
.B(n_356),
.C(n_358),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2320),
.B(n_358),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2320),
.B(n_359),
.Y(n_2374)
);

NAND2x1p5_ASAP7_75t_L g2375 ( 
.A(n_2288),
.B(n_360),
.Y(n_2375)
);

OR2x2_ASAP7_75t_L g2376 ( 
.A(n_2322),
.B(n_360),
.Y(n_2376)
);

NOR2x1p5_ASAP7_75t_L g2377 ( 
.A(n_2291),
.B(n_361),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2320),
.B(n_2098),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2293),
.Y(n_2379)
);

NOR2x1_ASAP7_75t_L g2380 ( 
.A(n_2288),
.B(n_361),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2320),
.B(n_362),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2289),
.A2(n_2106),
.B1(n_2069),
.B2(n_2049),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2322),
.B(n_362),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2288),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2294),
.B(n_363),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2380),
.B(n_363),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2368),
.B(n_364),
.Y(n_2387)
);

NAND3xp33_ASAP7_75t_L g2388 ( 
.A(n_2360),
.B(n_364),
.C(n_365),
.Y(n_2388)
);

NOR3xp33_ASAP7_75t_L g2389 ( 
.A(n_2354),
.B(n_366),
.C(n_367),
.Y(n_2389)
);

XNOR2xp5_ASAP7_75t_L g2390 ( 
.A(n_2328),
.B(n_367),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2369),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2369),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2367),
.B(n_368),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2368),
.Y(n_2394)
);

OAI322xp33_ASAP7_75t_L g2395 ( 
.A1(n_2327),
.A2(n_369),
.A3(n_370),
.B1(n_371),
.B2(n_372),
.C1(n_373),
.C2(n_374),
.Y(n_2395)
);

OR5x1_ASAP7_75t_L g2396 ( 
.A(n_2351),
.B(n_371),
.C(n_372),
.D(n_373),
.E(n_374),
.Y(n_2396)
);

NAND3x1_ASAP7_75t_L g2397 ( 
.A(n_2334),
.B(n_375),
.C(n_376),
.Y(n_2397)
);

AO22x2_ASAP7_75t_L g2398 ( 
.A1(n_2363),
.A2(n_2379),
.B1(n_2344),
.B2(n_2347),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2365),
.B(n_378),
.Y(n_2399)
);

NAND4xp75_ASAP7_75t_L g2400 ( 
.A(n_2338),
.B(n_2336),
.C(n_2350),
.D(n_2329),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2370),
.A2(n_2106),
.B1(n_2069),
.B2(n_2049),
.Y(n_2401)
);

BUFx2_ASAP7_75t_L g2402 ( 
.A(n_2340),
.Y(n_2402)
);

AOI211xp5_ASAP7_75t_L g2403 ( 
.A1(n_2348),
.A2(n_378),
.B(n_379),
.C(n_380),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2375),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2337),
.B(n_379),
.Y(n_2405)
);

XOR2x2_ASAP7_75t_L g2406 ( 
.A(n_2324),
.B(n_2366),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2373),
.B(n_380),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2352),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2374),
.A2(n_2031),
.B1(n_2091),
.B2(n_2083),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2341),
.B(n_2381),
.Y(n_2410)
);

NAND2x1p5_ASAP7_75t_L g2411 ( 
.A(n_2337),
.B(n_381),
.Y(n_2411)
);

NAND5xp2_ASAP7_75t_L g2412 ( 
.A(n_2371),
.B(n_381),
.C(n_382),
.D(n_383),
.E(n_384),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2335),
.B(n_382),
.Y(n_2413)
);

NAND4xp25_ASAP7_75t_L g2414 ( 
.A(n_2361),
.B(n_383),
.C(n_384),
.D(n_385),
.Y(n_2414)
);

AND3x4_ASAP7_75t_L g2415 ( 
.A(n_2346),
.B(n_386),
.C(n_387),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2372),
.B(n_386),
.C(n_387),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2384),
.Y(n_2417)
);

BUFx12f_ASAP7_75t_L g2418 ( 
.A(n_2364),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2332),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2325),
.Y(n_2420)
);

NAND2x1p5_ASAP7_75t_L g2421 ( 
.A(n_2377),
.B(n_389),
.Y(n_2421)
);

NOR3xp33_ASAP7_75t_L g2422 ( 
.A(n_2353),
.B(n_389),
.C(n_390),
.Y(n_2422)
);

OAI21xp5_ASAP7_75t_SL g2423 ( 
.A1(n_2385),
.A2(n_390),
.B(n_391),
.Y(n_2423)
);

NAND2x1p5_ASAP7_75t_L g2424 ( 
.A(n_2376),
.B(n_391),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2339),
.B(n_392),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2358),
.B(n_392),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2355),
.B(n_2357),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2383),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2355),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2326),
.B(n_393),
.Y(n_2430)
);

NOR3xp33_ASAP7_75t_L g2431 ( 
.A(n_2343),
.B(n_394),
.C(n_395),
.Y(n_2431)
);

NOR3xp33_ASAP7_75t_SL g2432 ( 
.A(n_2345),
.B(n_394),
.C(n_395),
.Y(n_2432)
);

OR2x2_ASAP7_75t_L g2433 ( 
.A(n_2331),
.B(n_397),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2349),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_SL g2435 ( 
.A1(n_2342),
.A2(n_397),
.B(n_398),
.Y(n_2435)
);

NOR3xp33_ASAP7_75t_L g2436 ( 
.A(n_2359),
.B(n_398),
.C(n_399),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2333),
.B(n_399),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2330),
.B(n_400),
.Y(n_2438)
);

NOR3xp33_ASAP7_75t_L g2439 ( 
.A(n_2356),
.B(n_400),
.C(n_401),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2362),
.B(n_401),
.Y(n_2440)
);

NAND5xp2_ASAP7_75t_L g2441 ( 
.A(n_2378),
.B(n_402),
.C(n_403),
.D(n_404),
.E(n_405),
.Y(n_2441)
);

OAI211xp5_ASAP7_75t_L g2442 ( 
.A1(n_2382),
.A2(n_403),
.B(n_404),
.C(n_405),
.Y(n_2442)
);

AND2x4_ASAP7_75t_L g2443 ( 
.A(n_2380),
.B(n_406),
.Y(n_2443)
);

NAND4xp75_ASAP7_75t_L g2444 ( 
.A(n_2334),
.B(n_406),
.C(n_407),
.D(n_408),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2368),
.B(n_407),
.Y(n_2445)
);

AND4x1_ASAP7_75t_L g2446 ( 
.A(n_2338),
.B(n_408),
.C(n_409),
.D(n_410),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2368),
.Y(n_2447)
);

AOI211xp5_ASAP7_75t_L g2448 ( 
.A1(n_2351),
.A2(n_409),
.B(n_410),
.C(n_411),
.Y(n_2448)
);

CKINVDCx20_ASAP7_75t_R g2449 ( 
.A(n_2370),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2368),
.B(n_411),
.Y(n_2450)
);

NOR2xp67_ASAP7_75t_L g2451 ( 
.A(n_2384),
.B(n_413),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2368),
.B(n_413),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_R g2453 ( 
.A(n_2449),
.B(n_414),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_R g2454 ( 
.A(n_2390),
.B(n_415),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_2405),
.B(n_416),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2451),
.B(n_416),
.Y(n_2456)
);

NAND3xp33_ASAP7_75t_SL g2457 ( 
.A(n_2415),
.B(n_417),
.C(n_418),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2405),
.B(n_417),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2413),
.B(n_419),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_R g2460 ( 
.A(n_2429),
.B(n_419),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_R g2461 ( 
.A(n_2402),
.B(n_420),
.Y(n_2461)
);

NAND2xp33_ASAP7_75t_SL g2462 ( 
.A(n_2432),
.B(n_420),
.Y(n_2462)
);

NAND2xp33_ASAP7_75t_SL g2463 ( 
.A(n_2387),
.B(n_421),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2386),
.B(n_422),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2404),
.B(n_422),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2386),
.B(n_423),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_R g2467 ( 
.A(n_2394),
.B(n_423),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2443),
.B(n_424),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_R g2469 ( 
.A(n_2447),
.B(n_424),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2443),
.B(n_425),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_R g2471 ( 
.A(n_2418),
.B(n_425),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2446),
.B(n_427),
.Y(n_2472)
);

XNOR2xp5_ASAP7_75t_L g2473 ( 
.A(n_2406),
.B(n_427),
.Y(n_2473)
);

XNOR2xp5_ASAP7_75t_L g2474 ( 
.A(n_2397),
.B(n_2396),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_SL g2475 ( 
.A(n_2411),
.B(n_428),
.C(n_429),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2448),
.B(n_428),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2403),
.B(n_2417),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2391),
.B(n_429),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_SL g2479 ( 
.A(n_2445),
.B(n_430),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_R g2480 ( 
.A(n_2434),
.B(n_430),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2393),
.B(n_431),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2407),
.B(n_431),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_SL g2483 ( 
.A(n_2444),
.B(n_432),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_R g2484 ( 
.A(n_2408),
.B(n_432),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_2392),
.B(n_433),
.Y(n_2485)
);

NAND3xp33_ASAP7_75t_L g2486 ( 
.A(n_2422),
.B(n_433),
.C(n_434),
.Y(n_2486)
);

NAND3xp33_ASAP7_75t_L g2487 ( 
.A(n_2431),
.B(n_2389),
.C(n_2436),
.Y(n_2487)
);

NAND2xp33_ASAP7_75t_SL g2488 ( 
.A(n_2450),
.B(n_2452),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2439),
.B(n_436),
.Y(n_2489)
);

NAND2x1_ASAP7_75t_SL g2490 ( 
.A(n_2430),
.B(n_436),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2424),
.B(n_437),
.Y(n_2491)
);

XNOR2xp5_ASAP7_75t_L g2492 ( 
.A(n_2398),
.B(n_437),
.Y(n_2492)
);

XNOR2xp5_ASAP7_75t_L g2493 ( 
.A(n_2398),
.B(n_438),
.Y(n_2493)
);

NAND2xp33_ASAP7_75t_SL g2494 ( 
.A(n_2438),
.B(n_2410),
.Y(n_2494)
);

NAND2xp33_ASAP7_75t_SL g2495 ( 
.A(n_2427),
.B(n_438),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_R g2496 ( 
.A(n_2426),
.B(n_439),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_R g2497 ( 
.A(n_2399),
.B(n_2420),
.Y(n_2497)
);

NAND3xp33_ASAP7_75t_L g2498 ( 
.A(n_2423),
.B(n_439),
.C(n_440),
.Y(n_2498)
);

NOR3xp33_ASAP7_75t_SL g2499 ( 
.A(n_2400),
.B(n_2412),
.C(n_2414),
.Y(n_2499)
);

NAND2xp33_ASAP7_75t_SL g2500 ( 
.A(n_2425),
.B(n_440),
.Y(n_2500)
);

NAND3xp33_ASAP7_75t_SL g2501 ( 
.A(n_2421),
.B(n_441),
.C(n_442),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2435),
.B(n_441),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_R g2503 ( 
.A(n_2428),
.B(n_442),
.Y(n_2503)
);

NAND2xp33_ASAP7_75t_SL g2504 ( 
.A(n_2437),
.B(n_443),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2388),
.B(n_444),
.Y(n_2505)
);

NAND2xp33_ASAP7_75t_SL g2506 ( 
.A(n_2440),
.B(n_444),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2416),
.B(n_445),
.Y(n_2507)
);

XNOR2xp5_ASAP7_75t_L g2508 ( 
.A(n_2419),
.B(n_445),
.Y(n_2508)
);

OAI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2492),
.A2(n_2442),
.B1(n_2433),
.B2(n_2409),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2493),
.A2(n_2401),
.B1(n_2441),
.B2(n_2395),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2473),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2490),
.Y(n_2512)
);

INVxp67_ASAP7_75t_L g2513 ( 
.A(n_2483),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2508),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2471),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2464),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2466),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2470),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2456),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2502),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2459),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2455),
.Y(n_2522)
);

OAI211xp5_ASAP7_75t_L g2523 ( 
.A1(n_2460),
.A2(n_446),
.B(n_447),
.C(n_448),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2458),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2491),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2478),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2485),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2474),
.Y(n_2528)
);

AO22x1_ASAP7_75t_L g2529 ( 
.A1(n_2481),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_2529)
);

BUFx3_ASAP7_75t_L g2530 ( 
.A(n_2482),
.Y(n_2530)
);

BUFx2_ASAP7_75t_L g2531 ( 
.A(n_2467),
.Y(n_2531)
);

INVxp67_ASAP7_75t_L g2532 ( 
.A(n_2468),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2499),
.B(n_1943),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2489),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2472),
.Y(n_2535)
);

AO22x1_ASAP7_75t_L g2536 ( 
.A1(n_2495),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_2536)
);

OAI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2498),
.A2(n_2091),
.B1(n_2069),
.B2(n_2043),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2475),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2469),
.Y(n_2539)
);

AND2x4_ASAP7_75t_L g2540 ( 
.A(n_2486),
.B(n_449),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2461),
.Y(n_2541)
);

OAI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2487),
.A2(n_2476),
.B1(n_2477),
.B2(n_2505),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2501),
.Y(n_2543)
);

OA22x2_ASAP7_75t_L g2544 ( 
.A1(n_2507),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2453),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2465),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2494),
.A2(n_452),
.B1(n_453),
.B2(n_455),
.Y(n_2547)
);

OA22x2_ASAP7_75t_L g2548 ( 
.A1(n_2463),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2480),
.A2(n_2454),
.B1(n_2462),
.B2(n_2457),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2484),
.Y(n_2550)
);

XNOR2xp5_ASAP7_75t_L g2551 ( 
.A(n_2528),
.B(n_2504),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2548),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2544),
.Y(n_2553)
);

OAI22x1_ASAP7_75t_L g2554 ( 
.A1(n_2512),
.A2(n_2496),
.B1(n_2479),
.B2(n_2506),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2536),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_SL g2556 ( 
.A1(n_2540),
.A2(n_2500),
.B1(n_2503),
.B2(n_2488),
.Y(n_2556)
);

OAI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2513),
.A2(n_2497),
.B1(n_2503),
.B2(n_459),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_SL g2558 ( 
.A1(n_2533),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2529),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2515),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_2560)
);

INVx4_ASAP7_75t_L g2561 ( 
.A(n_2531),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2529),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2538),
.B(n_460),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2539),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2523),
.Y(n_2565)
);

OAI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2532),
.A2(n_2543),
.B1(n_2511),
.B2(n_2535),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_SL g2567 ( 
.A1(n_2541),
.A2(n_461),
.B1(n_462),
.B2(n_463),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2540),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2510),
.Y(n_2569)
);

XOR2xp5_ASAP7_75t_L g2570 ( 
.A(n_2549),
.B(n_463),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2546),
.Y(n_2571)
);

NAND4xp25_ASAP7_75t_L g2572 ( 
.A(n_2542),
.B(n_464),
.C(n_465),
.D(n_466),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2522),
.Y(n_2573)
);

OAI22x1_ASAP7_75t_L g2574 ( 
.A1(n_2547),
.A2(n_464),
.B1(n_465),
.B2(n_466),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2524),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2526),
.B(n_467),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2550),
.Y(n_2577)
);

OAI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2527),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2545),
.Y(n_2579)
);

OR3x2_ASAP7_75t_L g2580 ( 
.A(n_2573),
.B(n_2520),
.C(n_2518),
.Y(n_2580)
);

OAI22x1_ASAP7_75t_L g2581 ( 
.A1(n_2570),
.A2(n_2514),
.B1(n_2517),
.B2(n_2525),
.Y(n_2581)
);

OAI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2551),
.A2(n_2509),
.B(n_2516),
.Y(n_2582)
);

AOI22xp33_ASAP7_75t_L g2583 ( 
.A1(n_2561),
.A2(n_2530),
.B1(n_2521),
.B2(n_2519),
.Y(n_2583)
);

BUFx2_ASAP7_75t_L g2584 ( 
.A(n_2562),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2557),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2555),
.Y(n_2586)
);

CKINVDCx20_ASAP7_75t_R g2587 ( 
.A(n_2569),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2574),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2559),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2552),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2579),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2576),
.Y(n_2592)
);

NAND3xp33_ASAP7_75t_L g2593 ( 
.A(n_2558),
.B(n_2534),
.C(n_2537),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2556),
.B(n_470),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2553),
.B(n_471),
.Y(n_2595)
);

OA21x2_ASAP7_75t_L g2596 ( 
.A1(n_2575),
.A2(n_472),
.B(n_473),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2563),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2572),
.B(n_472),
.Y(n_2598)
);

INVx2_ASAP7_75t_SL g2599 ( 
.A(n_2592),
.Y(n_2599)
);

CKINVDCx20_ASAP7_75t_R g2600 ( 
.A(n_2587),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2584),
.A2(n_2564),
.B1(n_2577),
.B2(n_2571),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2591),
.A2(n_2590),
.B1(n_2586),
.B2(n_2566),
.Y(n_2602)
);

OAI22xp5_ASAP7_75t_L g2603 ( 
.A1(n_2583),
.A2(n_2565),
.B1(n_2568),
.B2(n_2560),
.Y(n_2603)
);

OAI22x1_ASAP7_75t_L g2604 ( 
.A1(n_2588),
.A2(n_2589),
.B1(n_2595),
.B2(n_2594),
.Y(n_2604)
);

OA22x2_ASAP7_75t_L g2605 ( 
.A1(n_2582),
.A2(n_2554),
.B1(n_2567),
.B2(n_2578),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2598),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2580),
.A2(n_2576),
.B1(n_475),
.B2(n_476),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2581),
.A2(n_2593),
.B(n_2585),
.Y(n_2608)
);

INVx3_ASAP7_75t_SL g2609 ( 
.A(n_2597),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2596),
.A2(n_473),
.B1(n_476),
.B2(n_477),
.Y(n_2610)
);

AOI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2600),
.A2(n_2596),
.B1(n_478),
.B2(n_479),
.Y(n_2611)
);

OA22x2_ASAP7_75t_L g2612 ( 
.A1(n_2607),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_2612)
);

AOI21xp33_ASAP7_75t_L g2613 ( 
.A1(n_2599),
.A2(n_480),
.B(n_481),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2602),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_L g2615 ( 
.A(n_2601),
.B(n_2608),
.C(n_2603),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2605),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_2616)
);

OAI22x1_ASAP7_75t_L g2617 ( 
.A1(n_2609),
.A2(n_2606),
.B1(n_2604),
.B2(n_2610),
.Y(n_2617)
);

OAI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2608),
.A2(n_482),
.B(n_483),
.Y(n_2618)
);

OAI21xp5_ASAP7_75t_L g2619 ( 
.A1(n_2615),
.A2(n_483),
.B(n_484),
.Y(n_2619)
);

CKINVDCx20_ASAP7_75t_R g2620 ( 
.A(n_2614),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2618),
.B(n_486),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2612),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2611),
.B(n_2616),
.Y(n_2623)
);

INVxp33_ASAP7_75t_L g2624 ( 
.A(n_2617),
.Y(n_2624)
);

NAND5xp2_ASAP7_75t_L g2625 ( 
.A(n_2624),
.B(n_2613),
.C(n_487),
.D(n_488),
.E(n_489),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2620),
.A2(n_486),
.B1(n_487),
.B2(n_490),
.Y(n_2626)
);

XNOR2xp5_ASAP7_75t_L g2627 ( 
.A(n_2621),
.B(n_491),
.Y(n_2627)
);

OAI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2619),
.A2(n_2622),
.B1(n_2623),
.B2(n_495),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2627),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_SL g2630 ( 
.A1(n_2628),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2630)
);

NAND3xp33_ASAP7_75t_L g2631 ( 
.A(n_2629),
.B(n_2626),
.C(n_2625),
.Y(n_2631)
);

OAI31xp33_ASAP7_75t_L g2632 ( 
.A1(n_2631),
.A2(n_2630),
.A3(n_497),
.B(n_499),
.Y(n_2632)
);

AOI221xp5_ASAP7_75t_L g2633 ( 
.A1(n_2632),
.A2(n_496),
.B1(n_499),
.B2(n_500),
.C(n_501),
.Y(n_2633)
);

AOI221xp5_ASAP7_75t_L g2634 ( 
.A1(n_2633),
.A2(n_501),
.B1(n_502),
.B2(n_504),
.C(n_505),
.Y(n_2634)
);

AOI211xp5_ASAP7_75t_L g2635 ( 
.A1(n_2634),
.A2(n_504),
.B(n_505),
.C(n_506),
.Y(n_2635)
);


endmodule