module fake_netlist_5_2483_n_572 (n_10, n_24, n_61, n_75, n_65, n_78, n_74, n_57, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_38, n_80, n_4, n_35, n_73, n_17, n_19, n_30, n_5, n_33, n_14, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_27, n_64, n_77, n_81, n_28, n_70, n_68, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_572);

input n_10;
input n_24;
input n_61;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_70;
input n_68;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;

output n_572;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_82;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_124;
wire n_146;
wire n_86;
wire n_136;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_111;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_116;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_551;
wire n_382;
wire n_554;
wire n_254;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_100;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_119;
wire n_497;
wire n_559;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_87;
wire n_150;
wire n_530;
wire n_556;
wire n_106;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_93;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_90;
wire n_546;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_94;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_95;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_104;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_145;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_88;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_98;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_107;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_92;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_84;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_112;
wire n_542;
wire n_85;
wire n_463;
wire n_488;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_102;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_91;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_83;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_487;
wire n_495;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_99;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_89;
wire n_438;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;
wire n_110;

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVxp33_ASAP7_75t_SL g92 ( 
.A(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_7),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_76),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_61),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_10),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_46),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_5),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_2),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

BUFx8_ASAP7_75t_SL g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_11),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_15),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_32),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_24),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_36),
.Y(n_143)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_1),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_30),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_50),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_19),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_9),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_27),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_15),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_35),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_47),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_85),
.B(n_3),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_4),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_6),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_91),
.B(n_6),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_91),
.B(n_9),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_R g188 ( 
.A(n_108),
.B(n_13),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_R g190 ( 
.A(n_108),
.B(n_13),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

NAND2x1p5_ASAP7_75t_L g194 ( 
.A(n_99),
.B(n_39),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_14),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_14),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_153),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_98),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_101),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_144),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_102),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_137),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_99),
.B(n_110),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_99),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_124),
.B(n_18),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_R g229 ( 
.A(n_117),
.B(n_23),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_86),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_173),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

AO22x2_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_110),
.B1(n_93),
.B2(n_82),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

AO22x2_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_93),
.B1(n_120),
.B2(n_96),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_138),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_165),
.Y(n_248)
);

AO22x2_ASAP7_75t_L g249 ( 
.A1(n_163),
.A2(n_122),
.B1(n_156),
.B2(n_151),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_138),
.B1(n_124),
.B2(n_149),
.Y(n_250)
);

NAND3x1_ASAP7_75t_L g251 ( 
.A(n_169),
.B(n_118),
.C(n_150),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_186),
.A2(n_112),
.B1(n_88),
.B2(n_84),
.C(n_157),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_167),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_166),
.B(n_147),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

OR2x2_ASAP7_75t_SL g258 ( 
.A(n_206),
.B(n_143),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_140),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_182),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_160),
.B(n_136),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_163),
.B(n_106),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_206),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_94),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_199),
.B(n_107),
.Y(n_275)
);

NAND2x1p5_ASAP7_75t_L g276 ( 
.A(n_198),
.B(n_134),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_135),
.Y(n_278)
);

NAND3x1_ASAP7_75t_L g279 ( 
.A(n_169),
.B(n_162),
.C(n_128),
.Y(n_279)
);

OAI221xp5_ASAP7_75t_L g280 ( 
.A1(n_173),
.A2(n_126),
.B1(n_121),
.B2(n_119),
.C(n_42),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_199),
.B(n_28),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_195),
.B(n_31),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_41),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_174),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_53),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_222),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_194),
.B1(n_222),
.B2(n_197),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_222),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_254),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_244),
.B(n_194),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_217),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g299 ( 
.A(n_252),
.B(n_215),
.C(n_214),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_189),
.B1(n_197),
.B2(n_212),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_185),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_244),
.B(n_208),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_272),
.A2(n_205),
.B(n_217),
.Y(n_304)
);

AND3x2_ASAP7_75t_SL g305 ( 
.A(n_239),
.B(n_219),
.C(n_216),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_216),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_205),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_185),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_248),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_201),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_201),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_SL g323 ( 
.A(n_264),
.B(n_161),
.C(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_259),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_267),
.B(n_229),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_264),
.B(n_255),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_229),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_196),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_255),
.B(n_190),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_262),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_239),
.A2(n_183),
.B1(n_192),
.B2(n_191),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_247),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_233),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_248),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_231),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_276),
.B(n_184),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_237),
.B(n_164),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_271),
.B(n_172),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_340),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_279),
.B1(n_237),
.B2(n_258),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_234),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

BUFx4f_ASAP7_75t_SL g354 ( 
.A(n_312),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_237),
.B(n_278),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_307),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_261),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_295),
.A2(n_250),
.B1(n_280),
.B2(n_235),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_311),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_316),
.A2(n_175),
.B1(n_176),
.B2(n_288),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_291),
.B(n_288),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_249),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_249),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_280),
.B1(n_251),
.B2(n_249),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_234),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_314),
.B(n_273),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_303),
.B(n_277),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_240),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_236),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_243),
.Y(n_386)
);

O2A1O1Ixp5_ASAP7_75t_SL g387 ( 
.A1(n_315),
.A2(n_230),
.B(n_232),
.C(n_179),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_193),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_290),
.A2(n_278),
.B(n_285),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_297),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_318),
.B(n_263),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_270),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_292),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

O2A1O1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_327),
.A2(n_282),
.B(n_188),
.C(n_190),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_313),
.A2(n_287),
.B(n_274),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_188),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_322),
.B(n_274),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_274),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_335),
.A2(n_274),
.B1(n_287),
.B2(n_73),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_304),
.A2(n_287),
.B(n_79),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_309),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_365),
.A2(n_291),
.B1(n_335),
.B2(n_322),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

AOI221xp5_ASAP7_75t_SL g416 ( 
.A1(n_350),
.A2(n_301),
.B1(n_342),
.B2(n_305),
.C(n_326),
.Y(n_416)
);

AOI221xp5_ASAP7_75t_L g417 ( 
.A1(n_360),
.A2(n_301),
.B1(n_299),
.B2(n_305),
.C(n_323),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_339),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_363),
.B(n_294),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_400),
.B(n_294),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_296),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_397),
.A2(n_296),
.B(n_300),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_365),
.A2(n_383),
.B1(n_366),
.B2(n_371),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_300),
.B1(n_317),
.B2(n_333),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_357),
.B(n_389),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_362),
.B(n_317),
.Y(n_428)
);

CKINVDCx10_ASAP7_75t_R g429 ( 
.A(n_354),
.Y(n_429)
);

OR2x6_ASAP7_75t_SL g430 ( 
.A(n_368),
.B(n_330),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_383),
.A2(n_333),
.B1(n_321),
.B2(n_330),
.Y(n_431)
);

AO21x2_ASAP7_75t_L g432 ( 
.A1(n_357),
.A2(n_344),
.B(n_321),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_348),
.B(n_321),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_355),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_383),
.A2(n_321),
.B1(n_344),
.B2(n_287),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_347),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_359),
.A2(n_364),
.B1(n_381),
.B2(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_404),
.A2(n_394),
.B1(n_348),
.B2(n_359),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_384),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_408),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_393),
.A2(n_385),
.B(n_402),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_377),
.B(n_408),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_349),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_SL g449 ( 
.A(n_379),
.B(n_404),
.C(n_396),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_356),
.B(n_386),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_348),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_R g455 ( 
.A(n_370),
.B(n_378),
.Y(n_455)
);

AOI221xp5_ASAP7_75t_L g456 ( 
.A1(n_375),
.A2(n_390),
.B1(n_398),
.B2(n_378),
.C(n_396),
.Y(n_456)
);

CKINVDCx11_ASAP7_75t_R g457 ( 
.A(n_401),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_367),
.B(n_369),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_383),
.A2(n_348),
.B1(n_374),
.B2(n_389),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_401),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_354),
.A2(n_382),
.B1(n_395),
.B2(n_391),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_423),
.A2(n_397),
.B(n_405),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_380),
.Y(n_469)
);

AOI221xp5_ASAP7_75t_L g470 ( 
.A1(n_417),
.A2(n_405),
.B1(n_380),
.B2(n_409),
.C(n_411),
.Y(n_470)
);

AOI21xp33_ASAP7_75t_L g471 ( 
.A1(n_440),
.A2(n_395),
.B(n_380),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_423),
.A2(n_409),
.B(n_411),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_449),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_427),
.B(n_442),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_413),
.A2(n_412),
.B(n_416),
.C(n_436),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_412),
.B(n_425),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_424),
.A2(n_456),
.B1(n_463),
.B2(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_451),
.B1(n_422),
.B2(n_464),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_425),
.A2(n_448),
.B(n_415),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_433),
.A2(n_420),
.B(n_435),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_421),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_434),
.B(n_444),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_465),
.A2(n_418),
.B(n_466),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_421),
.A2(n_464),
.B1(n_460),
.B2(n_418),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_454),
.Y(n_490)
);

AOI21xp33_ASAP7_75t_L g491 ( 
.A1(n_444),
.A2(n_447),
.B(n_452),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_422),
.B(n_447),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_431),
.A2(n_443),
.B(n_459),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_446),
.B1(n_441),
.B2(n_453),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_458),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_432),
.A2(n_419),
.B(n_467),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_437),
.A2(n_441),
.B1(n_446),
.B2(n_453),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_458),
.A2(n_459),
.B(n_450),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

AOI222xp33_ASAP7_75t_L g502 ( 
.A1(n_426),
.A2(n_438),
.B1(n_457),
.B2(n_439),
.C1(n_454),
.C2(n_419),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_472),
.A2(n_450),
.B(n_467),
.Y(n_503)
);

OAI31xp33_ASAP7_75t_L g504 ( 
.A1(n_471),
.A2(n_426),
.A3(n_454),
.B(n_428),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

OAI211xp5_ASAP7_75t_SL g506 ( 
.A1(n_491),
.A2(n_428),
.B(n_430),
.C(n_438),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_497),
.A2(n_432),
.B(n_419),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_439),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

OAI221xp5_ASAP7_75t_L g512 ( 
.A1(n_488),
.A2(n_429),
.B1(n_430),
.B2(n_432),
.C(n_481),
.Y(n_512)
);

NOR2x1_ASAP7_75t_SL g513 ( 
.A(n_499),
.B(n_429),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_492),
.B1(n_482),
.B2(n_483),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_469),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_496),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_490),
.A2(n_474),
.B1(n_486),
.B2(n_502),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_490),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_495),
.A2(n_498),
.B1(n_470),
.B2(n_490),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_475),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_501),
.B1(n_475),
.B2(n_479),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_484),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_510),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_501),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_512),
.A2(n_485),
.B1(n_480),
.B2(n_500),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_507),
.B(n_479),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_516),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_484),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_473),
.C(n_484),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_476),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_505),
.Y(n_533)
);

NAND2x1_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_480),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_520),
.Y(n_535)
);

NAND4xp25_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_504),
.C(n_514),
.D(n_517),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_533),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_534),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_509),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_528),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_522),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_511),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_513),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_526),
.C(n_531),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_530),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_519),
.B1(n_523),
.B2(n_534),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_536),
.A2(n_519),
.B(n_518),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_541),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_525),
.C(n_521),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_537),
.A2(n_509),
.B(n_523),
.C(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_545),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_549),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_552),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_551),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_550),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_557),
.A2(n_547),
.B(n_546),
.Y(n_558)
);

OAI322xp33_ASAP7_75t_L g559 ( 
.A1(n_553),
.A2(n_546),
.A3(n_541),
.B1(n_542),
.B2(n_511),
.C1(n_538),
.C2(n_524),
.Y(n_559)
);

AOI211xp5_ASAP7_75t_L g560 ( 
.A1(n_554),
.A2(n_556),
.B(n_555),
.C(n_542),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_555),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_538),
.B1(n_554),
.B2(n_530),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_538),
.C(n_509),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_560),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_563),
.B(n_562),
.C(n_559),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_R g566 ( 
.A1(n_565),
.A2(n_513),
.B1(n_509),
.B2(n_508),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_565),
.A2(n_510),
.B1(n_468),
.B2(n_503),
.Y(n_567)
);

NAND4xp25_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_566),
.C(n_510),
.D(n_508),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_568),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_569),
.A2(n_510),
.B1(n_468),
.B2(n_494),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_570),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_503),
.B(n_494),
.Y(n_572)
);


endmodule