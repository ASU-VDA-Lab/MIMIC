module fake_netlist_1_12293_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_9), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_7), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
NOR3xp33_ASAP7_75t_L g24 ( .A(n_16), .B(n_0), .C(n_1), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_20), .B(n_1), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_17), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_17), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_27) );
OAI21x1_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_21), .B(n_20), .Y(n_28) );
OA21x2_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_22), .B(n_19), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_24), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_30), .Y(n_34) );
OAI221xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_27), .B1(n_30), .B2(n_29), .C(n_31), .Y(n_35) );
NAND3xp33_ASAP7_75t_SL g36 ( .A(n_35), .B(n_18), .C(n_33), .Y(n_36) );
OAI31xp33_ASAP7_75t_SL g37 ( .A1(n_34), .A2(n_29), .A3(n_4), .B(n_5), .Y(n_37) );
AOI221xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_23), .B1(n_21), .B2(n_6), .C(n_3), .Y(n_38) );
NAND2x1p5_ASAP7_75t_L g39 ( .A(n_37), .B(n_23), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
AOI21xp33_ASAP7_75t_L g41 ( .A1(n_36), .A2(n_23), .B(n_5), .Y(n_41) );
INVx2_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_39), .Y(n_43) );
OAI22xp5_ASAP7_75t_SL g44 ( .A1(n_43), .A2(n_40), .B1(n_23), .B2(n_41), .Y(n_44) );
AOI322xp5_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_42), .A3(n_11), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_8), .Y(n_45) );
endmodule