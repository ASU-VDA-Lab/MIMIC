module fake_jpeg_129_n_141 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_42),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_6),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_29),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_63),
.C(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_60),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_31),
.B1(n_43),
.B2(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_14),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_25),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_82),
.B(n_61),
.Y(n_85)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_64),
.B1(n_47),
.B2(n_54),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_14),
.B(n_1),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_96),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_59),
.B1(n_64),
.B2(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_49),
.B1(n_65),
.B2(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_56),
.C(n_65),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_72),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_73),
.B(n_83),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_85),
.B1(n_95),
.B2(n_94),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_92),
.B(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_96),
.C(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_107),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_116),
.B1(n_106),
.B2(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_94),
.B1(n_86),
.B2(n_98),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_108),
.B(n_79),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_104),
.A3(n_106),
.B1(n_108),
.B2(n_107),
.C(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_124),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_79),
.C(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_118),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_65),
.B1(n_2),
.B2(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_131),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_7),
.B(n_9),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_130),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_120),
.A3(n_121),
.B1(n_126),
.B2(n_125),
.C1(n_10),
.C2(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_135),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_134),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

AOI21x1_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_0),
.B(n_2),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_137),
.Y(n_141)
);


endmodule