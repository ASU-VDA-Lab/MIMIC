module fake_ariane_2455_n_33 (n_8, n_3, n_2, n_11, n_7, n_5, n_1, n_0, n_12, n_6, n_9, n_4, n_10, n_33);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_5;
input n_1;
input n_0;
input n_12;
input n_6;
input n_9;
input n_4;
input n_10;

output n_33;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_27;
wire n_29;
wire n_17;
wire n_18;
wire n_32;
wire n_28;
wire n_26;
wire n_14;
wire n_19;
wire n_30;
wire n_31;
wire n_16;
wire n_15;
wire n_21;
wire n_23;
wire n_25;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_0),
.A2(n_2),
.B1(n_10),
.B2(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_19),
.Y(n_23)
);

AO21x2_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_16),
.B(n_17),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_18),
.B1(n_15),
.B2(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_18),
.B1(n_15),
.B2(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_23),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_24),
.Y(n_29)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_28),
.A3(n_23),
.B1(n_15),
.B2(n_1),
.C1(n_4),
.C2(n_2),
.Y(n_30)
);

AO22x2_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_1),
.B1(n_7),
.B2(n_12),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_31),
.Y(n_33)
);


endmodule