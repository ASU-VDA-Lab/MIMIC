module fake_jpeg_15748_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_4),
.B(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_60),
.B1(n_55),
.B2(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_57),
.B1(n_61),
.B2(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_49),
.B1(n_45),
.B2(n_51),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_53),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_99)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_64),
.B1(n_49),
.B2(n_48),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_90),
.B1(n_95),
.B2(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_53),
.C(n_58),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_7),
.C(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_72),
.Y(n_87)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_89),
.B(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_82),
.B1(n_54),
.B2(n_75),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_96),
.Y(n_106)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_25),
.B1(n_41),
.B2(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_1),
.Y(n_96)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_27),
.B1(n_10),
.B2(n_11),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_8),
.B1(n_22),
.B2(n_23),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_30),
.C(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_114),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_99),
.B(n_97),
.C(n_93),
.D(n_18),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_112),
.B(n_115),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_99),
.B(n_13),
.C(n_17),
.D(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_101),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_107),
.B1(n_103),
.B2(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_119),
.Y(n_123)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_108),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_124),
.C(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_122),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_126),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_121),
.B(n_31),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_28),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_32),
.B(n_33),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_34),
.B(n_35),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_102),
.Y(n_136)
);


endmodule