module fake_jpeg_28396_n_79 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_1),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_56),
.B1(n_58),
.B2(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_35),
.C(n_13),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_12),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_14),
.B1(n_29),
.B2(n_5),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_65),
.C(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_60),
.B(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_71),
.CI(n_4),
.CON(n_74),
.SN(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_3),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_74),
.C(n_4),
.Y(n_76)
);

AOI332xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_3),
.A3(n_6),
.B1(n_8),
.B2(n_10),
.B3(n_11),
.C1(n_21),
.C2(n_22),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_54),
.C(n_57),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_26),
.A3(n_27),
.B1(n_30),
.B2(n_59),
.C1(n_66),
.C2(n_75),
.Y(n_79)
);


endmodule