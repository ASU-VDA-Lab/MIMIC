module fake_jpeg_2975_n_548 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_548);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_548;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_61),
.B(n_69),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_63),
.Y(n_159)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_9),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_24),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_70),
.B(n_92),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_81),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_19),
.A2(n_57),
.B(n_38),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_122),
.B(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_48),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_93),
.Y(n_165)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx9p33_ASAP7_75t_R g179 ( 
.A(n_95),
.Y(n_179)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_28),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_111),
.Y(n_138)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_105),
.Y(n_166)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_35),
.B(n_8),
.Y(n_111)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_116),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_35),
.B(n_10),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_40),
.B(n_10),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_42),
.Y(n_143)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_44),
.B(n_7),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_123),
.B(n_18),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_19),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_19),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_66),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_128),
.B(n_142),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_33),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_131),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_60),
.A2(n_37),
.B1(n_32),
.B2(n_43),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_135),
.A2(n_137),
.B1(n_174),
.B2(n_197),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_72),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_143),
.B(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_43),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_76),
.B(n_27),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_190),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_73),
.A2(n_32),
.B1(n_42),
.B2(n_27),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_167),
.A2(n_63),
.B1(n_45),
.B2(n_2),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_68),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_85),
.A2(n_42),
.B1(n_33),
.B2(n_57),
.Y(n_170)
);

OA22x2_ASAP7_75t_SL g228 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_62),
.A2(n_23),
.B1(n_41),
.B2(n_38),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_189),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_93),
.A2(n_51),
.B1(n_49),
.B2(n_57),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_194),
.B1(n_206),
.B2(n_131),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_82),
.B(n_41),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_77),
.B(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_74),
.B(n_41),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_200),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_51),
.B1(n_38),
.B2(n_23),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_58),
.B(n_23),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_196),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_95),
.A2(n_26),
.B(n_54),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_64),
.A2(n_56),
.B1(n_54),
.B2(n_52),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_95),
.A2(n_56),
.B(n_54),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_0),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_99),
.B(n_52),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_209),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_102),
.B(n_13),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_124),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_205),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_90),
.A2(n_56),
.B1(n_52),
.B2(n_45),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_125),
.A2(n_12),
.B(n_18),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_67),
.B1(n_97),
.B2(n_105),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_213),
.A2(n_220),
.B1(n_226),
.B2(n_257),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_115),
.A3(n_121),
.B1(n_112),
.B2(n_107),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_217),
.A2(n_274),
.B(n_228),
.C(n_235),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_130),
.A2(n_98),
.B1(n_88),
.B2(n_113),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_218),
.A2(n_245),
.B1(n_269),
.B2(n_237),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_141),
.A2(n_108),
.B1(n_104),
.B2(n_100),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_161),
.A2(n_117),
.B1(n_116),
.B2(n_94),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_128),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

AO22x2_ASAP7_75t_L g294 ( 
.A1(n_228),
.A2(n_154),
.B1(n_173),
.B2(n_210),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_151),
.B(n_3),
.C(n_5),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_250),
.C(n_238),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_5),
.B1(n_6),
.B2(n_14),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_234),
.A2(n_240),
.B1(n_251),
.B2(n_226),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_236),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_177),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_237),
.A2(n_255),
.B1(n_258),
.B2(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_163),
.A2(n_5),
.B1(n_6),
.B2(n_14),
.Y(n_240)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_243),
.A2(n_252),
.B1(n_259),
.B2(n_260),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_138),
.A2(n_16),
.B1(n_18),
.B2(n_136),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_131),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_247),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_129),
.Y(n_248)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_16),
.C(n_158),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_180),
.A2(n_16),
.B1(n_191),
.B2(n_166),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_131),
.A2(n_133),
.B1(n_171),
.B2(n_202),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_169),
.A2(n_172),
.B1(n_178),
.B2(n_152),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_256),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_169),
.A2(n_178),
.B1(n_172),
.B2(n_181),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_152),
.A2(n_133),
.B1(n_180),
.B2(n_157),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_133),
.A2(n_171),
.B1(n_201),
.B2(n_157),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_157),
.A2(n_198),
.B1(n_175),
.B2(n_139),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_170),
.B(n_183),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_264),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_185),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_145),
.B(n_182),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_271),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_188),
.A2(n_182),
.B1(n_211),
.B2(n_153),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_198),
.A2(n_139),
.B1(n_175),
.B2(n_188),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_270),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_127),
.B(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_127),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_181),
.A2(n_187),
.B1(n_207),
.B2(n_146),
.Y(n_273)
);

AO21x2_ASAP7_75t_SL g320 ( 
.A1(n_273),
.A2(n_231),
.B(n_249),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_165),
.B(n_144),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_275),
.Y(n_323)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_SL g276 ( 
.A(n_159),
.B(n_150),
.C(n_148),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_276),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_144),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_153),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_279),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_146),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_164),
.A2(n_162),
.B1(n_210),
.B2(n_173),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_148),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_214),
.B(n_208),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_316),
.C(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_239),
.A2(n_208),
.B1(n_150),
.B2(n_147),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_299),
.B1(n_301),
.B2(n_306),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_294),
.B(n_314),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_160),
.B1(n_173),
.B2(n_210),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_297),
.A2(n_318),
.B1(n_324),
.B2(n_277),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_216),
.A2(n_126),
.B1(n_147),
.B2(n_160),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_126),
.B1(n_160),
.B2(n_229),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_303),
.B1(n_325),
.B2(n_335),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_220),
.B1(n_213),
.B2(n_229),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_214),
.A2(n_230),
.B1(n_242),
.B2(n_244),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_331),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_222),
.A2(n_268),
.B1(n_242),
.B2(n_246),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_268),
.A2(n_228),
.B(n_212),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_328),
.B(n_329),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_268),
.A2(n_225),
.B1(n_224),
.B2(n_258),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_313),
.A2(n_286),
.B1(n_324),
.B2(n_285),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_221),
.B(n_228),
.C(n_219),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_315),
.B(n_330),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_223),
.Y(n_316)
);

AO21x2_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_332),
.B(n_325),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_321),
.A2(n_302),
.B1(n_296),
.B2(n_291),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_271),
.A2(n_217),
.B1(n_279),
.B2(n_255),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_273),
.B1(n_248),
.B2(n_227),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_273),
.B(n_250),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_282),
.B(n_236),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_233),
.A2(n_272),
.B(n_253),
.C(n_247),
.Y(n_330)
);

AOI32xp33_ASAP7_75t_L g331 ( 
.A1(n_281),
.A2(n_254),
.A3(n_267),
.B1(n_241),
.B2(n_283),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_257),
.A2(n_256),
.B1(n_277),
.B2(n_215),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_265),
.A2(n_261),
.B1(n_239),
.B2(n_268),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_214),
.C(n_216),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_317),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_343),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_305),
.B(n_303),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_340),
.B(n_358),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_342),
.B1(n_353),
.B2(n_363),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_316),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_350),
.Y(n_393)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_302),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_291),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_371),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_301),
.A2(n_296),
.B1(n_314),
.B2(n_300),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_292),
.B(n_304),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_359),
.C(n_362),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_315),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_361),
.Y(n_404)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_288),
.B(n_284),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_306),
.B(n_288),
.C(n_308),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_284),
.B(n_330),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_284),
.B(n_313),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_286),
.A2(n_328),
.B1(n_289),
.B2(n_320),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_312),
.B(n_335),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_365),
.B(n_287),
.Y(n_382)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_318),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_370),
.C(n_374),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_312),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_293),
.C(n_310),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_290),
.B(n_310),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_294),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_294),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_289),
.C(n_290),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_287),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_326),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_374),
.A2(n_320),
.B1(n_294),
.B2(n_332),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_379),
.A2(n_408),
.B1(n_342),
.B2(n_372),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_350),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_398),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_356),
.C(n_377),
.Y(n_411)
);

XNOR2x2_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_294),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_386),
.A2(n_394),
.B(n_399),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_331),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_399),
.B(n_394),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_309),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_359),
.C(n_338),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_349),
.A2(n_376),
.B(n_375),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_311),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_352),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_345),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_311),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_403),
.B(n_375),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_309),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_406),
.C(n_362),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_307),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_363),
.A2(n_326),
.B1(n_322),
.B2(n_327),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_409),
.B(n_322),
.Y(n_433)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_383),
.A2(n_353),
.B1(n_342),
.B2(n_349),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_412),
.A2(n_414),
.B1(n_416),
.B2(n_423),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_418),
.C(n_428),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_367),
.B1(n_342),
.B2(n_357),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_381),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_424),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_402),
.A2(n_342),
.B1(n_376),
.B2(n_348),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_387),
.A2(n_348),
.B1(n_368),
.B2(n_373),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_398),
.B(n_340),
.Y(n_425)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_344),
.Y(n_427)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_343),
.C(n_370),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_366),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_435),
.C(n_407),
.Y(n_443)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_433),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_410),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_391),
.C(n_401),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_436),
.A2(n_439),
.B1(n_390),
.B2(n_410),
.Y(n_463)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_385),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_392),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_438),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_380),
.B(n_389),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_445),
.C(n_454),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_406),
.C(n_407),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_383),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_462),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_406),
.C(n_378),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_455),
.B(n_382),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_418),
.C(n_428),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_399),
.C(n_403),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_438),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_461),
.B(n_417),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_404),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_463),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_404),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_439),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_466),
.B(n_469),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_448),
.A2(n_416),
.B1(n_414),
.B2(n_412),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_468),
.A2(n_448),
.B1(n_424),
.B2(n_449),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_456),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_450),
.B(n_425),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_470),
.B(n_475),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_429),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_476),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_464),
.A2(n_411),
.B1(n_423),
.B2(n_421),
.Y(n_472)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_478),
.C(n_481),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_389),
.C(n_403),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_482),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_434),
.C(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_420),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_486),
.C(n_442),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_456),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_484),
.Y(n_498)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_452),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_436),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_468),
.A2(n_449),
.B1(n_440),
.B2(n_460),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_490),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_447),
.B(n_441),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_470),
.A2(n_440),
.B1(n_387),
.B2(n_457),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_491),
.A2(n_419),
.B1(n_444),
.B2(n_482),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_441),
.B(n_463),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_501),
.Y(n_509)
);

OAI321xp33_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_422),
.A3(n_415),
.B1(n_446),
.B2(n_433),
.C(n_390),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_474),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_504),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_481),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_471),
.C(n_474),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_506),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_467),
.C(n_486),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_507),
.A2(n_508),
.B1(n_485),
.B2(n_488),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_467),
.C(n_454),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_512),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_478),
.C(n_462),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_483),
.C(n_476),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_444),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_495),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_515),
.B(n_518),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_502),
.A2(n_492),
.B1(n_487),
.B2(n_489),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_516),
.B(n_521),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_509),
.A2(n_491),
.B1(n_387),
.B2(n_379),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_520),
.B(n_499),
.Y(n_526)
);

AOI21x1_ASAP7_75t_SL g520 ( 
.A1(n_509),
.A2(n_488),
.B(n_495),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_465),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_499),
.B(n_498),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_510),
.B(n_397),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_528),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_523),
.A2(n_500),
.B(n_506),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_527),
.A2(n_532),
.B(n_519),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_480),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_530),
.B(n_531),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_479),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_522),
.B(n_393),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_525),
.C(n_521),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_535),
.A2(n_536),
.B(n_539),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_533),
.A2(n_520),
.B(n_515),
.Y(n_536)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_537),
.Y(n_541)
);

A2O1A1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_533),
.A2(n_518),
.B(n_516),
.C(n_393),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_534),
.A2(n_452),
.B(n_437),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_431),
.B(n_395),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_538),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_397),
.Y(n_545)
);

AOI322xp5_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_545),
.A3(n_388),
.B1(n_541),
.B2(n_540),
.C1(n_395),
.C2(n_432),
.Y(n_546)
);

AOI21x1_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_388),
.B(n_408),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_390),
.Y(n_548)
);


endmodule