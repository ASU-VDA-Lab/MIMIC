module fake_jpeg_25537_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_18),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_25),
.B(n_24),
.C(n_15),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_37),
.B(n_39),
.C(n_45),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_17),
.B1(n_26),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_13),
.B1(n_18),
.B2(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_17),
.B1(n_26),
.B2(n_23),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_13),
.B1(n_24),
.B2(n_25),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_56),
.Y(n_80)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_59),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_18),
.A3(n_13),
.B1(n_15),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_36),
.B1(n_15),
.B2(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_22),
.B1(n_27),
.B2(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_14),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_71),
.B1(n_81),
.B2(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_47),
.B1(n_43),
.B2(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_63),
.B(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_2),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_10),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_51),
.B1(n_62),
.B2(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_30),
.B1(n_40),
.B2(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_62),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_30),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_72),
.B1(n_74),
.B2(n_66),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_77),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_40),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_68),
.C(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_101),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_2),
.B(n_3),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_70),
.B1(n_80),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_85),
.B1(n_91),
.B2(n_84),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_80),
.B1(n_66),
.B2(n_4),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_102),
.B1(n_97),
.B2(n_99),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_114),
.B(n_120),
.C(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_96),
.C(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_111),
.B1(n_106),
.B2(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_116),
.B(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.C(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_7),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_6),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_6),
.B1(n_7),
.B2(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_129),
.Y(n_137)
);


endmodule