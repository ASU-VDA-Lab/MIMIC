module fake_jpeg_16345_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_60),
.B1(n_43),
.B2(n_52),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_80),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_48),
.C(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_60),
.B1(n_52),
.B2(n_43),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_61),
.B1(n_59),
.B2(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_1),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_44),
.B1(n_49),
.B2(n_56),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_23),
.B1(n_22),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_76),
.B1(n_78),
.B2(n_4),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_61),
.B1(n_46),
.B2(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_97),
.Y(n_103)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_95),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_74),
.B1(n_71),
.B2(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_96),
.B1(n_90),
.B2(n_91),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_57),
.C(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_5),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_85),
.B1(n_83),
.B2(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_25),
.B1(n_36),
.B2(n_35),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_6),
.B(n_8),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_102),
.C(n_106),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_118),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_103),
.C(n_107),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_111),
.B1(n_116),
.B2(n_117),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_86),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_120),
.B1(n_113),
.B2(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_122),
.B1(n_123),
.B2(n_26),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_18),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_21),
.A3(n_30),
.B1(n_29),
.B2(n_28),
.C1(n_27),
.C2(n_32),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_8),
.B(n_9),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_11),
.C(n_13),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_11),
.Y(n_135)
);


endmodule