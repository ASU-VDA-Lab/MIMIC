module real_jpeg_26079_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_1),
.A2(n_62),
.B(n_162),
.C(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_57),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_59),
.B(n_73),
.C(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_27),
.C(n_38),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_1),
.B(n_127),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_1),
.B(n_11),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_1),
.B(n_36),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_31),
.B1(n_58),
.B2(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_31),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_65),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_11),
.Y(n_167)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_274),
.B1(n_288),
.B2(n_289),
.Y(n_13)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_14),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_131),
.B(n_273),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_108),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_16),
.B(n_108),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_89),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_17),
.B(n_82),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_48),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_18),
.B(n_49),
.C(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_19),
.B(n_34),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_20),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_21),
.B(n_218),
.Y(n_223)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_22),
.A2(n_24),
.B(n_32),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_24),
.B(n_32),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_27),
.B(n_229),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_28),
.A2(n_59),
.B(n_61),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_28),
.A2(n_41),
.B(n_75),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_29),
.A2(n_93),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_29),
.B(n_223),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_32),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_32),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B(n_44),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_35),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_35),
.A2(n_86),
.B(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_36),
.B(n_193),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_46)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_42),
.B(n_206),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_44),
.B(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_45),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_68),
.B2(n_69),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_52),
.B(n_66),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_53),
.Y(n_163)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_64),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_57),
.B(n_105),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_73),
.B2(n_75),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_63),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_70),
.B(n_153),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_70),
.A2(n_78),
.B(n_126),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_71),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_79),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_72),
.B(n_101),
.Y(n_155)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_77),
.B(n_146),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_79),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_88),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_83),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_83),
.A2(n_88),
.B1(n_188),
.B2(n_245),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_83),
.A2(n_112),
.B(n_114),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_87),
.B(n_192),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_90),
.A2(n_91),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_95),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_98),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_100),
.A2(n_102),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_102),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_130),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_119),
.B2(n_120),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_110),
.B(n_120),
.C(n_130),
.Y(n_286)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_125),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_129),
.B(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_268),
.B(n_272),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_181),
.B(n_254),
.C(n_267),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_169),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_134),
.B(n_169),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_150),
.B2(n_168),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_148),
.B2(n_149),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_137),
.B(n_149),
.C(n_168),
.Y(n_255)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_140),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_141),
.B(n_157),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_142),
.A2(n_143),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_152),
.B(n_159),
.C(n_160),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_171),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_176),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_253),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_197),
.B(n_252),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_184),
.B(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_185),
.B(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_190),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_188),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_247),
.B(n_251),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_238),
.B(n_246),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_220),
.B(n_237),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_201),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_214),
.B2(n_219),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_213),
.C(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_226),
.B(n_236),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_232),
.B(n_235),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_243),
.C(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_264),
.B2(n_265),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_287),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_286),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);


endmodule