module fake_jpeg_3034_n_366 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_45),
.Y(n_124)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_47),
.B(n_53),
.Y(n_139)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_48),
.Y(n_146)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_14),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_27),
.A2(n_33),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_61),
.B(n_66),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_12),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_85),
.Y(n_112)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_99),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_23),
.B(n_10),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_90),
.Y(n_132)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_18),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_94),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_96),
.Y(n_140)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_50),
.B1(n_55),
.B2(n_72),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_111),
.A2(n_122),
.B1(n_151),
.B2(n_79),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_44),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_66),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_64),
.A2(n_44),
.B1(n_43),
.B2(n_34),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_34),
.C(n_31),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_127),
.B(n_124),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_53),
.A2(n_31),
.B(n_2),
.C(n_3),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_137),
.B(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_121),
.B1(n_140),
.B2(n_123),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_51),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_107),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_155),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_90),
.B1(n_108),
.B2(n_109),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g223 ( 
.A1(n_157),
.A2(n_194),
.B(n_107),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_158),
.A2(n_106),
.B1(n_125),
.B2(n_133),
.Y(n_222)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_171),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_96),
.B1(n_95),
.B2(n_93),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_170),
.B1(n_185),
.B2(n_189),
.Y(n_203)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_92),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_59),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_62),
.B1(n_83),
.B2(n_56),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_183),
.B1(n_150),
.B2(n_103),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_176),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_70),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_187),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_73),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_122),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_139),
.B(n_9),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_184),
.Y(n_196)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_109),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_191),
.Y(n_219)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_190),
.A2(n_147),
.B1(n_135),
.B2(n_146),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_138),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_119),
.B(n_138),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_193),
.B1(n_124),
.B2(n_128),
.Y(n_208)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_141),
.A2(n_144),
.B1(n_130),
.B2(n_134),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_152),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_134),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_205),
.C(n_187),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_214),
.B1(n_221),
.B2(n_194),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_148),
.B1(n_131),
.B2(n_126),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_157),
.A2(n_118),
.B1(n_131),
.B2(n_126),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_148),
.B1(n_118),
.B2(n_147),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_163),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_186),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_166),
.Y(n_232)
);

INVx2_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_247),
.B(n_248),
.C(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_237),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_243),
.Y(n_249)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_157),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_182),
.Y(n_238)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_183),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_189),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_219),
.B1(n_225),
.B2(n_196),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_175),
.B1(n_187),
.B2(n_194),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_223),
.B1(n_214),
.B2(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_175),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_238),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_217),
.C(n_198),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_260),
.C(n_243),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_268),
.B1(n_269),
.B2(n_235),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_217),
.C(n_203),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_223),
.B(n_204),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_248),
.B(n_247),
.Y(n_271)
);

OAI22x1_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_223),
.B1(n_221),
.B2(n_160),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_233),
.B(n_248),
.C(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_196),
.B1(n_224),
.B2(n_202),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_229),
.A2(n_202),
.B1(n_161),
.B2(n_197),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_276),
.B1(n_286),
.B2(n_255),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_281),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_229),
.B1(n_228),
.B2(n_245),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_282),
.B1(n_285),
.B2(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_251),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_256),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_233),
.B1(n_244),
.B2(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_258),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_264),
.B(n_236),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_257),
.B(n_227),
.Y(n_284)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_251),
.B(n_261),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_242),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_240),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_253),
.C(n_240),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_249),
.A2(n_246),
.B1(n_238),
.B2(n_230),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_259),
.B1(n_262),
.B2(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_290),
.C(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_255),
.C(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_265),
.B1(n_276),
.B2(n_246),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_295),
.B1(n_305),
.B2(n_275),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_266),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_286),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_267),
.C(n_226),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_267),
.C(n_263),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_275),
.C(n_281),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_317),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_320),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_270),
.B1(n_283),
.B2(n_263),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_278),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_318),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.C(n_305),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_263),
.C(n_197),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_276),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_325),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_309),
.C(n_319),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_298),
.Y(n_330)
);

OAI221xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_304),
.B1(n_295),
.B2(n_309),
.C(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_318),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_334),
.Y(n_344)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_324),
.B1(n_327),
.B2(n_316),
.C(n_297),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_236),
.B1(n_174),
.B2(n_165),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_307),
.B1(n_317),
.B2(n_297),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_335),
.B(n_336),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_297),
.B1(n_276),
.B2(n_200),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_340),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_200),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_326),
.C(n_216),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_343),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_326),
.C(n_216),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_210),
.C(n_276),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_345),
.B(n_347),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_210),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_162),
.C(n_155),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_335),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_354),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_346),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_351),
.A2(n_352),
.B1(n_102),
.B2(n_128),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_180),
.C(n_156),
.Y(n_354)
);

AOI31xp67_ASAP7_75t_L g356 ( 
.A1(n_354),
.A2(n_342),
.A3(n_185),
.B(n_102),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_179),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_358),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_349),
.C(n_352),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_360),
.A2(n_129),
.B(n_125),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.C(n_359),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g363 ( 
.A1(n_361),
.A2(n_135),
.B(n_102),
.Y(n_363)
);

O2A1O1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_364),
.A2(n_106),
.B(n_114),
.C(n_159),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_365),
.Y(n_366)
);


endmodule