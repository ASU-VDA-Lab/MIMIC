module fake_ariane_3353_n_1667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1667;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_63),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_43),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_54),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_27),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_0),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_64),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_81),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_32),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_62),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_74),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_34),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_10),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_42),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_102),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_32),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_58),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_26),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_37),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_46),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_31),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_57),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_90),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_51),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_33),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_15),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_53),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_69),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_16),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_137),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_30),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_80),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_72),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_56),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_66),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_129),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_21),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_13),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_18),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_88),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_7),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_17),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_50),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_5),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_42),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_46),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_36),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_99),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_130),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_95),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_44),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_92),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_100),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_97),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_111),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_25),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_89),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_107),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_40),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_39),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_101),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_12),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_22),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_91),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_61),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_116),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_113),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_40),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_117),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_45),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_134),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_140),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_93),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_114),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_77),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_55),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_28),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_20),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_52),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_248),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_161),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_162),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_165),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_225),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_165),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_R g309 ( 
.A(n_153),
.B(n_70),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_248),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_270),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_2),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_276),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_152),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_165),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_185),
.B(n_4),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_185),
.B(n_5),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_207),
.B(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_295),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_158),
.B(n_6),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_207),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_182),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_164),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_183),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_186),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_241),
.B(n_8),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_155),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_188),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_241),
.B(n_8),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_269),
.B(n_9),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_269),
.B(n_10),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_288),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_279),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_279),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_179),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_193),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_265),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_179),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_221),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_200),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_155),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_151),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_201),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_157),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_151),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_168),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_202),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_203),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_187),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_168),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_209),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_157),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_174),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_174),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_214),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_215),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_178),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_217),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_234),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_152),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_208),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_271),
.B(n_159),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_160),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_175),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_300),
.B(n_271),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_301),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_302),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_381),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_306),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_323),
.A2(n_189),
.B(n_176),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_307),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_307),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_308),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_310),
.B(n_198),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_336),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_329),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_315),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_305),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_190),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_360),
.A2(n_195),
.B(n_191),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_322),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_364),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_341),
.B(n_184),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_363),
.B(n_208),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_314),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_364),
.B(n_197),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_318),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_324),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_353),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_358),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_355),
.B(n_250),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_334),
.B(n_198),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_368),
.A2(n_285),
.B(n_257),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_361),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_354),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_365),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_366),
.B(n_152),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_303),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_373),
.B(n_226),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_380),
.B(n_371),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_400),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_359),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_436),
.B(n_374),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_384),
.A2(n_313),
.B1(n_344),
.B2(n_321),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_383),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_316),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_384),
.A2(n_340),
.B1(n_311),
.B2(n_345),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_384),
.A2(n_311),
.B1(n_319),
.B2(n_320),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_384),
.A2(n_309),
.B1(n_378),
.B2(n_376),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_440),
.B(n_319),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_448),
.B(n_320),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_451),
.B(n_345),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_400),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_348),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_454),
.B(n_346),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_404),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_400),
.B(n_371),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_383),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_441),
.A2(n_160),
.B1(n_258),
.B2(n_169),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_326),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_393),
.A2(n_331),
.B1(n_367),
.B2(n_247),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_454),
.B(n_257),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_372),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_441),
.B(n_153),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_169),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_455),
.B(n_379),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_387),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_450),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_445),
.B(n_285),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_259),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_352),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_397),
.B(n_154),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_402),
.B(n_405),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_449),
.B(n_259),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_421),
.B(n_177),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_372),
.Y(n_515)
);

AND3x2_ASAP7_75t_L g516 ( 
.A(n_431),
.B(n_235),
.C(n_194),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_393),
.B(n_416),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_439),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_375),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_393),
.B(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_392),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_431),
.B(n_154),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_388),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_418),
.A2(n_218),
.B1(n_291),
.B2(n_280),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_427),
.B(n_259),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_398),
.B(n_177),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_377),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_401),
.B(n_156),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_204),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_394),
.B(n_205),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_406),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_385),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_413),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_409),
.B(n_420),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_395),
.B(n_272),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_425),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_396),
.B(n_352),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_396),
.B(n_259),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_399),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_427),
.B(n_356),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_399),
.B(n_156),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_403),
.B(n_163),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_403),
.B(n_163),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_407),
.B(n_356),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_411),
.B(n_166),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_411),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_166),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_433),
.B(n_167),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_415),
.B(n_210),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_415),
.B(n_417),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_427),
.A2(n_251),
.B1(n_192),
.B2(n_196),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_417),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_419),
.B(n_211),
.C(n_298),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_419),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_427),
.B(n_167),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_429),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_446),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_SL g571 ( 
.A1(n_429),
.A2(n_231),
.B(n_199),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_427),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_434),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_406),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_442),
.B(n_170),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_425),
.B(n_170),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_425),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_408),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_443),
.B(n_171),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_443),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_408),
.B(n_443),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_414),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_414),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_414),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_443),
.B(n_172),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_443),
.B(n_172),
.Y(n_591)
);

AND2x2_ASAP7_75t_SL g592 ( 
.A(n_443),
.B(n_228),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_386),
.B(n_357),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_386),
.B(n_212),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_386),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_492),
.B(n_514),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_462),
.B(n_173),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_476),
.B(n_246),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_496),
.B(n_173),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_460),
.B(n_253),
.C(n_255),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_503),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_482),
.Y(n_603)
);

NAND3xp33_ASAP7_75t_L g604 ( 
.A(n_470),
.B(n_255),
.C(n_258),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_464),
.B(n_180),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_512),
.B(n_261),
.C(n_274),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_489),
.B(n_180),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_465),
.B(n_181),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_503),
.B(n_261),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_476),
.B(n_236),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_471),
.B(n_181),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_496),
.B(n_254),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_274),
.C(n_275),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_459),
.B(n_262),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_237),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_505),
.A2(n_226),
.B1(n_250),
.B2(n_184),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_482),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_592),
.B(n_264),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_592),
.B(n_521),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_238),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_486),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_492),
.B(n_382),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_463),
.A2(n_275),
.B1(n_296),
.B2(n_297),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_493),
.B(n_264),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_478),
.B(n_273),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_521),
.B(n_273),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_521),
.B(n_292),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_239),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_514),
.B(n_382),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_500),
.B(n_243),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_533),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_488),
.B(n_244),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_486),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_508),
.B(n_250),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_535),
.B(n_245),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_505),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_498),
.B(n_252),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_508),
.B(n_357),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_494),
.B(n_296),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_456),
.B(n_266),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_297),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_505),
.A2(n_226),
.B1(n_224),
.B2(n_223),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_483),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_509),
.B(n_227),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_540),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_457),
.B(n_230),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_507),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_534),
.B(n_542),
.Y(n_654)
);

BUFx5_ASAP7_75t_L g655 ( 
.A(n_531),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_588),
.Y(n_656)
);

A2O1A1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_537),
.A2(n_232),
.B(n_278),
.C(n_287),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_457),
.B(n_293),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_511),
.A2(n_294),
.B(n_18),
.C(n_20),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_501),
.B(n_11),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_541),
.B(n_240),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_524),
.B(n_11),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_528),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_507),
.B(n_467),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_472),
.B(n_22),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_588),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_511),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_468),
.B(n_242),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_563),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_566),
.B(n_233),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_566),
.B(n_268),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_569),
.B(n_229),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_545),
.B(n_222),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_SL g675 ( 
.A(n_541),
.B(n_281),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_545),
.B(n_220),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_517),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_533),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_527),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_556),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_553),
.B(n_284),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_553),
.B(n_219),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_556),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_567),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_480),
.B(n_28),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_495),
.B(n_290),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_502),
.B(n_29),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_523),
.B(n_547),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_554),
.B(n_289),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_216),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_549),
.B(n_213),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_473),
.B(n_474),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_466),
.B(n_469),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

AND2x6_ASAP7_75t_SL g696 ( 
.A(n_504),
.B(n_29),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_550),
.B(n_206),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_552),
.B(n_412),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_466),
.B(n_412),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_481),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_573),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_555),
.B(n_412),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_573),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_574),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_574),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_412),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_484),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_461),
.B(n_412),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_593),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_469),
.B(n_412),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_530),
.A2(n_385),
.B1(n_406),
.B2(n_39),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_501),
.B(n_35),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_35),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_548),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_580),
.B(n_36),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_582),
.B(n_41),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_557),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_491),
.B(n_41),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_590),
.A2(n_406),
.B1(n_44),
.B2(n_43),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_559),
.B(n_406),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_475),
.B(n_68),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_595),
.A2(n_75),
.B(n_78),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_475),
.B(n_79),
.Y(n_725)
);

XNOR2xp5_ASAP7_75t_L g726 ( 
.A(n_516),
.B(n_82),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_475),
.B(n_86),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_557),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_544),
.B(n_87),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_518),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_544),
.B(n_103),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_557),
.B(n_104),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_490),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_577),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_497),
.B(n_149),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_565),
.B(n_106),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_497),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_662),
.A2(n_585),
.B(n_571),
.C(n_558),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_635),
.B(n_577),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_694),
.A2(n_479),
.B(n_477),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_694),
.A2(n_479),
.B(n_477),
.Y(n_741)
);

AO21x1_ASAP7_75t_L g742 ( 
.A1(n_722),
.A2(n_522),
.B(n_594),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_654),
.B(n_525),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_707),
.B(n_525),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_638),
.B(n_570),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_647),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_625),
.A2(n_714),
.B(n_632),
.C(n_719),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_596),
.Y(n_748)
);

OAI21xp33_ASAP7_75t_L g749 ( 
.A1(n_610),
.A2(n_591),
.B(n_578),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_662),
.A2(n_568),
.B(n_558),
.C(n_584),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_610),
.B(n_506),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_723),
.B(n_526),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_698),
.A2(n_583),
.B(n_584),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_702),
.A2(n_584),
.B(n_581),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_706),
.A2(n_581),
.B(n_564),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_722),
.A2(n_458),
.B(n_526),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_608),
.B(n_642),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_679),
.B(n_548),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_600),
.A2(n_568),
.B1(n_548),
.B2(n_526),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_725),
.A2(n_458),
.B(n_529),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_600),
.B(n_487),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_612),
.B(n_487),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_616),
.B(n_562),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_628),
.A2(n_519),
.B(n_506),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_627),
.B(n_529),
.Y(n_766)
);

INVx11_ASAP7_75t_L g767 ( 
.A(n_602),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_611),
.B(n_570),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_597),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_663),
.B(n_577),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_630),
.A2(n_575),
.B(n_551),
.C(n_538),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_597),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_649),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_629),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_678),
.A2(n_575),
.B(n_551),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_587),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_587),
.Y(n_777)
);

OAI321xp33_ASAP7_75t_L g778 ( 
.A1(n_616),
.A2(n_532),
.A3(n_546),
.B1(n_513),
.B2(n_587),
.C(n_572),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_597),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_711),
.A2(n_699),
.B(n_689),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_648),
.A2(n_532),
.B(n_539),
.C(n_572),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_575),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_605),
.B(n_572),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_615),
.B(n_539),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_727),
.A2(n_538),
.B(n_539),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_622),
.B(n_539),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_623),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_622),
.B(n_539),
.Y(n_789)
);

BUFx4f_ASAP7_75t_L g790 ( 
.A(n_728),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_637),
.A2(n_546),
.B1(n_513),
.B2(n_121),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_SL g792 ( 
.A(n_640),
.B(n_652),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_601),
.A2(n_598),
.B(n_636),
.C(n_641),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_709),
.A2(n_546),
.B(n_513),
.C(n_123),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_624),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_650),
.A2(n_546),
.B1(n_513),
.B2(n_128),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_710),
.B(n_546),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_715),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_692),
.A2(n_513),
.B(n_115),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_607),
.B(n_513),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_640),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_697),
.A2(n_673),
.B(n_671),
.Y(n_802)
);

CKINVDCx11_ASAP7_75t_R g803 ( 
.A(n_696),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_667),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_672),
.A2(n_138),
.B(n_139),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_599),
.B(n_715),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_648),
.A2(n_143),
.B1(n_147),
.B2(n_619),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_633),
.B(n_599),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_653),
.B(n_677),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_604),
.B(n_626),
.Y(n_810)
);

BUFx4f_ASAP7_75t_L g811 ( 
.A(n_732),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_736),
.B(n_680),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_681),
.A2(n_705),
.B(n_684),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_685),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_597),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_674),
.B(n_676),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_621),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_660),
.B(n_713),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_639),
.B(n_718),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_613),
.B(n_639),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_682),
.A2(n_683),
.B(n_606),
.C(n_619),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_695),
.A2(n_701),
.B(n_704),
.C(n_703),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_634),
.B(n_693),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_687),
.A2(n_690),
.B(n_691),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_670),
.B(n_634),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_659),
.A2(n_657),
.B(n_668),
.C(n_614),
.Y(n_826)
);

OR2x6_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_609),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_665),
.B(n_686),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_665),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_700),
.Y(n_830)
);

AND2x6_ASAP7_75t_L g831 ( 
.A(n_631),
.B(n_730),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_656),
.B(n_666),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_733),
.Y(n_833)
);

BUFx4_ASAP7_75t_SL g834 ( 
.A(n_688),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_643),
.B(n_646),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_646),
.B(n_693),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_675),
.B(n_686),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_708),
.A2(n_737),
.B(n_734),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_734),
.A2(n_735),
.B(n_620),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_631),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_631),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_712),
.A2(n_720),
.B1(n_664),
.B2(n_717),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_631),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_669),
.B(n_645),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_620),
.B(n_730),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_734),
.A2(n_644),
.B(n_651),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_730),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_651),
.A2(n_658),
.B(n_716),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_730),
.B(n_734),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_726),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_712),
.B(n_658),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_644),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_655),
.B(n_721),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_729),
.B(n_731),
.C(n_724),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_655),
.A2(n_694),
.B(n_698),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_655),
.A2(n_725),
.B(n_722),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_654),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_662),
.A2(n_460),
.B(n_714),
.C(n_648),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_603),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_654),
.B(n_464),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_694),
.A2(n_702),
.B(n_698),
.Y(n_861)
);

NOR2x1p5_ASAP7_75t_L g862 ( 
.A(n_602),
.B(n_503),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_600),
.A2(n_496),
.B1(n_612),
.B2(n_619),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_638),
.B(n_492),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_600),
.A2(n_496),
.B1(n_612),
.B2(n_460),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_694),
.A2(n_702),
.B(n_698),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_603),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_638),
.B(n_492),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_654),
.B(n_464),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_661),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_638),
.B(n_492),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_654),
.B(n_464),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_600),
.A2(n_496),
.B1(n_612),
.B2(n_460),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_735),
.A2(n_479),
.B(n_477),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_600),
.A2(n_496),
.B1(n_612),
.B2(n_460),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_662),
.A2(n_460),
.B(n_714),
.C(n_648),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_638),
.B(n_492),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_625),
.A2(n_460),
.B(n_714),
.C(n_632),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_707),
.A2(n_603),
.B1(n_623),
.B2(n_618),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_599),
.B(n_476),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_599),
.B(n_476),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_694),
.A2(n_702),
.B(n_698),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_602),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_654),
.B(n_464),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_654),
.B(n_464),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_603),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_661),
.B(n_496),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_603),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_597),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_654),
.Y(n_890)
);

OA21x2_ASAP7_75t_L g891 ( 
.A1(n_678),
.A2(n_479),
.B(n_477),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_694),
.A2(n_702),
.B(n_698),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_617),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_652),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_858),
.A2(n_876),
.B(n_878),
.C(n_747),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_806),
.B(n_827),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_808),
.B(n_864),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_SL g898 ( 
.A(n_865),
.B(n_875),
.C(n_873),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_785),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_841),
.Y(n_900)
);

NAND2x1_ASAP7_75t_SL g901 ( 
.A(n_746),
.B(n_868),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_801),
.B(n_849),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_769),
.Y(n_903)
);

AND2x6_ASAP7_75t_SL g904 ( 
.A(n_819),
.B(n_823),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_871),
.B(n_877),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_773),
.Y(n_906)
);

AO31x2_ASAP7_75t_L g907 ( 
.A1(n_742),
.A2(n_842),
.A3(n_882),
.B(n_892),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_L g908 ( 
.A1(n_816),
.A2(n_758),
.B(n_857),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_753),
.A2(n_890),
.B(n_857),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_890),
.B(n_860),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_748),
.B(n_795),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_870),
.B(n_869),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_856),
.A2(n_802),
.B(n_824),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_855),
.A2(n_839),
.B(n_861),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_872),
.A2(n_885),
.B(n_884),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_752),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_743),
.B(n_879),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_751),
.A2(n_757),
.B(n_738),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_767),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_806),
.B(n_790),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_814),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_757),
.A2(n_763),
.B(n_762),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_790),
.B(n_748),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_821),
.A2(n_856),
.B(n_793),
.C(n_810),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_859),
.Y(n_926)
);

AOI21xp33_ASAP7_75t_L g927 ( 
.A1(n_836),
.A2(n_764),
.B(n_826),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_879),
.B(n_809),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_867),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_880),
.B(n_881),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_863),
.A2(n_818),
.B1(n_809),
.B2(n_837),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_780),
.A2(n_765),
.B(n_750),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_883),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_881),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_849),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_842),
.A2(n_807),
.B(n_853),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_854),
.A2(n_891),
.B(n_789),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_813),
.B(n_886),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_803),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_838),
.A2(n_755),
.B(n_756),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_786),
.A2(n_754),
.B(n_846),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_888),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_744),
.B(n_817),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_833),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_766),
.A2(n_768),
.B(n_777),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_798),
.B(n_887),
.Y(n_946)
);

INVx6_ASAP7_75t_L g947 ( 
.A(n_769),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_817),
.B(n_812),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_827),
.B(n_798),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_891),
.A2(n_775),
.B(n_848),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_812),
.B(n_745),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_783),
.B(n_805),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_812),
.A2(n_828),
.B1(n_804),
.B2(n_820),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_774),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_801),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_812),
.B(n_844),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

OAI22x1_ASAP7_75t_L g958 ( 
.A1(n_829),
.A2(n_850),
.B1(n_825),
.B2(n_852),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_851),
.B(n_835),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_799),
.A2(n_800),
.B(n_797),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_L g961 ( 
.A(n_831),
.B(n_749),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_811),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_822),
.A2(n_792),
.B(n_782),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_827),
.B(n_759),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_847),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_834),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_894),
.B(n_893),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_840),
.A2(n_894),
.B(n_794),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_831),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_770),
.A2(n_739),
.B(n_832),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_SL g971 ( 
.A1(n_760),
.A2(n_776),
.B(n_845),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_792),
.A2(n_831),
.B1(n_843),
.B2(n_779),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_831),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_772),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_781),
.A2(n_778),
.B(n_791),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_830),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_772),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_791),
.A2(n_796),
.B(n_843),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_778),
.A2(n_889),
.B(n_779),
.C(n_815),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_889),
.A2(n_741),
.B(n_740),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_808),
.B(n_864),
.Y(n_981)
);

BUFx4_ASAP7_75t_SL g982 ( 
.A(n_883),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_801),
.B(n_849),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_849),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_857),
.B(n_890),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_857),
.B(n_890),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_857),
.B(n_890),
.Y(n_987)
);

BUFx10_ASAP7_75t_L g988 ( 
.A(n_883),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_857),
.B(n_890),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_858),
.A2(n_876),
.B1(n_865),
.B2(n_875),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_856),
.A2(n_802),
.B(n_824),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_767),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_857),
.B(n_890),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_806),
.B(n_827),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_740),
.A2(n_741),
.B(n_874),
.Y(n_995)
);

AOI21x1_ASAP7_75t_SL g996 ( 
.A1(n_837),
.A2(n_787),
.B(n_784),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_823),
.B(n_496),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_856),
.A2(n_802),
.B(n_824),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_823),
.A2(n_503),
.B1(n_460),
.B2(n_496),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_746),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_856),
.A2(n_802),
.B(n_824),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_856),
.A2(n_802),
.B(n_824),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_857),
.B(n_890),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_806),
.B(n_827),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_823),
.A2(n_858),
.B(n_876),
.C(n_878),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_823),
.A2(n_858),
.B(n_876),
.C(n_878),
.Y(n_1006)
);

AO21x2_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_742),
.B(n_761),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_773),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_857),
.B(n_890),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_806),
.B(n_827),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_870),
.B(n_503),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_862),
.B(n_541),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_740),
.A2(n_741),
.B(n_874),
.Y(n_1013)
);

AO31x2_ASAP7_75t_L g1014 ( 
.A1(n_742),
.A2(n_842),
.A3(n_866),
.B(n_861),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_857),
.B(n_890),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_808),
.B(n_864),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_808),
.B(n_864),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_858),
.A2(n_876),
.B(n_753),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_785),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_764),
.A2(n_496),
.B1(n_612),
.B2(n_600),
.Y(n_1020)
);

AO31x2_ASAP7_75t_L g1021 ( 
.A1(n_742),
.A2(n_842),
.A3(n_866),
.B(n_861),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_857),
.B(n_890),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_969),
.B(n_973),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_969),
.B(n_896),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_913),
.A2(n_998),
.B(n_991),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_999),
.A2(n_1006),
.B(n_1005),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_896),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_966),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_992),
.B(n_933),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_985),
.B(n_986),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_994),
.B(n_1004),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_990),
.A2(n_895),
.B(n_925),
.Y(n_1032)
);

CKINVDCx11_ASAP7_75t_R g1033 ( 
.A(n_939),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_911),
.B(n_905),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_1008),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_920),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_906),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_928),
.A2(n_1022),
.B1(n_985),
.B2(n_1015),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_913),
.A2(n_998),
.B(n_991),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_897),
.B(n_981),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_928),
.A2(n_1022),
.B1(n_986),
.B2(n_1015),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_SL g1042 ( 
.A1(n_1020),
.A2(n_904),
.B1(n_993),
.B2(n_1009),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_1010),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_901),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_987),
.B(n_989),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_900),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1016),
.B(n_1017),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_919),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_1000),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_895),
.A2(n_997),
.B(n_1018),
.C(n_898),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_1010),
.Y(n_1051)
);

BUFx10_ASAP7_75t_L g1052 ( 
.A(n_900),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_SL g1053 ( 
.A(n_1011),
.B(n_898),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_918),
.A2(n_963),
.B(n_937),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1000),
.B(n_987),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_989),
.A2(n_1009),
.B(n_993),
.C(n_1003),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_908),
.A2(n_927),
.B(n_1020),
.C(n_910),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_916),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_918),
.A2(n_963),
.B(n_1003),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_934),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_921),
.B(n_930),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_964),
.B(n_962),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_912),
.B(n_933),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_910),
.B(n_909),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_924),
.B(n_953),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_931),
.A2(n_927),
.B(n_923),
.C(n_936),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_992),
.B(n_949),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_982),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_922),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_902),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_938),
.A2(n_915),
.B1(n_929),
.B2(n_1019),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_964),
.A2(n_949),
.B1(n_1012),
.B2(n_946),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_975),
.A2(n_961),
.B(n_932),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_926),
.B(n_942),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_944),
.B(n_935),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_959),
.B(n_938),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_954),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_988),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_975),
.A2(n_956),
.B(n_971),
.C(n_951),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_935),
.B(n_984),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_900),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_982),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_951),
.A2(n_948),
.B1(n_943),
.B2(n_959),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_943),
.A2(n_979),
.B1(n_948),
.B2(n_972),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_955),
.B(n_977),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_945),
.B(n_976),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_903),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_965),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_903),
.Y(n_1089)
);

CKINVDCx11_ASAP7_75t_R g1090 ( 
.A(n_957),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1007),
.A2(n_914),
.B(n_940),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_947),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_967),
.B(n_977),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_941),
.A2(n_950),
.B(n_952),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_970),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_947),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_957),
.Y(n_1097)
);

OR2x2_ASAP7_75t_SL g1098 ( 
.A(n_947),
.B(n_957),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_958),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_983),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_955),
.B(n_907),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_907),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_978),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_SL g1105 ( 
.A1(n_960),
.A2(n_968),
.B1(n_980),
.B2(n_995),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_907),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1013),
.A2(n_996),
.B(n_1014),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1014),
.B(n_1021),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_1021),
.B(n_969),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1021),
.B(n_999),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1021),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_899),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_913),
.A2(n_856),
.B(n_991),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_899),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_896),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_939),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_917),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1020),
.A2(n_496),
.B1(n_314),
.B2(n_318),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_928),
.A2(n_999),
.B1(n_876),
.B2(n_858),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_913),
.A2(n_856),
.B(n_991),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_985),
.B(n_986),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1005),
.B(n_876),
.C(n_858),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_896),
.B(n_994),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_913),
.A2(n_856),
.B(n_991),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_911),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_906),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_906),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_982),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_917),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_899),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_985),
.B(n_986),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_969),
.B(n_973),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_966),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_911),
.B(n_748),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_896),
.B(n_994),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_982),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_969),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_985),
.B(n_986),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_969),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_899),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_911),
.B(n_748),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_982),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_982),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_897),
.B(n_981),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_985),
.B(n_986),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_969),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_982),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1139),
.B(n_1146),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1034),
.B(n_1125),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1053),
.A2(n_1032),
.B1(n_1119),
.B2(n_1122),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1074),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1032),
.A2(n_1122),
.B(n_1026),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1139),
.B(n_1146),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_SL g1154 ( 
.A1(n_1053),
.A2(n_1042),
.B1(n_1111),
.B2(n_1110),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1042),
.A2(n_1118),
.B1(n_1026),
.B2(n_1119),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1038),
.A2(n_1041),
.B1(n_1131),
.B2(n_1121),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1058),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1037),
.Y(n_1159)
);

BUFx8_ASAP7_75t_L g1160 ( 
.A(n_1028),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1102),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1069),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1112),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1035),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1114),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1130),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1103),
.Y(n_1168)
);

OAI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1038),
.A2(n_1041),
.B1(n_1121),
.B2(n_1030),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1140),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1045),
.B(n_1131),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1134),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1141),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1050),
.A2(n_1066),
.B(n_1073),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1077),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1025),
.A2(n_1039),
.B(n_1048),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1126),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1057),
.A2(n_1056),
.B(n_1059),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1045),
.B(n_1145),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1145),
.B(n_1055),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1144),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1065),
.A2(n_1061),
.B1(n_1072),
.B2(n_1044),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1071),
.A2(n_1064),
.B(n_1084),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1100),
.A2(n_1044),
.B1(n_1084),
.B2(n_1125),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1090),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1068),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1064),
.A2(n_1071),
.B1(n_1063),
.B2(n_1106),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1052),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1052),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1075),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1098),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1091),
.A2(n_1107),
.B(n_1094),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1036),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1108),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1083),
.A2(n_1060),
.B1(n_1076),
.B2(n_1117),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1088),
.B(n_1127),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1102),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1076),
.A2(n_1129),
.B1(n_1062),
.B2(n_1086),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1049),
.A2(n_1072),
.B1(n_1079),
.B2(n_1067),
.Y(n_1199)
);

BUFx2_ASAP7_75t_R g1200 ( 
.A(n_1142),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1113),
.A2(n_1120),
.B(n_1124),
.C(n_1054),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1029),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1093),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1089),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1109),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1082),
.A2(n_1128),
.B(n_1136),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1087),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1062),
.A2(n_1123),
.B1(n_1135),
.B2(n_1031),
.Y(n_1208)
);

CKINVDCx11_ASAP7_75t_R g1209 ( 
.A(n_1116),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1031),
.A2(n_1135),
.B1(n_1123),
.B2(n_1027),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1099),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1027),
.A2(n_1051),
.B1(n_1115),
.B2(n_1043),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1027),
.B(n_1115),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1109),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1104),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1097),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1024),
.A2(n_1115),
.B1(n_1043),
.B2(n_1051),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1097),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1092),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1137),
.B(n_1070),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1143),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1080),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1043),
.B(n_1051),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1101),
.B(n_1096),
.Y(n_1225)
);

AO21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1105),
.A2(n_1023),
.B(n_1132),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1046),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1085),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1081),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1081),
.A2(n_1078),
.B1(n_1133),
.B2(n_1033),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1081),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1147),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1102),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1095),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1037),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1040),
.B(n_1144),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1134),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1116),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1068),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1102),
.Y(n_1241)
);

BUFx2_ASAP7_75t_R g1242 ( 
.A(n_1068),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1025),
.A2(n_1039),
.B(n_1048),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1053),
.A2(n_999),
.B1(n_865),
.B2(n_875),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1052),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1040),
.B(n_1144),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1053),
.A2(n_496),
.B1(n_1042),
.B2(n_314),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1074),
.Y(n_1248)
);

AO21x1_ASAP7_75t_SL g1249 ( 
.A1(n_1032),
.A2(n_1026),
.B(n_928),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1052),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1215),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1219),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1219),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1162),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1194),
.B(n_1249),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1178),
.A2(n_1174),
.B(n_1201),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1162),
.B(n_1197),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1205),
.B(n_1214),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1197),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1209),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1183),
.A2(n_1201),
.A3(n_1168),
.B(n_1235),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1233),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1241),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1241),
.B(n_1176),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1176),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1169),
.B(n_1176),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1243),
.B(n_1152),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1169),
.B(n_1156),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1243),
.B(n_1180),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1156),
.B(n_1151),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1203),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1150),
.B(n_1190),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1192),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1177),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1158),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1196),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1163),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1164),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1175),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1166),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1248),
.B(n_1167),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1244),
.A2(n_1150),
.B(n_1170),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1226),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1149),
.B(n_1171),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1198),
.A2(n_1195),
.B(n_1155),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1207),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1179),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_1157),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1237),
.B(n_1246),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1198),
.A2(n_1155),
.B(n_1234),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1161),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1199),
.A2(n_1148),
.B(n_1153),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1161),
.B(n_1181),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1159),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1223),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1236),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1154),
.B(n_1228),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1244),
.A2(n_1182),
.B(n_1217),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1216),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1184),
.B(n_1247),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1218),
.B(n_1231),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1239),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1211),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1172),
.A2(n_1238),
.B1(n_1173),
.B2(n_1208),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1165),
.B(n_1229),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1221),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1225),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1269),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1287),
.B(n_1220),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1267),
.B(n_1232),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1267),
.B(n_1232),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1254),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1283),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1267),
.B(n_1193),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1269),
.B(n_1220),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1268),
.A2(n_1148),
.B(n_1153),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1279),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1265),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1264),
.B(n_1185),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1287),
.B(n_1227),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1265),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1264),
.B(n_1230),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1268),
.B(n_1206),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1264),
.B(n_1230),
.Y(n_1324)
);

INVx3_ASAP7_75t_SL g1325 ( 
.A(n_1283),
.Y(n_1325)
);

INVxp33_ASAP7_75t_L g1326 ( 
.A(n_1293),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1266),
.B(n_1213),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1269),
.B(n_1227),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1300),
.A2(n_1208),
.B1(n_1191),
.B2(n_1210),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1283),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1291),
.B(n_1204),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1305),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1255),
.B(n_1204),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1291),
.B(n_1250),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1257),
.B(n_1224),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_L g1336 ( 
.A(n_1256),
.B(n_1202),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1283),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1261),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1256),
.B(n_1245),
.Y(n_1339)
);

INVxp67_ASAP7_75t_SL g1340 ( 
.A(n_1254),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1259),
.Y(n_1341)
);

INVx4_ASAP7_75t_L g1342 ( 
.A(n_1283),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1261),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1261),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1259),
.B(n_1188),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1257),
.B(n_1189),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1261),
.B(n_1210),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1261),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1261),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1261),
.B(n_1212),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1277),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1277),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1322),
.B(n_1252),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1323),
.B(n_1303),
.C(n_1286),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1323),
.B(n_1303),
.C(n_1286),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1316),
.B(n_1283),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1338),
.A2(n_1300),
.B1(n_1288),
.B2(n_1270),
.C(n_1271),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1347),
.A2(n_1298),
.B1(n_1285),
.B2(n_1290),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1319),
.B(n_1276),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1319),
.B(n_1276),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1319),
.B(n_1296),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1339),
.B(n_1262),
.C(n_1263),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1322),
.B(n_1253),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1338),
.A2(n_1288),
.B1(n_1270),
.B2(n_1271),
.C(n_1278),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1322),
.B(n_1253),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1317),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1324),
.B(n_1253),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1347),
.A2(n_1285),
.B1(n_1298),
.B2(n_1290),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1324),
.B(n_1270),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1339),
.B(n_1296),
.C(n_1299),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1324),
.B(n_1289),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1314),
.B(n_1289),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_1274),
.Y(n_1373)
);

OAI221xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1338),
.A2(n_1288),
.B1(n_1272),
.B2(n_1304),
.C(n_1297),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1310),
.B(n_1274),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1310),
.B(n_1307),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1339),
.B(n_1263),
.C(n_1275),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1336),
.B(n_1299),
.C(n_1275),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1311),
.B(n_1294),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1311),
.B(n_1294),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1329),
.A2(n_1298),
.B1(n_1285),
.B2(n_1282),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1314),
.B(n_1289),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1309),
.B(n_1293),
.Y(n_1384)
);

AND2x2_ASAP7_75t_SL g1385 ( 
.A(n_1347),
.B(n_1285),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1309),
.B(n_1293),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1320),
.B(n_1281),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1314),
.B(n_1251),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1331),
.B(n_1273),
.C(n_1272),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1329),
.A2(n_1298),
.B1(n_1285),
.B2(n_1290),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1320),
.B(n_1308),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1327),
.B(n_1251),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1308),
.B(n_1281),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1331),
.B(n_1273),
.C(n_1272),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1336),
.B(n_1301),
.C(n_1295),
.Y(n_1395)
);

AND2x2_ASAP7_75t_SL g1396 ( 
.A(n_1350),
.B(n_1258),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_L g1397 ( 
.A(n_1345),
.B(n_1305),
.C(n_1306),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1327),
.B(n_1251),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1316),
.A2(n_1282),
.B(n_1292),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1308),
.B(n_1281),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1317),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1327),
.B(n_1251),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1334),
.B(n_1282),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1384),
.B(n_1260),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1403),
.B(n_1334),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1371),
.B(n_1312),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1395),
.B(n_1330),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1366),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1371),
.B(n_1312),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1401),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1401),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1385),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1395),
.B(n_1330),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1385),
.A2(n_1282),
.B1(n_1350),
.B2(n_1290),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1354),
.B(n_1340),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1372),
.B(n_1332),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1396),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1391),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1396),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1354),
.B(n_1340),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1372),
.B(n_1383),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1385),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1353),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1393),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1400),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1392),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1382),
.A2(n_1350),
.B1(n_1290),
.B2(n_1297),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1396),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1376),
.B(n_1335),
.Y(n_1432)
);

XOR2xp5_ASAP7_75t_L g1433 ( 
.A(n_1382),
.B(n_1239),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1383),
.B(n_1332),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1353),
.B(n_1326),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1362),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1355),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1379),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1355),
.B(n_1341),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1363),
.B(n_1326),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1363),
.B(n_1333),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1370),
.B(n_1341),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1365),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1380),
.B(n_1315),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1387),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1365),
.B(n_1367),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1367),
.B(n_1330),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1418),
.B(n_1392),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1418),
.B(n_1378),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1408),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1436),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1419),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1405),
.B(n_1419),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1418),
.B(n_1402),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1418),
.B(n_1378),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1438),
.B(n_1397),
.Y(n_1457)
);

NAND2x1p5_ASAP7_75t_L g1458 ( 
.A(n_1421),
.B(n_1356),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1421),
.B(n_1398),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1436),
.B(n_1386),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1404),
.B(n_1209),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1421),
.B(n_1313),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1433),
.B(n_1160),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_1402),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1433),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1437),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1429),
.B(n_1381),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1408),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1409),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1431),
.B(n_1398),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1437),
.B(n_1420),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1429),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1431),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1420),
.B(n_1359),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1431),
.B(n_1388),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1423),
.B(n_1388),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1443),
.A2(n_1368),
.B(n_1374),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1423),
.B(n_1360),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1430),
.A2(n_1357),
.B1(n_1390),
.B2(n_1364),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1415),
.A2(n_1424),
.B1(n_1413),
.B2(n_1358),
.C(n_1399),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1411),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1448),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1447),
.B(n_1373),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1411),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1432),
.B(n_1361),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1451),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1452),
.B(n_1416),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.B(n_1472),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1467),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1477),
.B(n_1447),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1453),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1453),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1450),
.B(n_1407),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1484),
.B(n_1442),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1451),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1422),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1469),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1469),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1484),
.B(n_1407),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1474),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1464),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1470),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1407),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1461),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1466),
.B(n_1302),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_L g1512 ( 
.A(n_1450),
.B(n_1407),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1480),
.A2(n_1424),
.B1(n_1413),
.B2(n_1443),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1460),
.B(n_1479),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1470),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1474),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1480),
.A2(n_1424),
.B1(n_1413),
.B2(n_1394),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_L g1518 ( 
.A(n_1456),
.B(n_1414),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1482),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1479),
.B(n_1439),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1439),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1478),
.B(n_1446),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1487),
.B(n_1446),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1482),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1483),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1481),
.A2(n_1348),
.B1(n_1349),
.B2(n_1344),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1456),
.B(n_1414),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1486),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1456),
.B(n_1414),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1456),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1521),
.B(n_1463),
.C(n_1483),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1522),
.A2(n_1349),
.B1(n_1338),
.B2(n_1348),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1507),
.B(n_1468),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1490),
.B(n_1485),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1528),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1510),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1488),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_1511),
.Y(n_1540)
);

AOI222xp33_ASAP7_75t_L g1541 ( 
.A1(n_1513),
.A2(n_1463),
.B1(n_1344),
.B2(n_1348),
.C1(n_1349),
.C2(n_1343),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1511),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.B(n_1449),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1506),
.B(n_1186),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1490),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1527),
.A2(n_1344),
.B1(n_1348),
.B2(n_1349),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1499),
.B(n_1475),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1502),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1512),
.B(n_1449),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1491),
.B(n_1463),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1503),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1463),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1468),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1523),
.B(n_1525),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.B(n_1486),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1508),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1489),
.B(n_1345),
.C(n_1414),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1516),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1519),
.Y(n_1565)
);

CKINVDCx16_ASAP7_75t_R g1566 ( 
.A(n_1528),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1532),
.A2(n_1517),
.B(n_1495),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1540),
.A2(n_1518),
.B1(n_1500),
.B2(n_1493),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

NAND2x1_ASAP7_75t_L g1570 ( 
.A(n_1537),
.B(n_1528),
.Y(n_1570)
);

OAI32xp33_ASAP7_75t_L g1571 ( 
.A1(n_1566),
.A2(n_1495),
.A3(n_1530),
.B1(n_1458),
.B2(n_1504),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1555),
.Y(n_1572)
);

AOI32xp33_ASAP7_75t_L g1573 ( 
.A1(n_1550),
.A2(n_1530),
.A3(n_1509),
.B1(n_1504),
.B2(n_1493),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1547),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1537),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1563),
.A2(n_1495),
.B(n_1505),
.C(n_1458),
.Y(n_1579)
);

OAI31xp33_ASAP7_75t_L g1580 ( 
.A1(n_1562),
.A2(n_1509),
.A3(n_1494),
.B(n_1500),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_SL g1581 ( 
.A1(n_1544),
.A2(n_1505),
.B(n_1160),
.C(n_1524),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1559),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1494),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1537),
.B(n_1459),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1536),
.B(n_1526),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1535),
.A2(n_1458),
.B1(n_1462),
.B2(n_1459),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1531),
.B(n_1529),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1556),
.A2(n_1553),
.B(n_1552),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1531),
.B(n_1465),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1559),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1543),
.B(n_1465),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1592),
.B(n_1533),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1577),
.B(n_1549),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1574),
.B(n_1558),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1558),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1569),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1583),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1587),
.B(n_1543),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1576),
.B(n_1552),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_L g1607 ( 
.A(n_1573),
.B(n_1186),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1591),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1591),
.B(n_1557),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1557),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1589),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1589),
.B(n_1539),
.Y(n_1612)
);

AOI222xp33_ASAP7_75t_L g1613 ( 
.A1(n_1599),
.A2(n_1534),
.B1(n_1548),
.B2(n_1571),
.C1(n_1564),
.C2(n_1561),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1603),
.A2(n_1567),
.B1(n_1580),
.B2(n_1579),
.C(n_1568),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1603),
.A2(n_1579),
.B1(n_1581),
.B2(n_1546),
.C(n_1551),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1606),
.A2(n_1581),
.B1(n_1565),
.B2(n_1586),
.C(n_1570),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1595),
.A2(n_1560),
.B1(n_1589),
.B2(n_1541),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1594),
.B(n_1584),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1608),
.A2(n_1560),
.B1(n_1462),
.B2(n_1344),
.Y(n_1619)
);

OAI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1596),
.A2(n_1462),
.B(n_1476),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1602),
.A2(n_1471),
.B1(n_1476),
.B2(n_1412),
.C(n_1426),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1597),
.B(n_1471),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1611),
.A2(n_1412),
.B(n_1448),
.C(n_1427),
.Y(n_1623)
);

OAI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1607),
.A2(n_1343),
.B1(n_1304),
.B2(n_1315),
.C(n_1328),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1617),
.A2(n_1612),
.B(n_1605),
.C(n_1601),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1615),
.A2(n_1598),
.B(n_1604),
.C(n_1600),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1618),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1622),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1623),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1614),
.B(n_1613),
.C(n_1616),
.Y(n_1630)
);

OAI21xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1624),
.A2(n_1609),
.B(n_1610),
.Y(n_1631)
);

NOR3xp33_ASAP7_75t_L g1632 ( 
.A(n_1619),
.B(n_1593),
.C(n_1240),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1621),
.B(n_1222),
.Y(n_1633)
);

NOR4xp25_ASAP7_75t_L g1634 ( 
.A(n_1620),
.B(n_1160),
.C(n_1406),
.D(n_1410),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1614),
.A2(n_1200),
.B(n_1242),
.C(n_1240),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1627),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_SL g1637 ( 
.A1(n_1625),
.A2(n_1222),
.B(n_1318),
.C(n_1321),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1629),
.A2(n_1428),
.B(n_1417),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1630),
.B(n_1448),
.Y(n_1639)
);

NAND4xp25_ASAP7_75t_L g1640 ( 
.A(n_1635),
.B(n_1626),
.C(n_1628),
.D(n_1633),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1427),
.Y(n_1641)
);

NOR2x2_ASAP7_75t_L g1642 ( 
.A(n_1640),
.B(n_1635),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1636),
.B(n_1634),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1641),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1638),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1637),
.A2(n_1632),
.B1(n_1448),
.B2(n_1435),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1636),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1647),
.B(n_1305),
.Y(n_1648)
);

OR3x1_ASAP7_75t_L g1649 ( 
.A(n_1644),
.B(n_1352),
.C(n_1351),
.Y(n_1649)
);

NOR4xp75_ASAP7_75t_L g1650 ( 
.A(n_1645),
.B(n_1375),
.C(n_1428),
.D(n_1417),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1643),
.B(n_1284),
.C(n_1315),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1434),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_L g1653 ( 
.A(n_1652),
.B(n_1651),
.Y(n_1653)
);

AOI31xp33_ASAP7_75t_L g1654 ( 
.A1(n_1648),
.A2(n_1646),
.A3(n_1346),
.B(n_1434),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1650),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1653),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1655),
.B(n_1654),
.C(n_1649),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1657),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_SL g1659 ( 
.A1(n_1657),
.A2(n_1342),
.B(n_1313),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1444),
.B(n_1425),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1441),
.B(n_1435),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1660),
.B(n_1445),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1661),
.A2(n_1444),
.B(n_1425),
.Y(n_1663)
);

XOR2xp5_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1284),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1663),
.B1(n_1280),
.B2(n_1278),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_R g1666 ( 
.A1(n_1665),
.A2(n_1325),
.B1(n_1313),
.B2(n_1342),
.C(n_1444),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1325),
.B(n_1337),
.C(n_1330),
.Y(n_1667)
);


endmodule