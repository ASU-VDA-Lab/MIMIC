module fake_jpeg_14144_n_519 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_52),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_54),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_8),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_8),
.C(n_1),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_87),
.B(n_38),
.C(n_42),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_73),
.Y(n_114)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_69),
.Y(n_147)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_8),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_82),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_0),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_29),
.B(n_45),
.Y(n_151)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_1),
.C(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_89),
.B(n_27),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_R g96 ( 
.A(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_43),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_40),
.Y(n_136)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_101),
.A2(n_106),
.B1(n_121),
.B2(n_122),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_50),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_43),
.B1(n_47),
.B2(n_27),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_64),
.A2(n_73),
.B1(n_59),
.B2(n_87),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_48),
.B1(n_32),
.B2(n_40),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_18),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_126),
.B(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_40),
.B1(n_48),
.B2(n_32),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_135),
.B1(n_137),
.B2(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_132),
.B(n_145),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_79),
.B1(n_68),
.B2(n_63),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_33),
.B1(n_44),
.B2(n_36),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_32),
.B1(n_49),
.B2(n_33),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_36),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_70),
.B1(n_49),
.B2(n_93),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_55),
.B1(n_84),
.B2(n_81),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_46),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_46),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_154),
.B(n_157),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_62),
.A2(n_45),
.B1(n_42),
.B2(n_38),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_56),
.B1(n_65),
.B2(n_52),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_79),
.B(n_91),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_161),
.B(n_189),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_72),
.A3(n_76),
.B1(n_67),
.B2(n_58),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_180),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_98),
.C(n_85),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_191),
.C(n_198),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_168),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_1),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_203),
.Y(n_222)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_171),
.Y(n_250)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_107),
.B(n_75),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_179),
.B(n_190),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_110),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_183),
.B1(n_205),
.B2(n_209),
.Y(n_224)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_92),
.B1(n_90),
.B2(n_71),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_185),
.B(n_186),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_108),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_74),
.B(n_3),
.C(n_4),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_122),
.B(n_15),
.C(n_17),
.Y(n_220)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_129),
.A2(n_118),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_111),
.B(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_5),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_101),
.B(n_5),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_210),
.C(n_198),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_200),
.B(n_204),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_141),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_179),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_128),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_6),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_116),
.B(n_7),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_138),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_217),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_123),
.B(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_212),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_140),
.B(n_17),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_12),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_210),
.Y(n_264)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

BUFx24_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_139),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_139),
.B1(n_124),
.B2(n_149),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_113),
.B1(n_109),
.B2(n_142),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_218),
.A2(n_234),
.B1(n_237),
.B2(n_254),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_238),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_227),
.A2(n_170),
.B1(n_171),
.B2(n_196),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_163),
.A2(n_142),
.B1(n_113),
.B2(n_159),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_233),
.A2(n_236),
.B1(n_244),
.B2(n_257),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_143),
.B1(n_158),
.B2(n_115),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_161),
.A2(n_158),
.B1(n_103),
.B2(n_120),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_169),
.A2(n_125),
.B1(n_120),
.B2(n_103),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_125),
.B1(n_115),
.B2(n_152),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_215),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_176),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_162),
.A2(n_13),
.B1(n_119),
.B2(n_180),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_193),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_164),
.A2(n_13),
.B1(n_211),
.B2(n_197),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_191),
.A2(n_198),
.B(n_184),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_259),
.B(n_242),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_208),
.A2(n_191),
.B1(n_213),
.B2(n_210),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_212),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_185),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_207),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_167),
.B(n_173),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_270),
.B(n_271),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_286),
.B1(n_313),
.B2(n_232),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_160),
.B1(n_174),
.B2(n_192),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_274),
.A2(n_302),
.B1(n_305),
.B2(n_225),
.Y(n_340)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_294),
.C(n_252),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_222),
.B(n_194),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_278),
.B(n_280),
.Y(n_331)
);

BUFx24_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_245),
.B(n_186),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_287),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_283),
.B(n_285),
.Y(n_354)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_248),
.B(n_177),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_228),
.A2(n_160),
.B1(n_195),
.B2(n_188),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_172),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_215),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_249),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_217),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_165),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_176),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_226),
.B(n_182),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_303),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_SL g347 ( 
.A(n_301),
.B(n_256),
.C(n_258),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_240),
.A2(n_175),
.B1(n_200),
.B2(n_178),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_176),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_223),
.A2(n_214),
.B(n_193),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_223),
.B(n_250),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_240),
.A2(n_193),
.B1(n_237),
.B2(n_252),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_307),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_222),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_311),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_257),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_244),
.B(n_229),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_320),
.A2(n_342),
.B(n_268),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_255),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_326),
.C(n_332),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_281),
.B(n_301),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_328),
.A2(n_339),
.B(n_295),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_292),
.A2(n_252),
.B1(n_220),
.B2(n_233),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_337),
.B1(n_350),
.B2(n_268),
.Y(n_365)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_275),
.A2(n_246),
.A3(n_224),
.B1(n_251),
.B2(n_256),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_347),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_292),
.A2(n_224),
.B1(n_231),
.B2(n_227),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_281),
.A2(n_250),
.B(n_229),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_346),
.B1(n_312),
.B2(n_289),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_281),
.B(n_274),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_269),
.A2(n_231),
.B1(n_262),
.B2(n_251),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_286),
.A2(n_219),
.B1(n_261),
.B2(n_258),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_239),
.C(n_225),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_307),
.C(n_288),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_271),
.Y(n_357)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_331),
.B(n_278),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_358),
.B(n_372),
.Y(n_406)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

XOR2x2_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_325),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_360),
.B(n_388),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_368),
.Y(n_400)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_365),
.A2(n_375),
.B1(n_347),
.B2(n_317),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_302),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_300),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_318),
.A3(n_354),
.B1(n_315),
.B2(n_328),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_369),
.A2(n_330),
.B1(n_343),
.B2(n_345),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_331),
.B(n_287),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_310),
.B(n_303),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_333),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_376),
.Y(n_411)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_337),
.A2(n_283),
.B1(n_309),
.B2(n_272),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_282),
.B(n_279),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_321),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_377),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_382),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_320),
.B1(n_318),
.B2(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_284),
.B(n_298),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_347),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_321),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_311),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_353),
.C(n_349),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_346),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_306),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_341),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_299),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_355),
.B(n_325),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_402),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_397),
.A2(n_356),
.B1(n_365),
.B2(n_385),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_332),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_399),
.C(n_403),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_355),
.B(n_360),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_338),
.C(n_354),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_372),
.C(n_362),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_410),
.C(n_415),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_371),
.B(n_323),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_416),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_349),
.C(n_351),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_413),
.A2(n_369),
.B1(n_361),
.B2(n_383),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_329),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_357),
.B(n_344),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_344),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_418),
.C(n_416),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_351),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_420),
.A2(n_437),
.B1(n_414),
.B2(n_397),
.Y(n_444)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_373),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_418),
.B(n_382),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_377),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_404),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_428),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_434),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_361),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_440),
.C(n_442),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_387),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_431),
.B(n_435),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_367),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_436),
.B(n_439),
.Y(n_463)
);

OAI21xp33_ASAP7_75t_SL g437 ( 
.A1(n_392),
.A2(n_370),
.B(n_376),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_438),
.A2(n_378),
.B1(n_405),
.B2(n_417),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_406),
.B(n_358),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_381),
.C(n_375),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_411),
.A2(n_356),
.B(n_366),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_441),
.A2(n_366),
.B(n_388),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

BUFx12_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_444),
.A2(n_450),
.B1(n_462),
.B2(n_445),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_413),
.B1(n_363),
.B2(n_391),
.Y(n_447)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_443),
.A2(n_401),
.B1(n_396),
.B2(n_408),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_449),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_420),
.A2(n_415),
.B1(n_366),
.B2(n_392),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_451),
.A2(n_352),
.B(n_335),
.Y(n_479)
);

NOR4xp25_ASAP7_75t_L g452 ( 
.A(n_433),
.B(n_407),
.C(n_402),
.D(n_389),
.Y(n_452)
);

OAI221xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_425),
.B1(n_433),
.B2(n_427),
.C(n_423),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_389),
.B1(n_380),
.B2(n_374),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_458),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_398),
.C(n_348),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_422),
.B1(n_424),
.B2(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_460),
.B(n_427),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_465),
.A2(n_474),
.B1(n_461),
.B2(n_457),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_430),
.B(n_435),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_466),
.A2(n_467),
.B(n_468),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_432),
.B(n_442),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_444),
.A2(n_432),
.B(n_421),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_448),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_469),
.B(n_472),
.Y(n_482)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_419),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_446),
.A2(n_429),
.B(n_322),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_473),
.A2(n_479),
.B(n_462),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_450),
.A2(n_317),
.B1(n_359),
.B2(n_350),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_447),
.B1(n_455),
.B2(n_449),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_335),
.Y(n_477)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_477),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_425),
.C(n_348),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_461),
.C(n_453),
.Y(n_491)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_475),
.A2(n_454),
.B1(n_462),
.B2(n_453),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_484),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_456),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_489),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_487),
.B(n_490),
.Y(n_494)
);

A2O1A1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_457),
.B(n_461),
.C(n_452),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_466),
.A2(n_456),
.B(n_457),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_476),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_493),
.A2(n_479),
.B1(n_467),
.B2(n_457),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_464),
.C(n_470),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_496),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_470),
.C(n_478),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_299),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_481),
.Y(n_506)
);

AOI31xp67_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_279),
.A3(n_352),
.B(n_276),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_279),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_488),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_504),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_507),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_495),
.B(n_480),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_496),
.C(n_497),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_513),
.C(n_500),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_499),
.C(n_480),
.Y(n_513)
);

OAI311xp33_ASAP7_75t_L g514 ( 
.A1(n_510),
.A2(n_489),
.A3(n_493),
.B1(n_504),
.C1(n_508),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_515),
.C(n_511),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_484),
.C(n_494),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_517),
.B(n_219),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_518),
.B(n_261),
.Y(n_519)
);


endmodule