module fake_jpeg_15778_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_3),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g103 ( 
.A(n_39),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_56),
.Y(n_66)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_2),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_SL g55 ( 
.A(n_25),
.B(n_2),
.C(n_6),
.Y(n_55)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_19),
.B1(n_32),
.B2(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_27),
.B(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_34),
.B1(n_22),
.B2(n_30),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_79),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_81),
.C(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_28),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_83),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_35),
.Y(n_82)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_85),
.B(n_91),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_88),
.Y(n_114)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_35),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_29),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_94),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_32),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_21),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_29),
.B1(n_20),
.B2(n_24),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_24),
.B1(n_21),
.B2(n_19),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_107),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_20),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_133),
.B1(n_83),
.B2(n_36),
.Y(n_162)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_72),
.B1(n_10),
.B2(n_14),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_50),
.B1(n_10),
.B2(n_13),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_76),
.B1(n_72),
.B2(n_73),
.Y(n_136)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_77),
.A2(n_19),
.B(n_36),
.C(n_62),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_87),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_31),
.C(n_37),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_37),
.C(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_136),
.B(n_153),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_89),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_158),
.C(n_163),
.Y(n_168)
);

OR2x6_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_103),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_141),
.Y(n_186)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_132),
.B1(n_113),
.B2(n_110),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_130),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_71),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_160),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_8),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_103),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_133),
.A3(n_118),
.B1(n_114),
.B2(n_112),
.Y(n_176)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_164),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_88),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_86),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_98),
.C(n_102),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_108),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_118),
.B1(n_105),
.B2(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_178),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_163),
.C(n_148),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_181),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_115),
.B1(n_121),
.B2(n_104),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_137),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_141),
.B(n_162),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_141),
.B(n_186),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_158),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_183),
.C(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_140),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

AO221x1_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_172),
.B1(n_167),
.B2(n_177),
.C(n_170),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_208),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_173),
.C(n_151),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_192),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_141),
.C(n_149),
.Y(n_211)
);

OAI321xp33_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_159),
.A3(n_182),
.B1(n_188),
.B2(n_196),
.C(n_198),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_173),
.B(n_184),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_201),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_171),
.B1(n_147),
.B2(n_150),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_167),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_222),
.B1(n_209),
.B2(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_225),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_197),
.B1(n_189),
.B2(n_203),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_189),
.B1(n_208),
.B2(n_211),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_200),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_188),
.B(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_210),
.C(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_226),
.C(n_221),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_233),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_231),
.B(n_223),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_165),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_237),
.C(n_221),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_230),
.C(n_179),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_234),
.B(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_241),
.B(n_36),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_166),
.B(n_106),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);


endmodule