module fake_jpeg_198_n_130 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_9),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp67_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_5),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_37),
.C(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_6),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_46),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_13),
.B1(n_12),
.B2(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_11),
.B1(n_27),
.B2(n_21),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_20),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_11),
.B1(n_13),
.B2(n_26),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_12),
.B1(n_22),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_3),
.B1(n_24),
.B2(n_38),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_3),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_65),
.C(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_83),
.B1(n_69),
.B2(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_44),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_70),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_64),
.B1(n_56),
.B2(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_86),
.B1(n_69),
.B2(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_67),
.B1(n_60),
.B2(n_66),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_55),
.B(n_65),
.C(n_68),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

BUFx12f_ASAP7_75t_SL g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_73),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_99),
.Y(n_101)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_84),
.B1(n_88),
.B2(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_74),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_75),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_75),
.C(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_98),
.C(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_92),
.B(n_94),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_98),
.C(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_101),
.A3(n_92),
.B1(n_97),
.B2(n_104),
.C(n_105),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_121),
.B1(n_115),
.B2(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_101),
.C(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_104),
.B(n_97),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_76),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_76),
.B(n_126),
.C(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_88),
.B(n_90),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_90),
.Y(n_130)
);


endmodule