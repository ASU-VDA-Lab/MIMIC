module real_aes_15600_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_0), .A2(n_58), .B1(n_497), .B2(n_501), .C(n_507), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_0), .A2(n_58), .B1(n_581), .B2(n_587), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_1), .A2(n_31), .B1(n_117), .B2(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g493 ( .A(n_2), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_2), .A2(n_73), .B1(n_567), .B2(n_573), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_3), .A2(n_71), .B1(n_468), .B2(n_471), .C(n_475), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_3), .A2(n_19), .B1(n_43), .B2(n_603), .C1(n_606), .C2(n_608), .Y(n_602) );
AND2x2_ASAP7_75t_L g464 ( .A(n_4), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g478 ( .A(n_4), .Y(n_478) );
AND2x2_ASAP7_75t_L g488 ( .A(n_4), .B(n_66), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_5), .A2(n_10), .B1(n_111), .B2(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_6), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_7), .A2(n_11), .B1(n_86), .B2(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_9), .Y(n_168) );
INVxp67_ASAP7_75t_SL g520 ( .A(n_12), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_12), .A2(n_71), .B1(n_622), .B2(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g540 ( .A(n_13), .Y(n_540) );
INVx1_ASAP7_75t_L g560 ( .A(n_13), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_14), .A2(n_76), .B1(n_111), .B2(n_113), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_15), .A2(n_27), .B1(n_159), .B2(n_160), .Y(n_158) );
INVx2_ASAP7_75t_L g548 ( .A(n_16), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_17), .B(n_112), .Y(n_178) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_18), .A2(n_42), .B(n_126), .Y(n_125) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_19), .A2(n_48), .B1(n_480), .B2(n_486), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_20), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_21), .A2(n_35), .B1(n_134), .B2(n_137), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_22), .A2(n_40), .B1(n_111), .B2(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_23), .Y(n_213) );
INVx1_ASAP7_75t_L g626 ( .A(n_24), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_25), .B(n_159), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_26), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_28), .A2(n_65), .B1(n_117), .B2(n_207), .Y(n_206) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_29), .A2(n_457), .B(n_466), .C(n_489), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_29), .A2(n_59), .B1(n_535), .B2(n_554), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_30), .A2(n_33), .B1(n_117), .B2(n_149), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_32), .A2(n_44), .B1(n_111), .B2(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_34), .Y(n_513) );
XNOR2xp5_ASAP7_75t_L g453 ( .A(n_36), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_37), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g564 ( .A(n_37), .Y(n_564) );
INVx1_ASAP7_75t_L g615 ( .A(n_37), .Y(n_615) );
INVx2_ASAP7_75t_L g665 ( .A(n_38), .Y(n_665) );
BUFx2_ASAP7_75t_L g646 ( .A(n_39), .Y(n_646) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_40), .Y(n_675) );
INVx1_ASAP7_75t_L g651 ( .A(n_41), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_43), .A2(n_61), .B1(n_522), .B2(n_523), .C(n_524), .Y(n_521) );
BUFx3_ASAP7_75t_L g542 ( .A(n_45), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_46), .A2(n_55), .B1(n_116), .B2(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_47), .A2(n_57), .B1(n_117), .B2(n_149), .Y(n_189) );
INVx1_ASAP7_75t_L g620 ( .A(n_48), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_49), .A2(n_74), .B1(n_111), .B2(n_147), .Y(n_188) );
AND2x4_ASAP7_75t_L g95 ( .A(n_50), .B(n_96), .Y(n_95) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_50), .Y(n_639) );
INVx1_ASAP7_75t_L g126 ( .A(n_51), .Y(n_126) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_52), .Y(n_461) );
INVx1_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_54), .Y(n_463) );
INVx1_ASAP7_75t_L g654 ( .A(n_56), .Y(n_654) );
INVx2_ASAP7_75t_L g92 ( .A(n_60), .Y(n_92) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_61), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_62), .A2(n_75), .B1(n_137), .B2(n_210), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_62), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_62), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_63), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_64), .Y(n_231) );
INVx1_ASAP7_75t_L g465 ( .A(n_66), .Y(n_465) );
BUFx3_ASAP7_75t_L g477 ( .A(n_66), .Y(n_477) );
INVx2_ASAP7_75t_L g531 ( .A(n_67), .Y(n_531) );
INVx1_ASAP7_75t_L g546 ( .A(n_67), .Y(n_546) );
INVx1_ASAP7_75t_L g586 ( .A(n_67), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_68), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g647 ( .A(n_69), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_70), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_72), .B(n_112), .Y(n_181) );
INVx1_ASAP7_75t_L g490 ( .A(n_73), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_97), .B(n_452), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
INVx4_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_93), .Y(n_82) );
AO21x2_ASAP7_75t_L g687 ( .A1(n_83), .A2(n_640), .B(n_688), .Y(n_687) );
NAND2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_90), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_89), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_89), .Y(n_114) );
INVx3_ASAP7_75t_L g117 ( .A(n_89), .Y(n_117) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
INVx1_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
INVx2_ASAP7_75t_L g208 ( .A(n_89), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_89), .Y(n_210) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_89), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_90), .A2(n_110), .B1(n_115), .B2(n_118), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_90), .A2(n_118), .B1(n_133), .B2(n_136), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g145 ( .A1(n_90), .A2(n_146), .B1(n_148), .B2(n_150), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_90), .A2(n_118), .B1(n_158), .B2(n_162), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_90), .A2(n_180), .B(n_181), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_90), .A2(n_150), .B1(n_188), .B2(n_189), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_90), .A2(n_206), .B1(n_209), .B2(n_211), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_90), .A2(n_118), .B1(n_226), .B2(n_228), .Y(n_225) );
INVx6_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
O2A1O1Ixp5_ASAP7_75t_L g176 ( .A1(n_91), .A2(n_149), .B(n_177), .C(n_178), .Y(n_176) );
BUFx8_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
INVx1_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AO31x2_ASAP7_75t_L g144 ( .A1(n_94), .A2(n_145), .A3(n_152), .B(n_154), .Y(n_144) );
AO31x2_ASAP7_75t_L g156 ( .A1(n_94), .A2(n_157), .A3(n_165), .B(n_167), .Y(n_156) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_94), .A2(n_225), .A3(n_229), .B(n_230), .Y(n_224) );
BUFx10_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_96), .Y(n_641) );
INVxp67_ASAP7_75t_R g97 ( .A(n_98), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND3x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_349), .C(n_427), .Y(n_99) );
NOR2x1_ASAP7_75t_L g100 ( .A(n_101), .B(n_292), .Y(n_100) );
NAND3xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_239), .C(n_262), .Y(n_101) );
AOI221x1_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_169), .B1(n_192), .B2(n_201), .C(n_214), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_142), .Y(n_103) );
AND2x4_ASAP7_75t_L g329 ( .A(n_104), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_130), .Y(n_105) );
INVx2_ASAP7_75t_L g288 ( .A(n_106), .Y(n_288) );
INVx1_ASAP7_75t_L g315 ( .A(n_106), .Y(n_315) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g195 ( .A(n_107), .Y(n_195) );
AND2x4_ASAP7_75t_L g266 ( .A(n_107), .B(n_196), .Y(n_266) );
AO31x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_109), .A3(n_121), .B(n_127), .Y(n_107) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_108), .A2(n_152), .A3(n_187), .B(n_190), .Y(n_186) );
INVx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
INVx4_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AO31x2_ASAP7_75t_L g131 ( .A1(n_121), .A2(n_132), .A3(n_138), .B(n_140), .Y(n_131) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_SL g154 ( .A(n_123), .B(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_123), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g129 ( .A(n_124), .Y(n_129) );
INVx2_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_125), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_129), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g348 ( .A(n_130), .Y(n_348) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g196 ( .A(n_131), .Y(n_196) );
AND2x4_ASAP7_75t_L g237 ( .A(n_131), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g257 ( .A(n_131), .B(n_156), .Y(n_257) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_131), .Y(n_309) );
INVx1_ASAP7_75t_L g402 ( .A(n_131), .Y(n_402) );
AND2x2_ASAP7_75t_L g448 ( .A(n_131), .B(n_144), .Y(n_448) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_138), .A2(n_165), .A3(n_205), .B(n_212), .Y(n_204) );
INVx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_SL g182 ( .A(n_139), .Y(n_182) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_143), .B(n_314), .Y(n_313) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_143), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g442 ( .A(n_143), .B(n_340), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_143), .B(n_396), .Y(n_446) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_156), .Y(n_143) );
INVx4_ASAP7_75t_SL g198 ( .A(n_144), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_144), .B(n_200), .Y(n_250) );
BUFx2_ASAP7_75t_L g334 ( .A(n_144), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_144), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
BUFx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
INVx2_ASAP7_75t_L g238 ( .A(n_156), .Y(n_238) );
AND2x2_ASAP7_75t_L g240 ( .A(n_156), .B(n_195), .Y(n_240) );
INVx1_ASAP7_75t_L g265 ( .A(n_156), .Y(n_265) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_156), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_156), .B(n_348), .Y(n_379) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_166), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_SL g174 ( .A(n_166), .Y(n_174) );
INVx4_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_166), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_166), .B(n_231), .Y(n_230) );
INVxp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g423 ( .A(n_171), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_185), .Y(n_171) );
AND2x4_ASAP7_75t_L g218 ( .A(n_172), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g280 ( .A(n_172), .B(n_223), .Y(n_280) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx2_ASAP7_75t_L g366 ( .A(n_173), .Y(n_366) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_183), .Y(n_173) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_174), .A2(n_175), .B(n_183), .Y(n_253) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B(n_182), .Y(n_175) );
INVx2_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
AND2x4_ASAP7_75t_L g278 ( .A(n_185), .B(n_204), .Y(n_278) );
INVx3_ASAP7_75t_L g301 ( .A(n_185), .Y(n_301) );
INVx2_ASAP7_75t_L g322 ( .A(n_185), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_185), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_185), .B(n_222), .Y(n_416) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g203 ( .A(n_186), .B(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g217 ( .A(n_186), .Y(n_217) );
AND2x2_ASAP7_75t_L g295 ( .A(n_186), .B(n_219), .Y(n_295) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_197), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx3_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
AND2x2_ASAP7_75t_L g308 ( .A(n_195), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g377 ( .A(n_195), .B(n_198), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_196), .B(n_198), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_197), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g236 ( .A(n_198), .Y(n_236) );
AND2x2_ASAP7_75t_L g264 ( .A(n_198), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g282 ( .A(n_198), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g324 ( .A(n_198), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_198), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g385 ( .A(n_198), .Y(n_385) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_203), .B(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_SL g259 ( .A(n_203), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g338 ( .A(n_203), .B(n_221), .Y(n_338) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_203), .Y(n_373) );
INVx2_ASAP7_75t_L g390 ( .A(n_203), .Y(n_390) );
INVx2_ASAP7_75t_L g219 ( .A(n_204), .Y(n_219) );
OR2x2_ASAP7_75t_L g270 ( .A(n_204), .B(n_261), .Y(n_270) );
INVx1_ASAP7_75t_L g291 ( .A(n_204), .Y(n_291) );
BUFx2_ASAP7_75t_L g306 ( .A(n_204), .Y(n_306) );
OR2x2_ASAP7_75t_L g375 ( .A(n_204), .B(n_224), .Y(n_375) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_220), .B(n_233), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_215), .A2(n_297), .B(n_342), .C(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g241 ( .A(n_216), .B(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_216), .A2(n_275), .B1(n_441), .B2(n_442), .Y(n_440) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_L g232 ( .A(n_218), .Y(n_232) );
AND2x4_ASAP7_75t_L g360 ( .A(n_218), .B(n_269), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_218), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_232), .Y(n_220) );
INVx1_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g260 ( .A(n_222), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_223), .B(n_253), .Y(n_303) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g252 ( .A(n_224), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g269 ( .A(n_224), .Y(n_269) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_224), .Y(n_344) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g255 ( .A(n_235), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_236), .B(n_315), .Y(n_354) );
INVx2_ASAP7_75t_L g246 ( .A(n_237), .Y(n_246) );
AND2x2_ASAP7_75t_L g323 ( .A(n_237), .B(n_324), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_237), .B(n_287), .Y(n_368) );
AND2x2_ASAP7_75t_L g405 ( .A(n_237), .B(n_377), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_251), .B1(n_254), .B2(n_258), .Y(n_243) );
NOR2x1_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g449 ( .A(n_246), .Y(n_449) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g289 ( .A(n_252), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_252), .B(n_301), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_252), .B(n_295), .Y(n_386) );
AND2x4_ASAP7_75t_L g432 ( .A(n_252), .B(n_278), .Y(n_432) );
INVx1_ASAP7_75t_L g261 ( .A(n_253), .Y(n_261) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g438 ( .A(n_256), .B(n_334), .Y(n_438) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g371 ( .A(n_257), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g399 ( .A(n_257), .B(n_273), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_258), .B(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g380 ( .A(n_260), .B(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B1(n_271), .B2(n_275), .C(n_281), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g297 ( .A(n_264), .Y(n_297) );
AND2x2_ASAP7_75t_L g421 ( .A(n_264), .B(n_287), .Y(n_421) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
INVx3_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_266), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g355 ( .A(n_266), .B(n_356), .Y(n_355) );
NOR2xp67_ASAP7_75t_SL g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g294 ( .A(n_268), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_268), .B(n_301), .Y(n_363) );
AOI322xp5_ASAP7_75t_L g369 ( .A1(n_268), .A2(n_355), .A3(n_370), .B1(n_373), .B2(n_374), .C1(n_376), .C2(n_380), .Y(n_369) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g311 ( .A(n_269), .B(n_278), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_270), .B(n_322), .Y(n_321) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_270), .B(n_420), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_271), .A2(n_413), .B1(n_417), .B2(n_421), .Y(n_412) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx4_ASAP7_75t_L g396 ( .A(n_273), .Y(n_396) );
OR2x2_ASAP7_75t_L g426 ( .A(n_273), .B(n_401), .Y(n_426) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g439 ( .A(n_278), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_279), .B(n_305), .Y(n_326) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI211x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B(n_289), .C(n_290), .Y(n_281) );
INVx2_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g346 ( .A(n_287), .Y(n_346) );
NAND2x1_ASAP7_75t_L g437 ( .A(n_287), .B(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g343 ( .A(n_288), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g408 ( .A(n_290), .Y(n_408) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_310), .C(n_325), .Y(n_292) );
OAI211xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B(n_298), .C(n_308), .Y(n_293) );
INVx1_ASAP7_75t_L g307 ( .A(n_294), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_295), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g365 ( .A(n_295), .B(n_366), .Y(n_365) );
NAND2xp33_ASAP7_75t_L g388 ( .A(n_295), .B(n_336), .Y(n_388) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_307), .Y(n_298) );
INVx1_ASAP7_75t_L g434 ( .A(n_299), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_300), .B(n_304), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g381 ( .A(n_301), .Y(n_381) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_303), .Y(n_411) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_316), .B2(n_317), .C(n_320), .Y(n_310) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NOR2x1p5_ASAP7_75t_L g374 ( .A(n_322), .B(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g330 ( .A(n_324), .Y(n_330) );
AOI211xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_331), .C(n_341), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B1(n_337), .B2(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g420 ( .A(n_344), .Y(n_420) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_382), .C(n_403), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_361), .C(n_369), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B(n_357), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g451 ( .A(n_358), .B(n_419), .Y(n_451) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_360), .A2(n_398), .B(n_400), .Y(n_397) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
OR2x2_ASAP7_75t_L g389 ( .A(n_366), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_378), .Y(n_441) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g384 ( .A(n_379), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g394 ( .A(n_379), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_387), .B2(n_391), .C(n_397), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_383), .A2(n_429), .B(n_433), .Y(n_428) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI32xp33_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_396), .A3(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_398), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B(n_412), .C(n_422), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_435), .C(n_443), .Y(n_427) );
INVxp33_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI21xp33_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_439), .B(n_440), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B(n_450), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_636), .B2(n_642), .C(n_681), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_454), .A2(n_673), .B1(n_682), .B2(n_685), .Y(n_681) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_496), .B(n_527), .C(n_532), .Y(n_455) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_464), .Y(n_458) );
BUFx2_ASAP7_75t_L g486 ( .A(n_459), .Y(n_486) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x2_ASAP7_75t_L g470 ( .A(n_461), .B(n_463), .Y(n_470) );
INVx2_ASAP7_75t_L g474 ( .A(n_461), .Y(n_474) );
INVx1_ASAP7_75t_L g485 ( .A(n_461), .Y(n_485) );
BUFx2_ASAP7_75t_L g505 ( .A(n_461), .Y(n_505) );
OR2x2_ASAP7_75t_L g512 ( .A(n_461), .B(n_463), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_461), .B(n_462), .Y(n_519) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g473 ( .A(n_463), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g484 ( .A(n_463), .Y(n_484) );
INVx1_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
AND2x2_ASAP7_75t_L g492 ( .A(n_464), .B(n_483), .Y(n_492) );
AND2x4_ASAP7_75t_L g494 ( .A(n_464), .B(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_SL g500 ( .A(n_464), .B(n_469), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_479), .B(n_487), .Y(n_466) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x6_ASAP7_75t_L g487 ( .A(n_469), .B(n_488), .Y(n_487) );
BUFx3_ASAP7_75t_L g523 ( .A(n_469), .Y(n_523) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_473), .Y(n_495) );
BUFx3_ASAP7_75t_L g522 ( .A(n_473), .Y(n_522) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g526 ( .A(n_477), .Y(n_526) );
AND2x4_ASAP7_75t_L g525 ( .A(n_478), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_483), .B(n_488), .Y(n_632) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g506 ( .A(n_488), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_488), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_493), .B2(n_494), .Y(n_489) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_513), .B1(n_514), .B2(n_520), .C(n_521), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_513), .A2(n_599), .B(n_602), .Y(n_598) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx8_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_579), .C(n_625), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_566), .Y(n_533) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_549), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g593 ( .A(n_540), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_540), .B(n_542), .Y(n_605) );
INVx2_ASAP7_75t_L g583 ( .A(n_541), .Y(n_583) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g557 ( .A(n_542), .Y(n_557) );
OR2x2_ASAP7_75t_L g570 ( .A(n_542), .B(n_559), .Y(n_570) );
AND2x4_ASAP7_75t_L g607 ( .A(n_542), .B(n_593), .Y(n_607) );
INVx1_ASAP7_75t_L g572 ( .A(n_543), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
OR2x2_ASAP7_75t_L g629 ( .A(n_543), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .Y(n_543) );
OR2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g553 ( .A(n_545), .Y(n_553) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g562 ( .A(n_548), .Y(n_562) );
NAND2xp33_ASAP7_75t_SL g597 ( .A(n_548), .B(n_564), .Y(n_597) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVxp67_ASAP7_75t_L g565 ( .A(n_553), .Y(n_565) );
OR2x6_ASAP7_75t_L g554 ( .A(n_555), .B(n_565), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
BUFx3_ASAP7_75t_L g601 ( .A(n_556), .Y(n_601) );
INVx8_ASAP7_75t_L g623 ( .A(n_556), .Y(n_623) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x4_ASAP7_75t_L g577 ( .A(n_557), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVxp67_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
AND2x4_ASAP7_75t_L g584 ( .A(n_561), .B(n_585), .Y(n_584) );
AND2x6_ASAP7_75t_L g664 ( .A(n_561), .B(n_582), .Y(n_664) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND3x1_ASAP7_75t_L g613 ( .A(n_562), .B(n_614), .C(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x6_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
BUFx8_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g609 ( .A(n_577), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_594), .Y(n_579) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_582), .B(n_667), .C(n_670), .Y(n_666) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g588 ( .A(n_584), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g634 ( .A(n_584), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g631 ( .A(n_585), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g614 ( .A(n_586), .Y(n_614) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_598), .B1(n_610), .B2(n_616), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g670 ( .A(n_597), .Y(n_670) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx3_ASAP7_75t_L g619 ( .A(n_603), .Y(n_619) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g630 ( .A(n_604), .Y(n_630) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g624 ( .A(n_607), .Y(n_624) );
BUFx2_ASAP7_75t_L g635 ( .A(n_607), .Y(n_635) );
INVx1_ASAP7_75t_L g617 ( .A(n_608), .Y(n_617) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_616) );
INVx8_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_633), .Y(n_625) );
INVx8_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g672 ( .A(n_639), .Y(n_672) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_641), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g688 ( .A(n_641), .B(n_672), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_659), .B1(n_673), .B2(n_676), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_643), .A2(n_673), .B1(n_683), .B2(n_684), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_650), .B2(n_658), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_645) );
INVx1_ASAP7_75t_L g649 ( .A(n_646), .Y(n_649) );
INVx1_ASAP7_75t_L g648 ( .A(n_647), .Y(n_648) );
INVx1_ASAP7_75t_L g658 ( .A(n_650), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_657), .Y(n_650) );
INVx1_ASAP7_75t_SL g657 ( .A(n_651), .Y(n_657) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_654), .Y(n_656) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx12f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx12f_ASAP7_75t_L g683 ( .A(n_661), .Y(n_683) );
BUFx8_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B(n_666), .C(n_671), .Y(n_662) );
AND2x2_ASAP7_75t_L g680 ( .A(n_663), .B(n_666), .Y(n_680) );
INVx4_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g669 ( .A(n_665), .Y(n_669) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g679 ( .A(n_671), .Y(n_679) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g684 ( .A(n_678), .Y(n_684) );
OR2x6_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_686), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
endmodule