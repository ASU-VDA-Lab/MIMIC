module fake_jpeg_3872_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_12),
.B(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_47),
.B1(n_28),
.B2(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_63),
.B1(n_24),
.B2(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_61),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_22),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_36),
.B1(n_33),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_47),
.B1(n_38),
.B2(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_87),
.B1(n_90),
.B2(n_52),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_28),
.B1(n_18),
.B2(n_38),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_18),
.B1(n_27),
.B2(n_19),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_26),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_88),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_86),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_26),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_43),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_44),
.C(n_41),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_32),
.B1(n_52),
.B2(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_100),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_105),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_107),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_24),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_121),
.B1(n_122),
.B2(n_100),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_112),
.B1(n_83),
.B2(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_120),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_59),
.B1(n_41),
.B2(n_39),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_39),
.B1(n_44),
.B2(n_21),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_74),
.A2(n_59),
.B1(n_21),
.B2(n_20),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_20),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_98),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_121),
.B1(n_129),
.B2(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_134),
.B1(n_142),
.B2(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_140),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_85),
.B1(n_84),
.B2(n_91),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_113),
.B1(n_126),
.B2(n_93),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_83),
.B(n_92),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_152),
.B(n_124),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_77),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_146),
.Y(n_173)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_121),
.C(n_127),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_95),
.C(n_20),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_0),
.Y(n_151)
);

FAx1_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_21),
.CI(n_20),
.CON(n_152),
.SN(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_111),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_155),
.CI(n_159),
.CON(n_180),
.SN(n_180)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_105),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_23),
.B(n_35),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_86),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_161),
.B(n_163),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_162),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_169),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_109),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_117),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_168),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_124),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_102),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_122),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_182),
.B(n_35),
.C(n_25),
.D(n_104),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_35),
.B(n_2),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_20),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_126),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_187),
.B1(n_167),
.B2(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_113),
.B1(n_23),
.B2(n_104),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_132),
.B1(n_152),
.B2(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_23),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_152),
.B1(n_144),
.B2(n_142),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_35),
.B1(n_2),
.B2(n_1),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_150),
.B(n_155),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_212),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_152),
.B1(n_151),
.B2(n_132),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_219),
.B(n_193),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_8),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_104),
.B1(n_23),
.B2(n_25),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_183),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_1),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_177),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_180),
.B1(n_184),
.B2(n_171),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_231),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_172),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_235),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_169),
.C(n_182),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_243),
.C(n_223),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_202),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_247),
.B1(n_210),
.B2(n_201),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_9),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_240),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_16),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_6),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_3),
.C(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_211),
.B1(n_204),
.B2(n_217),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_5),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_212),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_227),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_223),
.B1(n_219),
.B2(n_199),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_229),
.B1(n_243),
.B2(n_226),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_265),
.C(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_207),
.B1(n_221),
.B2(n_198),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_240),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_221),
.B1(n_198),
.B2(n_203),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_205),
.C(n_213),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_283),
.B1(n_263),
.B2(n_259),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_230),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_274),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_237),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_241),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_244),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_245),
.B1(n_229),
.B2(n_249),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_273),
.B(n_255),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_301),
.B(n_302),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_257),
.B1(n_262),
.B2(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_268),
.B1(n_261),
.B2(n_258),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_276),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_11),
.Y(n_312)
);

NAND2x1_ASAP7_75t_SL g301 ( 
.A(n_275),
.B(n_258),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_225),
.B(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_296),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_285),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_311),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_307),
.B(n_290),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_310),
.B(n_314),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_272),
.B(n_244),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_11),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_12),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_13),
.C(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_13),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_294),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_320),
.B(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_319),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_292),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_294),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_322),
.B(n_308),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_327),
.B(n_319),
.Y(n_331)
);

NAND2x1p5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_311),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_298),
.Y(n_329)
);

A2O1A1O1Ixp25_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_333),
.B(n_330),
.C(n_298),
.D(n_323),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_326),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_330),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_332),
.C(n_291),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_13),
.B(n_14),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_14),
.B(n_15),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_15),
.Y(n_339)
);


endmodule