module fake_aes_1255_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
INVxp67_ASAP7_75t_SL g14 ( .A(n_12), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_5), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_17), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
OAI21x1_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_15), .B(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
BUFx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_18), .B1(n_19), .B2(n_16), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B(n_10), .Y(n_24) );
NAND3xp33_ASAP7_75t_SL g25 ( .A(n_24), .B(n_0), .C(n_1), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_1), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_2), .B(n_3), .Y(n_27) );
AOI322xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_2), .A3(n_3), .B1(n_4), .B2(n_7), .C1(n_8), .C2(n_26), .Y(n_28) );
endmodule