module fake_jpeg_22664_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_6),
.B(n_2),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_24),
.C(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_11),
.A2(n_4),
.B1(n_14),
.B2(n_10),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_13),
.B(n_12),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_10),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_10),
.C(n_13),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_15),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_24),
.B1(n_14),
.B2(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_11),
.B1(n_13),
.B2(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_33),
.B1(n_32),
.B2(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_33),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_41),
.B1(n_39),
.B2(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_26),
.Y(n_46)
);

AOI332xp33_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_12),
.A3(n_27),
.B1(n_43),
.B2(n_46),
.B3(n_47),
.C1(n_29),
.C2(n_25),
.Y(n_49)
);


endmodule