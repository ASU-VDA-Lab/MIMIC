module fake_jpeg_30727_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_15),
.A2(n_2),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_21),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_77),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_49),
.C(n_46),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_54),
.C(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_56),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_17),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_25),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_1),
.C(n_3),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_54),
.B1(n_55),
.B2(n_48),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_81),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_85),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_51),
.B1(n_48),
.B2(n_22),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_7),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_48),
.B1(n_51),
.B2(n_6),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_20),
.B1(n_40),
.B2(n_37),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_94),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_18),
.A3(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_41),
.B(n_14),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_1),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_106),
.C(n_110),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.C(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_3),
.C(n_6),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_19),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_7),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_11),
.C(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_24),
.C(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_12),
.C(n_26),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_120),
.B(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_30),
.C(n_27),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_119),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_113),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_126),
.B(n_124),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_122),
.B(n_116),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);


endmodule