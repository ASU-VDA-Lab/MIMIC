module fake_jpeg_18060_n_17 (n_3, n_2, n_1, n_0, n_4, n_17);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_17;

wire n_13;
wire n_11;
wire n_14;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_4),
.B(n_0),
.Y(n_5)
);

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_7),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_5),
.C(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_8),
.B(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_11),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_2),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_11),
.B(n_5),
.Y(n_14)
);

A2O1A1O1Ixp25_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_15),
.B(n_9),
.C(n_6),
.D(n_7),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_6),
.B(n_7),
.C(n_12),
.D(n_14),
.Y(n_17)
);


endmodule