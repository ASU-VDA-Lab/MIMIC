module fake_netlist_1_11217_n_674 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_674);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_674;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_564;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_423;
wire n_621;
wire n_666;
wire n_342;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_498;
wire n_597;
wire n_349;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g85 ( .A(n_80), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_53), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_19), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_77), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_17), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_44), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_51), .Y(n_91) );
NOR2xp33_ASAP7_75t_L g92 ( .A(n_13), .B(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_22), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_2), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_30), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_3), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_56), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_49), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_73), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_70), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_37), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_33), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_58), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_36), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_75), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_65), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_31), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_101), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_123), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_101), .B(n_0), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_97), .B(n_1), .Y(n_129) );
NAND2xp33_ASAP7_75t_R g130 ( .A(n_88), .B(n_35), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_98), .B(n_1), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_123), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_96), .B(n_39), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_123), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_108), .B(n_34), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_113), .B(n_3), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_89), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_118), .A2(n_40), .B(n_83), .Y(n_144) );
CKINVDCx11_ASAP7_75t_R g145 ( .A(n_109), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_87), .B(n_4), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_85), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_94), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_103), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_104), .A2(n_42), .B(n_82), .Y(n_154) );
INVxp67_ASAP7_75t_SL g155 ( .A(n_136), .Y(n_155) );
BUFx10_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_150), .B(n_111), .Y(n_157) );
BUFx6f_ASAP7_75t_SL g158 ( .A(n_128), .Y(n_158) );
NOR2xp33_ASAP7_75t_R g159 ( .A(n_130), .B(n_122), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_128), .A2(n_106), .B1(n_120), .B2(n_107), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_142), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_128), .B(n_121), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_136), .B(n_94), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_150), .B(n_124), .Y(n_164) );
NAND2xp33_ASAP7_75t_L g165 ( .A(n_135), .B(n_121), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_124), .B(n_95), .Y(n_169) );
NAND2xp33_ASAP7_75t_R g170 ( .A(n_129), .B(n_95), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_124), .B(n_105), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_125), .B(n_105), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
INVx4_ASAP7_75t_SL g175 ( .A(n_135), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_125), .B(n_88), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_132), .B(n_90), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_132), .B(n_90), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_127), .B(n_91), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
AND3x2_ASAP7_75t_L g188 ( .A(n_129), .B(n_117), .C(n_99), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_132), .B(n_91), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_135), .B(n_116), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_131), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_173), .B(n_132), .Y(n_194) );
INVxp33_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_173), .A2(n_138), .B1(n_135), .B2(n_153), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_159), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_140), .B1(n_146), .B2(n_143), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_164), .B(n_127), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_174), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_179), .B(n_146), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_174), .B(n_146), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_167), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_172), .B(n_134), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_156), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_180), .B(n_140), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_165), .B1(n_160), .B2(n_169), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_158), .Y(n_209) );
AND2x6_ASAP7_75t_SL g210 ( .A(n_163), .B(n_145), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_178), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_156), .B(n_134), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
INVx5_ASAP7_75t_L g215 ( .A(n_156), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_147), .B(n_149), .C(n_143), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_181), .B(n_141), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_162), .A2(n_151), .B(n_141), .C(n_148), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_156), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_190), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_166), .B(n_153), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_157), .B(n_153), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_175), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_188), .B(n_147), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_151), .B1(n_135), .B2(n_138), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_166), .B(n_147), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_193), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_166), .B(n_147), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_166), .B(n_149), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_175), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_166), .A2(n_138), .B1(n_135), .B2(n_149), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_166), .B(n_148), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_184), .B(n_148), .Y(n_234) );
NOR2xp67_ASAP7_75t_L g235 ( .A(n_187), .B(n_131), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_184), .B(n_138), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_175), .B(n_100), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g239 ( .A(n_187), .B(n_131), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_175), .B(n_154), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_184), .Y(n_241) );
NOR2x2_ASAP7_75t_L g242 ( .A(n_184), .B(n_138), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_184), .A2(n_138), .B1(n_152), .B2(n_131), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_184), .B(n_115), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_225), .A2(n_154), .B(n_152), .C(n_112), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_195), .B(n_7), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_205), .A2(n_144), .B(n_154), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_236), .A2(n_144), .B(n_182), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_203), .A2(n_144), .B(n_182), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_212), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_195), .B(n_9), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_211), .B(n_212), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_200), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_110), .B1(n_114), .B2(n_144), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_214), .B(n_144), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_194), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_226), .A2(n_176), .B(n_177), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_228), .A2(n_176), .B(n_177), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_217), .A2(n_92), .B1(n_126), .B2(n_133), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_199), .B(n_9), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_202), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_218), .A2(n_191), .B(n_189), .C(n_186), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_219), .A2(n_191), .B(n_189), .Y(n_265) );
CKINVDCx11_ASAP7_75t_R g266 ( .A(n_210), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_206), .A2(n_186), .B(n_185), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_207), .B(n_10), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_202), .B(n_138), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_215), .B(n_161), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_206), .A2(n_185), .B(n_161), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_207), .A2(n_138), .B1(n_187), .B2(n_161), .Y(n_273) );
AOI21x1_ASAP7_75t_L g274 ( .A1(n_240), .A2(n_167), .B(n_133), .Y(n_274) );
OAI22xp5_ASAP7_75t_SL g275 ( .A1(n_197), .A2(n_138), .B1(n_11), .B2(n_12), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_202), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_196), .A2(n_183), .B(n_139), .C(n_137), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_222), .A2(n_183), .B(n_168), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_207), .B(n_10), .Y(n_280) );
BUFx8_ASAP7_75t_SL g281 ( .A(n_198), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_215), .B(n_183), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_224), .Y(n_283) );
NOR2xp67_ASAP7_75t_SL g284 ( .A(n_215), .B(n_168), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_198), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_240), .A2(n_168), .B(n_139), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_240), .A2(n_168), .B(n_139), .Y(n_287) );
AND2x6_ASAP7_75t_L g288 ( .A(n_213), .B(n_137), .Y(n_288) );
BUFx2_ASAP7_75t_SL g289 ( .A(n_215), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_208), .B(n_137), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g291 ( .A(n_214), .B(n_133), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_209), .B(n_126), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_252), .A2(n_230), .B1(n_232), .B2(n_220), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_250), .B(n_238), .Y(n_296) );
AO31x2_ASAP7_75t_L g297 ( .A1(n_254), .A2(n_126), .A3(n_244), .B(n_234), .Y(n_297) );
BUFx10_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_247), .A2(n_221), .B(n_233), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_262), .B(n_238), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_264), .A2(n_243), .B(n_227), .C(n_231), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_286), .A2(n_229), .B(n_213), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_287), .A2(n_201), .B(n_241), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_265), .A2(n_201), .B(n_241), .Y(n_306) );
NOR2xp33_ASAP7_75t_SL g307 ( .A(n_270), .B(n_230), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_277), .A2(n_239), .B1(n_235), .B2(n_204), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_281), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_268), .A2(n_204), .B1(n_223), .B2(n_237), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_279), .A2(n_237), .B(n_223), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_246), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_267), .A2(n_237), .B(n_242), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_245), .A2(n_242), .B(n_47), .C(n_48), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_260), .Y(n_316) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_254), .A2(n_43), .B(n_81), .Y(n_317) );
AO21x1_ASAP7_75t_L g318 ( .A1(n_255), .A2(n_41), .B(n_79), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_269), .A2(n_12), .B(n_13), .C(n_14), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_248), .A2(n_50), .B(n_76), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_276), .Y(n_322) );
AO32x2_ASAP7_75t_L g323 ( .A1(n_275), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .Y(n_323) );
BUFx10_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_16), .B1(n_18), .B2(n_20), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
OA21x2_ASAP7_75t_L g327 ( .A1(n_249), .A2(n_54), .B(n_21), .Y(n_327) );
AO31x2_ASAP7_75t_L g328 ( .A1(n_261), .A2(n_18), .A3(n_84), .B(n_24), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g329 ( .A(n_292), .B(n_283), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_312), .A2(n_261), .B1(n_251), .B2(n_290), .C(n_269), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
AO221x2_ASAP7_75t_L g333 ( .A1(n_325), .A2(n_290), .B1(n_266), .B2(n_292), .C(n_255), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_326), .B(n_273), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_316), .B(n_278), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_300), .A2(n_272), .B(n_257), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_296), .A2(n_288), .B1(n_293), .B2(n_291), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_314), .A2(n_259), .B(n_282), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_299), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_321), .A2(n_271), .B(n_284), .Y(n_342) );
AO21x2_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_291), .B(n_288), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_301), .B(n_288), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_327), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_314), .A2(n_288), .B(n_25), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_327), .A2(n_288), .B(n_26), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_296), .A2(n_23), .B(n_27), .C(n_28), .Y(n_350) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_32), .A3(n_52), .B(n_55), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_295), .B(n_59), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_322), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_307), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_302), .B(n_71), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_320), .A2(n_302), .B(n_313), .C(n_306), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_297), .A3(n_311), .B(n_304), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_345), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_328), .Y(n_359) );
INVxp33_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_335), .B(n_328), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_346), .A2(n_308), .B(n_305), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_348), .B(n_327), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_335), .B(n_328), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_341), .B(n_297), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_331), .A2(n_310), .B1(n_329), .B2(n_308), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_317), .B(n_297), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_341), .B(n_297), .Y(n_369) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_310), .B(n_328), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_345), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_357), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_357), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_334), .B(n_298), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_357), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_323), .B(n_298), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_334), .B(n_323), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_332), .B(n_323), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_332), .B(n_323), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_336), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_376), .B(n_357), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_373), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_371), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_367), .A2(n_333), .B1(n_344), .B2(n_352), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_372), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_376), .B(n_351), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_375), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_369), .B(n_333), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_358), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_358), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_355), .B(n_352), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_360), .B(n_333), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_375), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_361), .B(n_351), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_376), .B(n_351), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_382), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_360), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_370), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_361), .B(n_351), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_361), .B(n_351), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_375), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_416), .B(n_359), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_393), .B(n_374), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
OR2x6_ASAP7_75t_L g428 ( .A(n_397), .B(n_364), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_416), .B(n_359), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_386), .B(n_359), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_386), .B(n_365), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_393), .B(n_378), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_394), .B(n_384), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_394), .B(n_365), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_402), .B(n_378), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_400), .B(n_365), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_398), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_400), .B(n_381), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_387), .B(n_381), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_402), .B(n_378), .Y(n_445) );
HB1xp67_ASAP7_75t_SL g446 ( .A(n_397), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_397), .B(n_385), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_381), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_388), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_387), .B(n_383), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_397), .B(n_385), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_387), .B(n_383), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_387), .B(n_383), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_406), .B(n_384), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_424), .B(n_382), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_412), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_424), .B(n_324), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_387), .B(n_370), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_410), .B(n_370), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_410), .B(n_370), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_390), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_403), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_422), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_388), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_417), .B(n_380), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_410), .B(n_370), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_403), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_417), .B(n_380), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_419), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_408), .B(n_324), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_420), .B(n_368), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_401), .B(n_388), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_420), .B(n_368), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_389), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_389), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_368), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_432), .B(n_401), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_475), .B(n_401), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_461), .B(n_421), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_429), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_446), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_457), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_461), .B(n_421), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_432), .B(n_421), .Y(n_490) );
OAI33xp33_ASAP7_75t_L g491 ( .A1(n_468), .A2(n_408), .A3(n_367), .B1(n_377), .B2(n_415), .B3(n_337), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_425), .B(n_415), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_463), .B(n_413), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_435), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_425), .B(n_391), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_471), .A2(n_413), .B(n_418), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_440), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_431), .B(n_422), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_475), .B(n_431), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_430), .B(n_389), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_440), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_463), .B(n_418), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_443), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_428), .B(n_385), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_469), .B(n_418), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_439), .B(n_423), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_459), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_473), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_469), .B(n_418), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_449), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_439), .B(n_423), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_447), .B(n_409), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_470), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_470), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_447), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_466), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_433), .B(n_423), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_444), .B(n_413), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_444), .B(n_414), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_451), .B(n_414), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_451), .B(n_414), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_453), .B(n_414), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_448), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_458), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_414), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_433), .B(n_419), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_458), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_441), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_455), .B(n_392), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_448), .B(n_392), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_437), .B(n_419), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_460), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_501), .B(n_438), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_482), .B(n_438), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_484), .B(n_474), .Y(n_545) );
INVx5_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_484), .B(n_474), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_486), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_489), .B(n_479), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_492), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_512), .B(n_442), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_489), .B(n_479), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_522), .B(n_428), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_498), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_494), .B(n_504), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_532), .B(n_476), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_482), .B(n_445), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_504), .B(n_454), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_499), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_496), .A2(n_333), .B1(n_476), .B2(n_460), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_493), .B(n_437), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_509), .B(n_445), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_509), .B(n_426), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_480), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_506), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_513), .B(n_454), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_513), .B(n_442), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_510), .B(n_426), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_488), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_428), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_527), .B(n_442), .C(n_456), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_481), .B(n_441), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_480), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_436), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_488), .Y(n_584) );
AOI21xp5_ASAP7_75t_SL g585 ( .A1(n_518), .A2(n_428), .B(n_452), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_521), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_526), .B(n_428), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_517), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_491), .B(n_442), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_544), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_559), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_562), .A2(n_552), .B1(n_589), .B2(n_546), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_589), .B(n_490), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_590), .B(n_545), .Y(n_595) );
OAI22xp33_ASAP7_75t_SL g596 ( .A1(n_546), .A2(n_508), .B1(n_518), .B2(n_522), .Y(n_596) );
AOI322xp5_ASAP7_75t_L g597 ( .A1(n_546), .A2(n_511), .A3(n_500), .B1(n_536), .B2(n_523), .C1(n_524), .C2(n_540), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_552), .A2(n_530), .B1(n_528), .B2(n_529), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_555), .A2(n_452), .B(n_497), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g600 ( .A1(n_555), .A2(n_452), .B(n_529), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_567), .A2(n_528), .B1(n_530), .B2(n_531), .C(n_534), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_543), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_546), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_555), .A2(n_534), .B1(n_531), .B2(n_515), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_548), .B(n_535), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_585), .A2(n_538), .B1(n_525), .B2(n_539), .C(n_502), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_551), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_553), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_550), .B(n_533), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_554), .B(n_533), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_561), .Y(n_614) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_585), .B(n_379), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_558), .A2(n_434), .B(n_517), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_573), .A2(n_434), .B(n_409), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g619 ( .A1(n_578), .A2(n_567), .B(n_582), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_576), .B(n_462), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_SL g621 ( .A1(n_582), .A2(n_377), .B(n_385), .C(n_462), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_581), .B(n_396), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g623 ( .A1(n_542), .A2(n_472), .A3(n_478), .B1(n_477), .B2(n_450), .C1(n_467), .C2(n_355), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_593), .A2(n_564), .B1(n_566), .B2(n_563), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_594), .A2(n_587), .B1(n_573), .B2(n_583), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_591), .B(n_577), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_596), .A2(n_541), .B(n_586), .Y(n_627) );
NOR2xp67_ASAP7_75t_SL g628 ( .A(n_600), .B(n_309), .Y(n_628) );
AOI221x1_ASAP7_75t_L g629 ( .A1(n_619), .A2(n_568), .B1(n_569), .B2(n_580), .C(n_570), .Y(n_629) );
AOI321xp33_ASAP7_75t_L g630 ( .A1(n_608), .A2(n_541), .A3(n_557), .B1(n_571), .B2(n_572), .C(n_579), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_599), .A2(n_571), .B(n_560), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_597), .A2(n_574), .B(n_385), .C(n_588), .Y(n_632) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_620), .B(n_588), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_597), .A2(n_584), .B(n_575), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_602), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_592), .B(n_575), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_601), .B(n_584), .C(n_379), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_616), .B(n_396), .Y(n_638) );
AOI221x1_ASAP7_75t_SL g639 ( .A1(n_595), .A2(n_396), .B1(n_472), .B2(n_477), .C(n_467), .Y(n_639) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_603), .A2(n_336), .A3(n_349), .B1(n_478), .B2(n_450), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_615), .A2(n_349), .B(n_396), .C(n_347), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_618), .A2(n_396), .B1(n_379), .B2(n_368), .Y(n_642) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_611), .A2(n_349), .A3(n_392), .B1(n_405), .B2(n_404), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_637), .B(n_623), .C(n_617), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_630), .B(n_598), .C(n_604), .D(n_621), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_632), .A2(n_612), .A3(n_609), .B(n_614), .Y(n_646) );
AND4x1_ASAP7_75t_L g647 ( .A(n_628), .B(n_610), .C(n_606), .D(n_607), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_629), .B(n_613), .C(n_622), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_639), .A2(n_605), .B1(n_354), .B2(n_353), .C(n_350), .Y(n_649) );
OAI21xp33_ASAP7_75t_SL g650 ( .A1(n_627), .A2(n_364), .B(n_620), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_626), .B(n_379), .Y(n_651) );
AOI221x1_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_340), .B1(n_338), .B2(n_405), .C(n_404), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_624), .A2(n_379), .B(n_364), .C(n_343), .Y(n_653) );
OAI221xp5_ASAP7_75t_SL g654 ( .A1(n_631), .A2(n_364), .B1(n_339), .B2(n_405), .C(n_404), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_654), .B(n_624), .C(n_641), .D(n_642), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_645), .B(n_625), .C(n_640), .D(n_638), .Y(n_656) );
AND5x1_ASAP7_75t_L g657 ( .A(n_646), .B(n_643), .C(n_633), .D(n_636), .E(n_635), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_644), .B(n_379), .Y(n_658) );
AND3x2_ASAP7_75t_L g659 ( .A(n_647), .B(n_351), .C(n_399), .Y(n_659) );
OAI22xp5_ASAP7_75t_SL g660 ( .A1(n_650), .A2(n_364), .B1(n_363), .B2(n_399), .Y(n_660) );
NOR5xp2_ASAP7_75t_L g661 ( .A(n_656), .B(n_648), .C(n_653), .D(n_649), .E(n_652), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_660), .A2(n_651), .B1(n_364), .B2(n_399), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_658), .B(n_343), .C(n_364), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_659), .B(n_407), .Y(n_664) );
OR5x1_ASAP7_75t_L g665 ( .A(n_663), .B(n_655), .C(n_657), .D(n_343), .E(n_407), .Y(n_665) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_662), .B(n_363), .Y(n_666) );
INVx3_ASAP7_75t_SL g667 ( .A(n_665), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
AOI22xp33_ASAP7_75t_R g669 ( .A1(n_668), .A2(n_661), .B1(n_664), .B2(n_363), .Y(n_669) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_667), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_363), .B1(n_342), .B2(n_407), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_669), .B(n_342), .C(n_407), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_342), .B(n_363), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_363), .B(n_342), .Y(n_674) );
endmodule