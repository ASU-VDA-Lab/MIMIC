module real_jpeg_19990_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI21xp33_ASAP7_75t_SL g28 ( 
.A1(n_0),
.A2(n_4),
.B(n_29),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_5),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_0),
.A2(n_4),
.B1(n_20),
.B2(n_39),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_6),
.B1(n_27),
.B2(n_39),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_20),
.B(n_27),
.C(n_28),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_27),
.B(n_44),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_1),
.A2(n_4),
.B1(n_20),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_3),
.A2(n_4),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_23),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_7),
.B1(n_21),
.B2(n_52),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_3),
.A2(n_4),
.B(n_7),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_8),
.B1(n_20),
.B2(n_36),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_5),
.B(n_39),
.C(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_34),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_8),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_8),
.B1(n_36),
.B2(n_52),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_20),
.B(n_52),
.C(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_76),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_75),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_13)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_30),
.B2(n_31),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_18),
.B1(n_41),
.B2(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_17),
.A2(n_18),
.B1(n_84),
.B2(n_87),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_17),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_18),
.B1(n_73),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_32),
.C(n_41),
.Y(n_31)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_18),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_18),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_18),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_18),
.B(n_49),
.C(n_85),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_20),
.A2(n_35),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_20),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_21),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_40),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_63),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_49),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_49),
.B1(n_81),
.B2(n_98),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_48),
.A2(n_56),
.B(n_105),
.C(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_48),
.A2(n_49),
.B1(n_71),
.B2(n_72),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_67),
.C(n_71),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_68),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_107),
.B(n_114),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_100),
.B(n_106),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_99),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_83),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);


endmodule