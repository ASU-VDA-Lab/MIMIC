module fake_netlist_1_8188_n_1001 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1001);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1001;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_243;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_947;
wire n_924;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
BUFx10_ASAP7_75t_L g237 ( .A(n_53), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_232), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_51), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_234), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_222), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_39), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_153), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_80), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_214), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_199), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_136), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_101), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
INVxp33_ASAP7_75t_R g254 ( .A(n_84), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_48), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_58), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_151), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_3), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_163), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_103), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_133), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_225), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_207), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_198), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_189), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_125), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_10), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_141), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_60), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_3), .Y(n_272) );
BUFx10_ASAP7_75t_L g273 ( .A(n_80), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_138), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_152), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_220), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_184), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_139), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_108), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_233), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_20), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_200), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_93), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_201), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_159), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_100), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_102), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_208), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_145), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_29), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_223), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_119), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_35), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_122), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_45), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_114), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_58), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_127), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_192), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_92), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_187), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_155), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_219), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_212), .Y(n_306) );
BUFx10_ASAP7_75t_L g307 ( .A(n_178), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_96), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_76), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_197), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_211), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_142), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_180), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_166), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_85), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_34), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_37), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_104), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_209), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_164), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_99), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g322 ( .A(n_30), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_38), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_82), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_128), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_213), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_217), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_173), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_38), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_161), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_74), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_21), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_75), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_117), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_156), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_172), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_30), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_190), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_236), .Y(n_339) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_57), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_230), .Y(n_341) );
BUFx10_ASAP7_75t_L g342 ( .A(n_165), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_154), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_191), .Y(n_344) );
CKINVDCx14_ASAP7_75t_R g345 ( .A(n_22), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_22), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_177), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_162), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_88), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_160), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_231), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_157), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_188), .Y(n_353) );
BUFx10_ASAP7_75t_L g354 ( .A(n_216), .Y(n_354) );
BUFx10_ASAP7_75t_L g355 ( .A(n_86), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_137), .Y(n_356) );
BUFx8_ASAP7_75t_SL g357 ( .A(n_210), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_115), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_59), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_185), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_175), .Y(n_361) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_307), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_277), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_277), .B(n_0), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_277), .Y(n_365) );
INVx5_ASAP7_75t_L g366 ( .A(n_344), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_240), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_246), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_262), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_238), .Y(n_371) );
OA21x2_ASAP7_75t_L g372 ( .A1(n_238), .A2(n_89), .B(n_87), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_255), .B(n_0), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_340), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_245), .B(n_2), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_357), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_252), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_253), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_305), .Y(n_380) );
INVx5_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_328), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_257), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_279), .B(n_5), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_239), .Y(n_385) );
INVx6_ASAP7_75t_L g386 ( .A(n_307), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_246), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_239), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_242), .Y(n_390) );
CKINVDCx11_ASAP7_75t_R g391 ( .A(n_256), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_258), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_326), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_340), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_242), .A2(n_91), .B(n_90), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_326), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_302), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_259), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_345), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_268), .Y(n_400) );
OAI22x1_ASAP7_75t_R g401 ( .A1(n_256), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
BUFx12f_ASAP7_75t_L g403 ( .A(n_342), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_377), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_380), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_382), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_362), .Y(n_409) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_362), .B(n_314), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_364), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_364), .Y(n_412) );
NOR2xp33_ASAP7_75t_R g413 ( .A(n_399), .B(n_345), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_391), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_369), .B(n_356), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_389), .B(n_272), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_389), .Y(n_417) );
NOR2xp33_ASAP7_75t_R g418 ( .A(n_403), .B(n_248), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_389), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_389), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_369), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_401), .Y(n_424) );
OA22x2_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_247), .B1(n_269), .B2(n_260), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_363), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_386), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_363), .Y(n_428) );
AND3x2_ASAP7_75t_L g429 ( .A(n_401), .B(n_254), .C(n_384), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_386), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_386), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_369), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_369), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_402), .B(n_354), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_367), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_365), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_375), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_378), .B(n_379), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_374), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_376), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_368), .Y(n_445) );
INVxp33_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_439), .B(n_394), .C(n_322), .Y(n_447) );
AO221x1_ASAP7_75t_L g448 ( .A1(n_422), .A2(n_263), .B1(n_267), .B2(n_266), .C(n_248), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_437), .B(n_383), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_442), .B(n_247), .C(n_241), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_432), .B(n_392), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_411), .B(n_398), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_445), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_412), .B(n_398), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_420), .B(n_400), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_438), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_433), .B(n_249), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_421), .B(n_249), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_404), .B(n_368), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_430), .B(n_250), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_431), .B(n_251), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_434), .B(n_251), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_441), .B(n_415), .C(n_414), .Y(n_467) );
INVxp33_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
BUFx5_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_417), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_408), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_431), .B(n_349), .Y(n_472) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_409), .B(n_263), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_427), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_410), .B(n_396), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_427), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_425), .B(n_396), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_425), .B(n_396), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_419), .A2(n_397), .B(n_395), .C(n_385), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_406), .B(n_299), .C(n_296), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_407), .B(n_237), .Y(n_484) );
AND2x6_ASAP7_75t_L g485 ( .A(n_436), .B(n_270), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_405), .B(n_354), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_424), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_429), .B(n_316), .C(n_309), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_424), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
BUFx6f_ASAP7_75t_SL g491 ( .A(n_443), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_443), .B(n_355), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_422), .B(n_355), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_416), .Y(n_494) );
NOR2xp67_ASAP7_75t_L g495 ( .A(n_409), .B(n_371), .Y(n_495) );
INVxp33_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_439), .B(n_332), .C(n_329), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_422), .B(n_243), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_430), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_428), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_422), .Y(n_501) );
NAND2xp33_ASAP7_75t_L g502 ( .A(n_411), .B(n_244), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_440), .B(n_385), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_410), .B(n_267), .Y(n_504) );
INVxp33_ASAP7_75t_L g505 ( .A(n_418), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_442), .B(n_337), .C(n_333), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_440), .B(n_388), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_440), .B(n_388), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_422), .Y(n_509) );
BUFx5_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_428), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_445), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_418), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_445), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g515 ( .A(n_409), .B(n_390), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_440), .B(n_390), .Y(n_516) );
AO221x1_ASAP7_75t_L g517 ( .A1(n_418), .A2(n_288), .B1(n_351), .B2(n_311), .C(n_359), .Y(n_517) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_409), .B(n_397), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_494), .A2(n_359), .B1(n_311), .B2(n_351), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_499), .B(n_465), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_503), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_499), .B(n_288), .Y(n_522) );
OR2x2_ASAP7_75t_SL g523 ( .A(n_501), .B(n_372), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_449), .B(n_346), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_495), .B(n_271), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_449), .A2(n_397), .B1(n_291), .B2(n_294), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_515), .B(n_282), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_503), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_512), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_470), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_506), .B(n_274), .Y(n_531) );
CKINVDCx8_ASAP7_75t_R g532 ( .A(n_504), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_512), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_512), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_507), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_474), .Y(n_536) );
AND2x6_ASAP7_75t_SL g537 ( .A(n_504), .B(n_317), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_508), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_518), .B(n_323), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_461), .A2(n_395), .B(n_372), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_489), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_516), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_447), .A2(n_331), .B1(n_324), .B2(n_278), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
BUFx3_ASAP7_75t_L g547 ( .A(n_484), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_451), .B(n_273), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_478), .A2(n_275), .B1(n_285), .B2(n_284), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_456), .B(n_273), .Y(n_551) );
BUFx4f_ASAP7_75t_SL g552 ( .A(n_493), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_461), .A2(n_454), .B(n_452), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_476), .Y(n_555) );
BUFx12f_ASAP7_75t_L g556 ( .A(n_475), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_485), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_450), .B(n_8), .Y(n_558) );
CKINVDCx11_ASAP7_75t_R g559 ( .A(n_446), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
AO22x1_ASAP7_75t_L g561 ( .A1(n_496), .A2(n_264), .B1(n_265), .B2(n_261), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_479), .A2(n_393), .B1(n_293), .B2(n_298), .Y(n_562) );
CKINVDCx11_ASAP7_75t_R g563 ( .A(n_505), .Y(n_563) );
OR2x2_ASAP7_75t_SL g564 ( .A(n_448), .B(n_372), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_511), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_476), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_479), .B(n_276), .Y(n_567) );
BUFx8_ASAP7_75t_L g568 ( .A(n_491), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_485), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_498), .Y(n_570) );
BUFx8_ASAP7_75t_L g571 ( .A(n_491), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_466), .B(n_280), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_467), .B(n_482), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_455), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_458), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_468), .B(n_281), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_497), .A2(n_304), .B1(n_308), .B2(n_306), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_517), .A2(n_393), .B1(n_312), .B2(n_319), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_477), .A2(n_334), .B1(n_335), .B2(n_318), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_486), .B(n_9), .Y(n_581) );
BUFx4f_ASAP7_75t_L g582 ( .A(n_485), .Y(n_582) );
AO22x2_ASAP7_75t_L g583 ( .A1(n_488), .A2(n_339), .B1(n_347), .B2(n_341), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_459), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_502), .B(n_283), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_460), .B(n_286), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_462), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_464), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_472), .B(n_287), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_510), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_492), .Y(n_592) );
INVx5_ASAP7_75t_L g593 ( .A(n_471), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_480), .B(n_9), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_481), .A2(n_352), .B1(n_353), .B2(n_350), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_471), .Y(n_596) );
INVx8_ASAP7_75t_L g597 ( .A(n_471), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_483), .Y(n_598) );
NOR2x2_ASAP7_75t_L g599 ( .A(n_490), .B(n_11), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_499), .B(n_289), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_449), .B(n_290), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_503), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_449), .B(n_292), .Y(n_603) );
NOR2x2_ASAP7_75t_L g604 ( .A(n_473), .B(n_11), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_461), .A2(n_361), .B(n_360), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_465), .B(n_297), .C(n_295), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_503), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_494), .B(n_300), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_449), .B(n_301), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_503), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_463), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_512), .Y(n_613) );
AND3x1_ASAP7_75t_L g614 ( .A(n_488), .B(n_12), .C(n_13), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_449), .B(n_303), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_449), .B(n_310), .Y(n_616) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_512), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_449), .B(n_313), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g619 ( .A1(n_494), .A2(n_320), .B1(n_321), .B2(n_315), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_512), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_509), .B(n_393), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_451), .A2(n_393), .B(n_327), .C(n_330), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_449), .B(n_325), .Y(n_623) );
INVx5_ASAP7_75t_L g624 ( .A(n_512), .Y(n_624) );
NAND2xp33_ASAP7_75t_L g625 ( .A(n_469), .B(n_336), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_495), .B(n_12), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_449), .B(n_338), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_513), .Y(n_628) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_473), .B(n_13), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_473), .B(n_14), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_521), .B(n_343), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_553), .A2(n_373), .B(n_370), .C(n_348), .Y(n_632) );
INVx5_ASAP7_75t_L g633 ( .A(n_597), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_528), .A2(n_358), .B1(n_381), .B2(n_366), .Y(n_634) );
NOR2xp33_ASAP7_75t_SL g635 ( .A(n_629), .B(n_366), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_532), .B(n_15), .Y(n_636) );
AND2x6_ASAP7_75t_SL g637 ( .A(n_574), .B(n_16), .Y(n_637) );
OAI22x1_ASAP7_75t_L g638 ( .A1(n_604), .A2(n_19), .B1(n_17), .B2(n_18), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g639 ( .A(n_579), .B(n_17), .C(n_18), .Y(n_639) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_613), .Y(n_640) );
BUFx12f_ASAP7_75t_L g641 ( .A(n_559), .Y(n_641) );
AOI22x1_ASAP7_75t_L g642 ( .A1(n_594), .A2(n_605), .B1(n_541), .B2(n_592), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_535), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_613), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_567), .A2(n_381), .B(n_366), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_563), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_547), .B(n_20), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_538), .A2(n_545), .B1(n_602), .B2(n_543), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_568), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_536), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_607), .B(n_370), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_610), .B(n_23), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_612), .A2(n_373), .B1(n_26), .B2(n_24), .Y(n_653) );
AO32x1_ASAP7_75t_L g654 ( .A1(n_523), .A2(n_373), .A3(n_25), .B1(n_26), .B2(n_27), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_568), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_571), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_520), .B(n_24), .Y(n_657) );
OR2x6_ASAP7_75t_L g658 ( .A(n_539), .B(n_25), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_630), .B(n_373), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_549), .Y(n_660) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_613), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_522), .B(n_28), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_598), .A2(n_95), .B(n_94), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_619), .B(n_31), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_526), .B(n_32), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_582), .B(n_33), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_537), .B(n_33), .Y(n_667) );
AOI22xp5_ASAP7_75t_SL g668 ( .A1(n_628), .A2(n_36), .B1(n_39), .B2(n_40), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_582), .B(n_40), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_601), .A2(n_98), .B(n_97), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_546), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_537), .B(n_41), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_519), .B(n_42), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_560), .A2(n_43), .B(n_44), .C(n_45), .Y(n_674) );
INVx5_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_597), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_574), .B(n_46), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_624), .B(n_47), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_544), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_624), .B(n_49), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_603), .A2(n_106), .B(n_105), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_556), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_565), .B(n_50), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_530), .B(n_50), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_584), .B(n_52), .Y(n_685) );
AO21x1_ASAP7_75t_L g686 ( .A1(n_626), .A2(n_109), .B(n_107), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_609), .A2(n_111), .B(n_110), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_524), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_615), .A2(n_113), .B(n_112), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_616), .A2(n_118), .B(n_116), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_611), .Y(n_691) );
BUFx12f_ASAP7_75t_L g692 ( .A(n_542), .Y(n_692) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_588), .A2(n_121), .B(n_120), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_618), .A2(n_124), .B(n_123), .Y(n_694) );
HAxp5_ASAP7_75t_L g695 ( .A(n_599), .B(n_57), .CON(n_695), .SN(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_623), .A2(n_129), .B(n_126), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_570), .B(n_61), .Y(n_697) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_617), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_578), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_550), .B(n_63), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_557), .B(n_64), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_555), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_558), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_550), .A2(n_65), .B(n_66), .C(n_67), .Y(n_704) );
CKINVDCx11_ASAP7_75t_R g705 ( .A(n_589), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_548), .A2(n_65), .B(n_67), .C(n_68), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_551), .A2(n_68), .B(n_69), .C(n_70), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_552), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_587), .B(n_69), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g710 ( .A1(n_622), .A2(n_170), .B(n_229), .C(n_228), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_578), .B(n_71), .Y(n_711) );
INVx4_ASAP7_75t_L g712 ( .A(n_593), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_608), .B(n_71), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_627), .A2(n_171), .B(n_226), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_569), .B(n_72), .Y(n_715) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_617), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_540), .A2(n_73), .B(n_74), .C(n_75), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_525), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_525), .B(n_77), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_617), .Y(n_720) );
INVx3_ASAP7_75t_L g721 ( .A(n_620), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_527), .B(n_78), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_620), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_620), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_527), .B(n_79), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_581), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_566), .B(n_83), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_595), .B(n_130), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_606), .B(n_132), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_596), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_621), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_562), .A2(n_134), .B(n_135), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_583), .B(n_140), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_580), .B(n_143), .Y(n_734) );
NAND2xp33_ASAP7_75t_L g735 ( .A(n_596), .B(n_144), .Y(n_735) );
AND2x6_ASAP7_75t_L g736 ( .A(n_591), .B(n_146), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_625), .A2(n_147), .B(n_148), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_561), .B(n_149), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_575), .Y(n_739) );
INVx3_ASAP7_75t_L g740 ( .A(n_529), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_577), .B(n_150), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_576), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_531), .B(n_158), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_573), .A2(n_167), .B(n_168), .C(n_169), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_533), .Y(n_745) );
NOR2xp67_ASAP7_75t_L g746 ( .A(n_586), .B(n_174), .Y(n_746) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_596), .Y(n_747) );
OR2x6_ASAP7_75t_L g748 ( .A(n_583), .B(n_176), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_564), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_614), .B(n_182), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_590), .B(n_183), .C(n_186), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_600), .B(n_235), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_534), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_614), .B(n_193), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_534), .Y(n_755) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_585), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_554), .B(n_205), .Y(n_757) );
BUFx12f_ASAP7_75t_L g758 ( .A(n_656), .Y(n_758) );
AO21x2_ASAP7_75t_L g759 ( .A1(n_632), .A2(n_572), .B(n_554), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_643), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_730), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_648), .A2(n_572), .B(n_554), .Y(n_762) );
OAI21x1_ASAP7_75t_L g763 ( .A1(n_693), .A2(n_572), .B(n_206), .Y(n_763) );
INVx6_ASAP7_75t_L g764 ( .A(n_633), .Y(n_764) );
INVx5_ASAP7_75t_SL g765 ( .A(n_658), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_695), .B(n_215), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_660), .Y(n_767) );
NAND2x1p5_ASAP7_75t_L g768 ( .A(n_675), .B(n_218), .Y(n_768) );
BUFx12f_ASAP7_75t_L g769 ( .A(n_641), .Y(n_769) );
NAND2x1p5_ASAP7_75t_L g770 ( .A(n_676), .B(n_712), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_692), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g772 ( .A(n_655), .Y(n_772) );
BUFx2_ASAP7_75t_SL g773 ( .A(n_649), .Y(n_773) );
AO21x2_ASAP7_75t_L g774 ( .A1(n_663), .A2(n_659), .B(n_732), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g775 ( .A1(n_652), .A2(n_703), .B(n_665), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_676), .Y(n_776) );
AOI22x1_ASAP7_75t_L g777 ( .A1(n_687), .A2(n_689), .B1(n_694), .B2(n_714), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_721), .A2(n_737), .B(n_651), .Y(n_778) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_747), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_640), .Y(n_780) );
BUFx12f_ASAP7_75t_L g781 ( .A(n_646), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_739), .B(n_742), .Y(n_782) );
OR3x4_ASAP7_75t_SL g783 ( .A(n_637), .B(n_638), .C(n_668), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_708), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_700), .A2(n_683), .B(n_690), .Y(n_785) );
OA21x2_ASAP7_75t_L g786 ( .A1(n_749), .A2(n_743), .B(n_696), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_711), .B(n_673), .Y(n_787) );
OAI21x1_ASAP7_75t_L g788 ( .A1(n_720), .A2(n_724), .B(n_723), .Y(n_788) );
INVx6_ASAP7_75t_SL g789 ( .A(n_748), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_691), .Y(n_790) );
BUFx12f_ASAP7_75t_L g791 ( .A(n_682), .Y(n_791) );
OAI21x1_ASAP7_75t_SL g792 ( .A1(n_728), .A2(n_731), .B(n_738), .Y(n_792) );
BUFx4_ASAP7_75t_SL g793 ( .A(n_757), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_718), .B(n_650), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_671), .A2(n_645), .B(n_744), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_740), .A2(n_755), .B(n_751), .Y(n_796) );
AO21x2_ASAP7_75t_L g797 ( .A1(n_710), .A2(n_639), .B(n_746), .Y(n_797) );
INVx8_ASAP7_75t_L g798 ( .A(n_685), .Y(n_798) );
AND2x2_ASAP7_75t_SL g799 ( .A(n_635), .B(n_697), .Y(n_799) );
AO21x2_ASAP7_75t_L g800 ( .A1(n_735), .A2(n_715), .B(n_678), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_680), .Y(n_801) );
AO21x2_ASAP7_75t_L g802 ( .A1(n_674), .A2(n_727), .B(n_653), .Y(n_802) );
BUFx2_ASAP7_75t_L g803 ( .A(n_702), .Y(n_803) );
AOI22x1_ASAP7_75t_L g804 ( .A1(n_752), .A2(n_750), .B1(n_754), .B2(n_745), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_631), .B(n_677), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_697), .Y(n_806) );
INVx4_ASAP7_75t_L g807 ( .A(n_705), .Y(n_807) );
AO21x2_ASAP7_75t_L g808 ( .A1(n_719), .A2(n_725), .B(n_722), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_644), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_713), .B(n_657), .Y(n_810) );
AO21x2_ASAP7_75t_L g811 ( .A1(n_729), .A2(n_734), .B(n_704), .Y(n_811) );
INVx6_ASAP7_75t_L g812 ( .A(n_753), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_657), .Y(n_813) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_644), .Y(n_814) );
AO21x2_ASAP7_75t_L g815 ( .A1(n_717), .A2(n_701), .B(n_726), .Y(n_815) );
INVx6_ASAP7_75t_L g816 ( .A(n_753), .Y(n_816) );
OAI21x1_ASAP7_75t_L g817 ( .A1(n_634), .A2(n_707), .B(n_706), .Y(n_817) );
INVx8_ASAP7_75t_L g818 ( .A(n_661), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_667), .B(n_672), .Y(n_819) );
AO21x2_ASAP7_75t_L g820 ( .A1(n_666), .A2(n_669), .B(n_688), .Y(n_820) );
BUFx2_ASAP7_75t_SL g821 ( .A(n_736), .Y(n_821) );
BUFx8_ASAP7_75t_L g822 ( .A(n_733), .Y(n_822) );
AO21x2_ASAP7_75t_L g823 ( .A1(n_654), .A2(n_741), .B(n_699), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_698), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_698), .Y(n_825) );
INVx5_ASAP7_75t_SL g826 ( .A(n_716), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_636), .B(n_647), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_654), .A2(n_736), .B(n_664), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_679), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_662), .Y(n_830) );
BUFx4f_ASAP7_75t_L g831 ( .A(n_756), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_684), .A2(n_709), .B(n_642), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_633), .B(n_675), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_632), .A2(n_553), .B(n_594), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_711), .A2(n_630), .B1(n_629), .B2(n_748), .Y(n_835) );
NAND2x1p5_ASAP7_75t_L g836 ( .A(n_633), .B(n_675), .Y(n_836) );
OAI21x1_ASAP7_75t_SL g837 ( .A1(n_686), .A2(n_648), .B(n_663), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_643), .B(n_521), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_643), .B(n_521), .Y(n_839) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_730), .Y(n_840) );
AOI22x1_ASAP7_75t_L g841 ( .A1(n_670), .A2(n_681), .B1(n_689), .B2(n_687), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_632), .A2(n_553), .B(n_594), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_643), .B(n_521), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_790), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_831), .A2(n_835), .B1(n_789), .B2(n_829), .Y(n_845) );
BUFx12f_ASAP7_75t_L g846 ( .A(n_769), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_782), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_758), .Y(n_848) );
INVx6_ASAP7_75t_L g849 ( .A(n_764), .Y(n_849) );
INVx4_ASAP7_75t_L g850 ( .A(n_833), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_819), .B(n_838), .Y(n_851) );
AO21x2_ASAP7_75t_L g852 ( .A1(n_837), .A2(n_762), .B(n_792), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_805), .B(n_787), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_839), .Y(n_854) );
OR2x6_ASAP7_75t_L g855 ( .A(n_798), .B(n_821), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_822), .A2(n_799), .B1(n_830), .B2(n_810), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_843), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_767), .Y(n_858) );
INVx4_ASAP7_75t_L g859 ( .A(n_833), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_836), .Y(n_860) );
INVx2_ASAP7_75t_SL g861 ( .A(n_764), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_801), .B(n_767), .Y(n_862) );
BUFx4f_ASAP7_75t_SL g863 ( .A(n_781), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_760), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_813), .A2(n_765), .B1(n_827), .B2(n_804), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_803), .B(n_776), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_775), .A2(n_798), .B1(n_815), .B2(n_766), .Y(n_867) );
BUFx8_ASAP7_75t_SL g868 ( .A(n_771), .Y(n_868) );
CKINVDCx11_ASAP7_75t_R g869 ( .A(n_791), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_775), .A2(n_815), .B1(n_808), .B2(n_806), .Y(n_870) );
INVx4_ASAP7_75t_L g871 ( .A(n_770), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_793), .Y(n_872) );
CKINVDCx11_ASAP7_75t_R g873 ( .A(n_772), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_779), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_783), .A2(n_807), .B1(n_828), .B2(n_768), .Y(n_875) );
OA21x2_ASAP7_75t_L g876 ( .A1(n_796), .A2(n_832), .B(n_785), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_794), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_814), .Y(n_878) );
INVx8_ASAP7_75t_L g879 ( .A(n_818), .Y(n_879) );
CKINVDCx6p67_ASAP7_75t_R g880 ( .A(n_773), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_820), .A2(n_802), .B1(n_842), .B2(n_834), .Y(n_881) );
INVx5_ASAP7_75t_L g882 ( .A(n_818), .Y(n_882) );
OAI21x1_ASAP7_75t_L g883 ( .A1(n_795), .A2(n_763), .B(n_778), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_784), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_788), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_869), .Y(n_886) );
AO32x1_ASAP7_75t_L g887 ( .A1(n_885), .A2(n_824), .A3(n_809), .B1(n_823), .B2(n_786), .Y(n_887) );
CKINVDCx10_ASAP7_75t_R g888 ( .A(n_863), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_858), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_871), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_851), .B(n_826), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_847), .B(n_811), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_855), .B(n_780), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_853), .A2(n_800), .B1(n_774), .B2(n_817), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_856), .A2(n_812), .B1(n_816), .B2(n_780), .Y(n_895) );
CKINVDCx16_ASAP7_75t_R g896 ( .A(n_846), .Y(n_896) );
OR2x6_ASAP7_75t_L g897 ( .A(n_879), .B(n_816), .Y(n_897) );
BUFx3_ASAP7_75t_L g898 ( .A(n_880), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_877), .B(n_800), .Y(n_899) );
CKINVDCx16_ASAP7_75t_R g900 ( .A(n_872), .Y(n_900) );
NOR2xp33_ASAP7_75t_R g901 ( .A(n_873), .B(n_825), .Y(n_901) );
BUFx8_ASAP7_75t_SL g902 ( .A(n_868), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_868), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_866), .B(n_825), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_845), .A2(n_797), .B1(n_841), .B2(n_777), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_864), .Y(n_906) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_879), .Y(n_907) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_882), .Y(n_908) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_882), .Y(n_909) );
CKINVDCx16_ASAP7_75t_R g910 ( .A(n_850), .Y(n_910) );
NOR2xp33_ASAP7_75t_R g911 ( .A(n_884), .B(n_840), .Y(n_911) );
NAND2xp33_ASAP7_75t_L g912 ( .A(n_882), .B(n_761), .Y(n_912) );
NOR2xp33_ASAP7_75t_R g913 ( .A(n_848), .B(n_761), .Y(n_913) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_874), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_844), .Y(n_915) );
INVx4_ASAP7_75t_L g916 ( .A(n_882), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_914), .B(n_881), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_890), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_889), .B(n_852), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_889), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_899), .B(n_881), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_892), .B(n_870), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_906), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_902), .Y(n_924) );
OAI22xp5_ASAP7_75t_SL g925 ( .A1(n_900), .A2(n_875), .B1(n_865), .B2(n_859), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_915), .B(n_852), .Y(n_926) );
BUFx3_ASAP7_75t_L g927 ( .A(n_908), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_910), .A2(n_871), .B1(n_867), .B2(n_865), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_911), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_894), .B(n_878), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_904), .B(n_878), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_887), .Y(n_932) );
INVx2_ASAP7_75t_SL g933 ( .A(n_913), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_887), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_887), .Y(n_935) );
INVx3_ASAP7_75t_L g936 ( .A(n_916), .Y(n_936) );
AND2x4_ASAP7_75t_L g937 ( .A(n_919), .B(n_905), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_923), .Y(n_938) );
AND2x4_ASAP7_75t_L g939 ( .A(n_919), .B(n_883), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_921), .B(n_876), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_921), .B(n_876), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_920), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_918), .Y(n_943) );
BUFx2_ASAP7_75t_L g944 ( .A(n_918), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_925), .A2(n_891), .B1(n_862), .B2(n_895), .Y(n_945) );
CKINVDCx16_ASAP7_75t_R g946 ( .A(n_933), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_925), .A2(n_862), .B1(n_854), .B2(n_857), .Y(n_947) );
AND2x4_ASAP7_75t_L g948 ( .A(n_926), .B(n_893), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_922), .B(n_759), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_917), .B(n_759), .Y(n_950) );
NAND3xp33_ASAP7_75t_SL g951 ( .A(n_928), .B(n_903), .C(n_901), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_938), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_940), .B(n_930), .Y(n_953) );
NOR3xp33_ASAP7_75t_SL g954 ( .A(n_951), .B(n_896), .C(n_886), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_943), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_942), .Y(n_956) );
NAND2xp5_ASAP7_75t_SL g957 ( .A(n_946), .B(n_929), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_941), .B(n_931), .Y(n_958) );
CKINVDCx16_ASAP7_75t_R g959 ( .A(n_946), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_943), .Y(n_960) );
NAND2xp5_ASAP7_75t_SL g961 ( .A(n_945), .B(n_929), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_949), .B(n_931), .Y(n_962) );
AND2x4_ASAP7_75t_L g963 ( .A(n_939), .B(n_932), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_944), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_949), .B(n_934), .Y(n_965) );
AND2x4_ASAP7_75t_L g966 ( .A(n_939), .B(n_935), .Y(n_966) );
OAI211xp5_ASAP7_75t_L g967 ( .A1(n_961), .A2(n_957), .B(n_947), .C(n_954), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_952), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_952), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_963), .B(n_948), .Y(n_970) );
INVx1_ASAP7_75t_SL g971 ( .A(n_959), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_956), .Y(n_972) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_960), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_965), .B(n_950), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_956), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_972), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g977 ( .A1(n_967), .A2(n_964), .B(n_955), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_975), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_971), .A2(n_937), .B1(n_963), .B2(n_966), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_968), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_969), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_979), .B(n_970), .Y(n_982) );
O2A1O1Ixp33_ASAP7_75t_L g983 ( .A1(n_977), .A2(n_973), .B(n_898), .C(n_924), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_980), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_981), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_984), .Y(n_986) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_983), .Y(n_987) );
OA21x2_ASAP7_75t_L g988 ( .A1(n_987), .A2(n_985), .B(n_982), .Y(n_988) );
NOR2x1_ASAP7_75t_L g989 ( .A(n_986), .B(n_888), .Y(n_989) );
NOR3xp33_ASAP7_75t_L g990 ( .A(n_989), .B(n_916), .C(n_861), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_990), .B(n_988), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_991), .B(n_974), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_992), .B(n_976), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_993), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_994), .Y(n_995) );
AOI21xp5_ASAP7_75t_L g996 ( .A1(n_995), .A2(n_907), .B(n_978), .Y(n_996) );
AOI211xp5_ASAP7_75t_L g997 ( .A1(n_996), .A2(n_907), .B(n_909), .C(n_912), .Y(n_997) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_997), .B(n_909), .C(n_860), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_998), .A2(n_849), .B1(n_897), .B2(n_936), .Y(n_999) );
OR2x6_ASAP7_75t_L g1000 ( .A(n_999), .B(n_927), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_1000), .A2(n_958), .B1(n_953), .B2(n_962), .Y(n_1001) );
endmodule