module fake_jpeg_15430_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_6),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.C(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_4),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_46),
.B1(n_49),
.B2(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_5),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_7),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_7),
.B1(n_11),
.B2(n_9),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_13),
.B1(n_28),
.B2(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_33),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_19),
.B(n_14),
.Y(n_84)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_71),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_13),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_16),
.B1(n_19),
.B2(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_70),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_23),
.B(n_15),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_20),
.B(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_25),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_79),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_20),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_53),
.C(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_26),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_48),
.B1(n_19),
.B2(n_16),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_16),
.B1(n_19),
.B2(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_52),
.B1(n_58),
.B2(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_57),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_68),
.B1(n_56),
.B2(n_54),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_67),
.B(n_63),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_63),
.C(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_116),
.B1(n_117),
.B2(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_107),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_65),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_76),
.B1(n_71),
.B2(n_57),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_75),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_92),
.B1(n_91),
.B2(n_95),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_96),
.C(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_127),
.C(n_122),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_84),
.B(n_83),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_124),
.B(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_94),
.B1(n_86),
.B2(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_103),
.B1(n_111),
.B2(n_107),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_93),
.C(n_69),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_97),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_102),
.C(n_106),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_95),
.B(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_128),
.C(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_105),
.C(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_143),
.C(n_144),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_140),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_111),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_142),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_106),
.CI(n_120),
.CON(n_143),
.SN(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_102),
.C(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_148),
.A2(n_129),
.B(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_133),
.C(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_151),
.C(n_144),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_143),
.C(n_136),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_150),
.C(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_129),
.C(n_132),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_158),
.CI(n_159),
.CON(n_160),
.SN(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_153),
.C(n_149),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_160),
.Y(n_162)
);


endmodule