module fake_netlist_5_2458_n_1228 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1228);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1228;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_1222;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_1227;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_1110;
wire n_864;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_247;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_516;
wire n_498;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_640;
wire n_275;
wire n_624;
wire n_252;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_1049;
wire n_992;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1100;
wire n_1207;
wire n_1214;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_833;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_428;
wire n_297;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_1225;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_580;
wire n_290;
wire n_221;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_1223;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_1165;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1122;
wire n_1111;
wire n_1197;
wire n_1211;
wire n_1226;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_781;
wire n_711;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_846;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_1224;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_1116;
wire n_954;
wire n_627;
wire n_1212;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_647;
wire n_407;
wire n_527;
wire n_237;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_1089;
wire n_927;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1032;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_34),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_12),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_90),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_28),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_31),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_32),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_105),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_80),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_89),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_21),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_66),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_26),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_16),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_63),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_64),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_9),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_37),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_13),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_134),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_41),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_56),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_5),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_91),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_33),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_112),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_96),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_29),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_117),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_22),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_35),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_20),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_118),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_119),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_125),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_183),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_150),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_93),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_69),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_113),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_140),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_87),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_52),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_26),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_120),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_85),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_123),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_84),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_19),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_115),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_76),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_0),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_171),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_81),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_86),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_109),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_145),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_65),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_185),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_138),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_55),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_49),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_135),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_40),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_193),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_197),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_197),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_262),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_1),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_300),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_193),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_250),
.B(n_1),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_190),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_241),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_194),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_250),
.B(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_288),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_2),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_288),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_199),
.B(n_3),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_213),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_235),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_215),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_221),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_186),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_200),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_3),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_203),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_206),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_211),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_189),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_194),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_224),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_240),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_216),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_218),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_223),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_227),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_228),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_234),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_230),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_198),
.B(n_4),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_253),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_192),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_244),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_226),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_226),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_233),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_258),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_263),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_245),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_266),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_248),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_195),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_251),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_261),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_205),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_208),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_299),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_268),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_270),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_269),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_272),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_289),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_299),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_271),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_209),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_233),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_254),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_254),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_285),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_327),
.B(n_188),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_196),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_349),
.A2(n_323),
.B(n_321),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_339),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_352),
.B(n_196),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_188),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

XNOR2x2_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_187),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

OA21x2_ASAP7_75t_L g423 ( 
.A1(n_358),
.A2(n_295),
.B(n_292),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_359),
.B(n_201),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_345),
.B(n_232),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

OR2x2_ASAP7_75t_SL g430 ( 
.A(n_313),
.B(n_296),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_370),
.B(n_372),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_311),
.B(n_287),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_335),
.B(n_302),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_317),
.B(n_287),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_331),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_201),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_319),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_202),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_202),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_396),
.A2(n_286),
.B(n_283),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_332),
.Y(n_442)
);

XNOR2x2_ASAP7_75t_R g443 ( 
.A(n_308),
.B(n_4),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_331),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_324),
.B(n_287),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_287),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_334),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_336),
.A2(n_293),
.B(n_298),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_366),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_367),
.B(n_287),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_306),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_337),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_314),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_413),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_273),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

OAI21xp33_ASAP7_75t_SL g473 ( 
.A1(n_397),
.A2(n_312),
.B(n_329),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_357),
.C(n_212),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_434),
.B(n_240),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_414),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_SL g484 ( 
.A1(n_397),
.A2(n_434),
.B(n_426),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_420),
.A2(n_322),
.B1(n_382),
.B2(n_240),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_433),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_442),
.B(n_337),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_240),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g497 ( 
.A(n_423),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_240),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_413),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_390),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_240),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_403),
.Y(n_512)
);

AND2x2_ASAP7_75t_SL g513 ( 
.A(n_433),
.B(n_435),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_433),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g516 ( 
.A(n_446),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_442),
.B(n_338),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_413),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_442),
.B(n_421),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_418),
.B(n_322),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_433),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_423),
.B(n_240),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_442),
.B(n_338),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_404),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_433),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_418),
.B(n_378),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_432),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_404),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_442),
.B(n_348),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_441),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_398),
.B(n_382),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_488),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_486),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_467),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_514),
.B(n_442),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

NOR3xp33_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_484),
.C(n_473),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_534),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_514),
.B(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_469),
.B(n_406),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_514),
.B(n_513),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_501),
.B(n_458),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_484),
.B(n_514),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_513),
.B(n_442),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_473),
.A2(n_434),
.B(n_398),
.C(n_427),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_469),
.B(n_406),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_474),
.A2(n_430),
.B1(n_427),
.B2(n_346),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_406),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_469),
.B(n_441),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_502),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_533),
.A2(n_420),
.B1(n_441),
.B2(n_452),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_521),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_514),
.B(n_461),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_521),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_467),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_513),
.B(n_441),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_510),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_511),
.B(n_458),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_513),
.B(n_442),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_467),
.B(n_441),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_504),
.Y(n_574)
);

BUFx12f_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_489),
.B(n_353),
.C(n_348),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_446),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_474),
.B(n_210),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_467),
.B(n_441),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_480),
.A2(n_461),
.B1(n_452),
.B2(n_438),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_472),
.B(n_452),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_488),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_477),
.B(n_503),
.Y(n_585)
);

OR2x2_ASAP7_75t_SL g586 ( 
.A(n_489),
.B(n_443),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_472),
.B(n_452),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_528),
.Y(n_588)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_452),
.Y(n_590)
);

INVx8_ASAP7_75t_L g591 ( 
.A(n_528),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_480),
.A2(n_452),
.B1(n_438),
.B2(n_364),
.Y(n_592)
);

AND2x6_ASAP7_75t_SL g593 ( 
.A(n_503),
.B(n_207),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_472),
.B(n_433),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_438),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_503),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_477),
.B(n_430),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_476),
.B(n_471),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_533),
.A2(n_430),
.B1(n_360),
.B2(n_381),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_L g600 ( 
.A1(n_499),
.A2(n_207),
.B1(n_238),
.B2(n_294),
.C(n_214),
.Y(n_600)
);

BUFx5_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_493),
.B(n_380),
.Y(n_602)
);

NAND2x1_ASAP7_75t_L g603 ( 
.A(n_476),
.B(n_422),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_493),
.B(n_391),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_499),
.B(n_214),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_353),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_479),
.B(n_435),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_506),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_479),
.B(n_435),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_522),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_515),
.B(n_356),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_470),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_470),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_477),
.B(n_356),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_480),
.A2(n_439),
.B1(n_440),
.B2(n_437),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_515),
.B(n_458),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_494),
.B(n_361),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_480),
.A2(n_439),
.B1(n_440),
.B2(n_437),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_470),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_470),
.Y(n_622)
);

INVxp33_ASAP7_75t_L g623 ( 
.A(n_496),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_490),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_477),
.B(n_361),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_515),
.B(n_458),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_618),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_611),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_612),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_538),
.B(n_480),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_538),
.B(n_533),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_564),
.A2(n_527),
.B(n_523),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_575),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_564),
.A2(n_523),
.B(n_594),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_543),
.A2(n_518),
.B1(n_310),
.B2(n_316),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_601),
.B(n_478),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_543),
.B(n_478),
.Y(n_637)
);

BUFx4f_ASAP7_75t_L g638 ( 
.A(n_591),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_623),
.B(n_494),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_585),
.B(n_551),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_545),
.A2(n_497),
.B(n_519),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_614),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_559),
.A2(n_548),
.B1(n_598),
.B2(n_585),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_617),
.B(n_517),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_560),
.B(n_464),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_542),
.A2(n_525),
.B(n_517),
.C(n_532),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_559),
.A2(n_518),
.B1(n_326),
.B2(n_328),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_615),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_601),
.B(n_525),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_552),
.A2(n_497),
.B(n_519),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_620),
.B(n_601),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_601),
.B(n_566),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_563),
.B(n_389),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_309),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_371),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_573),
.A2(n_497),
.B(n_496),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_561),
.B(n_371),
.Y(n_657)
);

CKINVDCx10_ASAP7_75t_R g658 ( 
.A(n_593),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_554),
.A2(n_497),
.B(n_491),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_595),
.B(n_373),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_580),
.A2(n_497),
.B(n_498),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_582),
.A2(n_507),
.B(n_498),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_607),
.A2(n_491),
.B(n_481),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_601),
.B(n_470),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_597),
.A2(n_524),
.B(n_507),
.C(n_487),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_542),
.B(n_475),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_621),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_609),
.A2(n_491),
.B(n_481),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_491),
.B(n_481),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_590),
.A2(n_524),
.B(n_487),
.Y(n_670)
);

AO21x2_ASAP7_75t_L g671 ( 
.A1(n_555),
.A2(n_424),
.B(n_416),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_622),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_565),
.A2(n_487),
.B(n_475),
.Y(n_673)
);

OAI321xp33_ASAP7_75t_L g674 ( 
.A1(n_553),
.A2(n_307),
.A3(n_369),
.B1(n_387),
.B2(n_420),
.C(n_464),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_562),
.B(n_457),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_597),
.A2(n_487),
.B(n_475),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_548),
.A2(n_294),
.B1(n_238),
.B2(n_416),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_537),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_596),
.B(n_424),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_540),
.B(n_475),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_618),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_586),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_606),
.A2(n_475),
.B1(n_487),
.B2(n_508),
.Y(n_683)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_606),
.A2(n_625),
.B(n_616),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_549),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_561),
.B(n_373),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_556),
.B(n_482),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_626),
.A2(n_508),
.B(n_481),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_603),
.A2(n_544),
.B(n_539),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_616),
.A2(n_500),
.B(n_495),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_591),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_550),
.A2(n_520),
.B(n_508),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_374),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_600),
.A2(n_377),
.B(n_374),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_625),
.A2(n_500),
.B(n_495),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_422),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_547),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_550),
.A2(n_520),
.B(n_508),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_422),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_588),
.B(n_425),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_576),
.B(n_377),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_379),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_571),
.A2(n_530),
.B(n_520),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_570),
.B(n_422),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_571),
.A2(n_500),
.B(n_495),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_546),
.A2(n_530),
.B(n_520),
.Y(n_709)
);

OAI21xp33_ASAP7_75t_L g710 ( 
.A1(n_572),
.A2(n_383),
.B(n_379),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_547),
.A2(n_530),
.B(n_492),
.Y(n_711)
);

AO22x1_ASAP7_75t_L g712 ( 
.A1(n_572),
.A2(n_385),
.B1(n_383),
.B2(n_301),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_574),
.B(n_482),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_557),
.B(n_605),
.Y(n_715)
);

AO21x1_ASAP7_75t_L g716 ( 
.A1(n_579),
.A2(n_445),
.B(n_492),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_581),
.A2(n_530),
.B1(n_445),
.B2(n_385),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_619),
.B(n_425),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_674),
.A2(n_557),
.B(n_613),
.C(n_602),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_SL g720 ( 
.A1(n_657),
.A2(n_687),
.B(n_704),
.C(n_705),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_677),
.A2(n_604),
.B(n_608),
.C(n_568),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_690),
.B(n_568),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_630),
.A2(n_592),
.B1(n_558),
.B2(n_610),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_694),
.Y(n_724)
);

OAI22x1_ASAP7_75t_L g725 ( 
.A1(n_654),
.A2(n_304),
.B1(n_298),
.B2(n_301),
.Y(n_725)
);

AO22x1_ASAP7_75t_L g726 ( 
.A1(n_696),
.A2(n_304),
.B1(n_457),
.B2(n_460),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_635),
.B(n_535),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_684),
.A2(n_583),
.B(n_536),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_642),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_694),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_636),
.A2(n_492),
.B(n_624),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_714),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_630),
.A2(n_584),
.B1(n_290),
.B2(n_457),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_669),
.A2(n_659),
.B(n_650),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_677),
.A2(n_425),
.B1(n_445),
.B2(n_448),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_662),
.A2(n_492),
.B(n_529),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_648),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_637),
.A2(n_431),
.B(n_425),
.C(n_447),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_631),
.B(n_447),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_635),
.B(n_431),
.C(n_219),
.Y(n_740)
);

O2A1O1Ixp5_ASAP7_75t_L g741 ( 
.A1(n_716),
.A2(n_445),
.B(n_492),
.C(n_453),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_667),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_646),
.A2(n_456),
.B(n_448),
.C(n_445),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_631),
.A2(n_462),
.B1(n_460),
.B2(n_463),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_633),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_640),
.B(n_447),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_678),
.B(n_447),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_643),
.B(n_447),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_690),
.B(n_460),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_694),
.B(n_462),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_627),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_686),
.B(n_407),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_627),
.B(n_217),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_679),
.A2(n_462),
.B(n_463),
.C(n_417),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_627),
.B(n_529),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_660),
.A2(n_220),
.B1(n_222),
.B2(n_225),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_644),
.A2(n_463),
.B(n_456),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_675),
.B(n_407),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_634),
.A2(n_529),
.B(n_485),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_628),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_643),
.A2(n_465),
.B1(n_453),
.B2(n_466),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_713),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_715),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_665),
.A2(n_531),
.B(n_512),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_641),
.A2(n_512),
.B(n_509),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_SL g768 ( 
.A(n_647),
.B(n_236),
.C(n_229),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_688),
.B(n_237),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_SL g770 ( 
.A1(n_666),
.A2(n_482),
.B(n_485),
.C(n_509),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_672),
.Y(n_771)
);

OA22x2_ASAP7_75t_L g772 ( 
.A1(n_697),
.A2(n_436),
.B1(n_410),
.B2(n_412),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_675),
.B(n_407),
.Y(n_773)
);

OA22x2_ASAP7_75t_L g774 ( 
.A1(n_647),
.A2(n_436),
.B1(n_410),
.B2(n_412),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

INVx5_ASAP7_75t_L g776 ( 
.A(n_688),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_688),
.B(n_242),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_689),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_649),
.A2(n_661),
.B(n_656),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_682),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_R g782 ( 
.A(n_638),
.B(n_655),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_720),
.B(n_645),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_767),
.A2(n_692),
.B(n_709),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_761),
.A2(n_668),
.B(n_663),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_746),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_719),
.A2(n_651),
.B(n_639),
.C(n_710),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_780),
.A2(n_666),
.B(n_676),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_765),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_760),
.B(n_638),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_764),
.A2(n_681),
.B1(n_652),
.B2(n_700),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_749),
.A2(n_695),
.A3(n_701),
.B(n_706),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_745),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_743),
.A2(n_632),
.B(n_673),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_721),
.A2(n_703),
.B(n_718),
.C(n_645),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_781),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_762),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_725),
.A2(n_712),
.B1(n_449),
.B2(n_409),
.C(n_417),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_775),
.B(n_778),
.Y(n_800)
);

AO31x2_ASAP7_75t_L g801 ( 
.A1(n_749),
.A2(n_691),
.A3(n_711),
.B(n_689),
.Y(n_801)
);

AO31x2_ASAP7_75t_L g802 ( 
.A1(n_763),
.A2(n_707),
.A3(n_702),
.B(n_699),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_727),
.B(n_779),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_753),
.Y(n_804)
);

AO21x1_ASAP7_75t_L g805 ( 
.A1(n_723),
.A2(n_733),
.B(n_758),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_723),
.A2(n_717),
.B(n_683),
.Y(n_806)
);

AOI21xp33_ASAP7_75t_L g807 ( 
.A1(n_740),
.A2(n_671),
.B(n_680),
.Y(n_807)
);

AO31x2_ASAP7_75t_L g808 ( 
.A1(n_763),
.A2(n_664),
.A3(n_680),
.B(n_531),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_768),
.A2(n_449),
.B(n_409),
.C(n_465),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_755),
.A2(n_453),
.B(n_465),
.C(n_466),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_736),
.A2(n_698),
.B(n_693),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_SL g812 ( 
.A1(n_754),
.A2(n_664),
.B(n_708),
.C(n_670),
.Y(n_812)
);

AO32x2_ASAP7_75t_L g813 ( 
.A1(n_733),
.A2(n_744),
.A3(n_774),
.B1(n_728),
.B2(n_741),
.Y(n_813)
);

AO31x2_ASAP7_75t_L g814 ( 
.A1(n_747),
.A2(n_531),
.A3(n_512),
.B(n_509),
.Y(n_814)
);

AO21x1_ASAP7_75t_L g815 ( 
.A1(n_758),
.A2(n_456),
.B(n_448),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_776),
.B(n_681),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_747),
.A2(n_681),
.B(n_671),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_738),
.A2(n_681),
.B(n_456),
.C(n_448),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_722),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_751),
.B(n_453),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_729),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_744),
.A2(n_466),
.B(n_465),
.C(n_419),
.Y(n_822)
);

AOI31xp67_ASAP7_75t_L g823 ( 
.A1(n_774),
.A2(n_509),
.A3(n_512),
.B(n_526),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_751),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_739),
.A2(n_529),
.B(n_485),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_759),
.A2(n_485),
.B(n_482),
.Y(n_826)
);

AO32x2_ASAP7_75t_L g827 ( 
.A1(n_728),
.A2(n_658),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_773),
.A2(n_448),
.B(n_456),
.C(n_466),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_734),
.A2(n_731),
.B(n_766),
.Y(n_829)
);

AO31x2_ASAP7_75t_L g830 ( 
.A1(n_748),
.A2(n_526),
.A3(n_415),
.B(n_407),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_726),
.B(n_408),
.Y(n_831)
);

AO31x2_ASAP7_75t_L g832 ( 
.A1(n_737),
.A2(n_526),
.A3(n_415),
.B(n_408),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_448),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_742),
.Y(n_834)
);

CKINVDCx11_ASAP7_75t_R g835 ( 
.A(n_724),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_771),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_SL g837 ( 
.A1(n_806),
.A2(n_772),
.B1(n_776),
.B2(n_750),
.Y(n_837)
);

CKINVDCx11_ASAP7_75t_R g838 ( 
.A(n_835),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_808),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_788),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_SL g841 ( 
.A1(n_803),
.A2(n_772),
.B1(n_776),
.B2(n_750),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_790),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_800),
.A2(n_757),
.B1(n_776),
.B2(n_722),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_805),
.A2(n_777),
.B1(n_769),
.B2(n_735),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_808),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_823),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_816),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_820),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_824),
.B(n_752),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_783),
.A2(n_799),
.B1(n_833),
.B2(n_789),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_787),
.B(n_752),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_794),
.B(n_766),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_791),
.A2(n_797),
.B1(n_786),
.B2(n_819),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_792),
.A2(n_724),
.B1(n_730),
.B2(n_264),
.Y(n_854)
);

BUFx4f_ASAP7_75t_SL g855 ( 
.A(n_836),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_SL g856 ( 
.A1(n_798),
.A2(n_730),
.B1(n_724),
.B2(n_756),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_813),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_832),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_832),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_831),
.A2(n_730),
.B1(n_456),
.B2(n_756),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_821),
.A2(n_252),
.B1(n_255),
.B2(n_259),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_793),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_804),
.B(n_454),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_834),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_832),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_795),
.A2(n_756),
.B1(n_265),
.B2(n_275),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_813),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_804),
.A2(n_260),
.B1(n_277),
.B2(n_280),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_809),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_SL g871 ( 
.A1(n_796),
.A2(n_408),
.B(n_411),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_807),
.A2(n_756),
.B1(n_454),
.B2(n_455),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_815),
.A2(n_459),
.B1(n_454),
.B2(n_455),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_830),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_830),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_811),
.A2(n_827),
.B1(n_829),
.B2(n_817),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_812),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_818),
.A2(n_282),
.B1(n_291),
.B2(n_297),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_828),
.A2(n_428),
.B1(n_408),
.B2(n_411),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_814),
.Y(n_880)
);

CKINVDCx11_ASAP7_75t_R g881 ( 
.A(n_827),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_814),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_808),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_814),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_830),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_826),
.A2(n_419),
.B(n_411),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_801),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_810),
.Y(n_888)
);

HB1xp67_ASAP7_75t_SL g889 ( 
.A(n_827),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_801),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_785),
.A2(n_784),
.B1(n_825),
.B2(n_454),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_801),
.A2(n_454),
.B1(n_455),
.B2(n_459),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_802),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_875),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_874),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_857),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_862),
.A2(n_822),
.B(n_802),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_857),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_857),
.Y(n_899)
);

OAI21x1_ASAP7_75t_L g900 ( 
.A1(n_862),
.A2(n_802),
.B(n_793),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_880),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_862),
.B(n_793),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_880),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_875),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_857),
.B(n_5),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_882),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_857),
.B(n_411),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_852),
.B(n_770),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_887),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_863),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_887),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_863),
.B(n_6),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_884),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_884),
.Y(n_914)
);

CKINVDCx8_ASAP7_75t_R g915 ( 
.A(n_863),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_839),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_839),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_893),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_845),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_882),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_858),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_845),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_838),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_893),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_890),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_858),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_863),
.B(n_7),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_863),
.Y(n_930)
);

OA21x2_ASAP7_75t_L g931 ( 
.A1(n_900),
.A2(n_885),
.B(n_874),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_905),
.B(n_848),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_908),
.B(n_852),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_910),
.B(n_868),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_905),
.A2(n_844),
.B(n_850),
.C(n_853),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_897),
.A2(n_867),
.B(n_871),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_923),
.A2(n_843),
.B1(n_870),
.B2(n_881),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_916),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_923),
.A2(n_870),
.B1(n_881),
.B2(n_855),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_896),
.B(n_842),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_905),
.B(n_848),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_916),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_905),
.A2(n_889),
.B(n_851),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_910),
.B(n_868),
.Y(n_944)
);

AO32x2_ASAP7_75t_L g945 ( 
.A1(n_910),
.A2(n_868),
.A3(n_876),
.B1(n_878),
.B2(n_885),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

NOR2x1_ASAP7_75t_SL g947 ( 
.A(n_918),
.B(n_851),
.Y(n_947)
);

AO21x2_ASAP7_75t_L g948 ( 
.A1(n_900),
.A2(n_866),
.B(n_859),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_912),
.B(n_848),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_917),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_912),
.A2(n_837),
.B(n_869),
.C(n_841),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_908),
.B(n_868),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_912),
.B(n_848),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_896),
.B(n_842),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_912),
.B(n_838),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_930),
.B(n_907),
.Y(n_956)
);

INVx8_ASAP7_75t_L g957 ( 
.A(n_929),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_896),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_929),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_929),
.A2(n_888),
.B(n_854),
.C(n_865),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_929),
.A2(n_856),
.B(n_847),
.C(n_849),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_908),
.A2(n_847),
.B(n_849),
.C(n_860),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_907),
.B(n_848),
.Y(n_963)
);

AOI21xp33_ASAP7_75t_L g964 ( 
.A1(n_907),
.A2(n_868),
.B(n_840),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_930),
.B(n_840),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_896),
.B(n_849),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_917),
.B(n_877),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_897),
.A2(n_847),
.B(n_872),
.C(n_870),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_900),
.A2(n_859),
.B(n_866),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_907),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_938),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_959),
.B(n_930),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_942),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_955),
.B(n_939),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_933),
.B(n_926),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_934),
.B(n_895),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_946),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_950),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_965),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_935),
.A2(n_915),
.B1(n_895),
.B2(n_873),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_943),
.A2(n_904),
.B1(n_877),
.B2(n_898),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_937),
.A2(n_904),
.B1(n_877),
.B2(n_898),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_958),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_947),
.B(n_896),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_944),
.B(n_895),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_969),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_940),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_933),
.B(n_926),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_969),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_967),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_967),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_952),
.B(n_926),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_956),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_952),
.B(n_898),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_948),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_977),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

OAI211xp5_ASAP7_75t_L g998 ( 
.A1(n_981),
.A2(n_951),
.B(n_960),
.C(n_968),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_984),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_977),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_976),
.B(n_898),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_977),
.Y(n_1002)
);

AND2x4_ASAP7_75t_SL g1003 ( 
.A(n_984),
.B(n_940),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_978),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_976),
.B(n_898),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_971),
.Y(n_1006)
);

OAI211xp5_ASAP7_75t_SL g1007 ( 
.A1(n_990),
.A2(n_991),
.B(n_982),
.C(n_974),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_990),
.Y(n_1008)
);

AOI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_980),
.A2(n_953),
.B1(n_957),
.B2(n_964),
.C(n_936),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_991),
.B(n_954),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_984),
.B(n_945),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_985),
.B(n_993),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_979),
.B(n_954),
.Y(n_1013)
);

NAND4xp25_ASAP7_75t_L g1014 ( 
.A(n_980),
.B(n_961),
.C(n_962),
.D(n_953),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_978),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_993),
.B(n_932),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_985),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_999),
.B(n_987),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_999),
.B(n_987),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_R g1020 ( 
.A(n_1011),
.B(n_970),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_996),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_997),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_996),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1010),
.B(n_979),
.Y(n_1024)
);

NAND2x1_ASAP7_75t_L g1025 ( 
.A(n_996),
.B(n_983),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1011),
.B(n_987),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1000),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_1018),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.B(n_1007),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1024),
.B(n_1008),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1022),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1023),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1017),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1029),
.B(n_1018),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1031),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1028),
.B(n_1026),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1035),
.B(n_1034),
.Y(n_1040)
);

OAI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_1038),
.A2(n_998),
.B1(n_1014),
.B2(n_1009),
.C(n_1020),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1036),
.A2(n_1019),
.B1(n_1026),
.B2(n_1033),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_1036),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_1035),
.B(n_1032),
.C(n_1033),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1037),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1035),
.B(n_1019),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_1035),
.A2(n_1025),
.B(n_936),
.C(n_957),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1035),
.B(n_1003),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_SL g1050 ( 
.A1(n_1041),
.A2(n_10),
.B(n_11),
.Y(n_1050)
);

OAI32xp33_ASAP7_75t_L g1051 ( 
.A1(n_1042),
.A2(n_1021),
.A3(n_1017),
.B1(n_997),
.B2(n_1006),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1047),
.A2(n_1021),
.B1(n_1003),
.B2(n_1006),
.Y(n_1052)
);

OAI221xp5_ASAP7_75t_SL g1053 ( 
.A1(n_1039),
.A2(n_1012),
.B1(n_995),
.B2(n_1005),
.C(n_1001),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1040),
.B(n_1027),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1044),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_1027),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1044),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1049),
.B(n_1016),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1045),
.B(n_1021),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1043),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1048),
.B(n_1013),
.Y(n_1062)
);

AOI222xp33_ASAP7_75t_L g1063 ( 
.A1(n_1041),
.A2(n_957),
.B1(n_995),
.B2(n_983),
.C1(n_941),
.C2(n_949),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1044),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.B(n_861),
.Y(n_1066)
);

AOI222xp33_ASAP7_75t_L g1067 ( 
.A1(n_1060),
.A2(n_983),
.B1(n_988),
.B2(n_975),
.C1(n_972),
.C2(n_992),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_1059),
.A2(n_10),
.B(n_13),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_1059),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1050),
.B(n_1015),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1057),
.B(n_1000),
.Y(n_1071)
);

XOR2x2_ASAP7_75t_L g1072 ( 
.A(n_1058),
.B(n_14),
.Y(n_1072)
);

XOR2x2_ASAP7_75t_L g1073 ( 
.A(n_1062),
.B(n_15),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_1064),
.B(n_15),
.C(n_16),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_1061),
.A2(n_988),
.B(n_975),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1054),
.B(n_1002),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1051),
.A2(n_1004),
.B(n_1002),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1056),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1063),
.B(n_1004),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1052),
.A2(n_1053),
.B1(n_1065),
.B2(n_1005),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1053),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1055),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1062),
.A2(n_963),
.B1(n_992),
.B2(n_966),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1055),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1084),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1073),
.A2(n_973),
.B(n_450),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1082),
.Y(n_1087)
);

OR3x1_ASAP7_75t_L g1088 ( 
.A(n_1068),
.B(n_964),
.C(n_973),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1072),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1069),
.B(n_1001),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_17),
.C(n_18),
.Y(n_1091)
);

NAND4xp25_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_994),
.C(n_972),
.D(n_450),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1066),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_1078),
.B(n_994),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1070),
.B(n_978),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1079),
.A2(n_904),
.B1(n_899),
.B2(n_894),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1074),
.B(n_17),
.Y(n_1097)
);

NAND4xp25_ASAP7_75t_L g1098 ( 
.A(n_1080),
.B(n_444),
.C(n_450),
.D(n_451),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1071),
.B(n_18),
.Y(n_1099)
);

OAI211xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1083),
.A2(n_415),
.B(n_419),
.C(n_428),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1075),
.B(n_20),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1089),
.A2(n_1076),
.B1(n_1077),
.B2(n_1067),
.C(n_25),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_L g1103 ( 
.A(n_1091),
.B(n_444),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1093),
.B(n_21),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1091),
.A2(n_915),
.B1(n_989),
.B2(n_986),
.C(n_444),
.Y(n_1105)
);

OAI322xp33_ASAP7_75t_L g1106 ( 
.A1(n_1085),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1097),
.A2(n_904),
.B1(n_986),
.B2(n_989),
.Y(n_1107)
);

NAND4xp25_ASAP7_75t_L g1108 ( 
.A(n_1090),
.B(n_444),
.C(n_450),
.D(n_451),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1094),
.B(n_1086),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1087),
.B(n_451),
.C(n_419),
.D(n_428),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1099),
.B(n_24),
.Y(n_1111)
);

OAI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1096),
.A2(n_915),
.B1(n_986),
.B2(n_989),
.C(n_451),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1092),
.B(n_30),
.Y(n_1113)
);

NAND4xp25_ASAP7_75t_L g1114 ( 
.A(n_1101),
.B(n_428),
.C(n_415),
.D(n_33),
.Y(n_1114)
);

AOI322xp5_ASAP7_75t_L g1115 ( 
.A1(n_1095),
.A2(n_899),
.A3(n_894),
.B1(n_945),
.B2(n_924),
.C1(n_904),
.C2(n_925),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1100),
.B(n_30),
.C(n_32),
.Y(n_1116)
);

NOR4xp25_ASAP7_75t_L g1117 ( 
.A(n_1098),
.B(n_34),
.C(n_35),
.D(n_36),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_1088),
.A2(n_36),
.B(n_37),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1089),
.A2(n_38),
.B(n_39),
.Y(n_1119)
);

AOI211xp5_ASAP7_75t_L g1120 ( 
.A1(n_1091),
.A2(n_39),
.B(n_40),
.C(n_42),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1089),
.A2(n_915),
.B1(n_894),
.B2(n_904),
.C(n_45),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1091),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1122)
);

AOI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1089),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1089),
.A2(n_46),
.B(n_47),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1093),
.Y(n_1125)
);

OAI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_1102),
.A2(n_899),
.B(n_904),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_1119),
.A2(n_48),
.B(n_50),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1125),
.Y(n_1128)
);

OAI22x1_ASAP7_75t_L g1129 ( 
.A1(n_1109),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1118),
.A2(n_459),
.B1(n_455),
.B2(n_454),
.C(n_904),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_1122),
.A2(n_459),
.B(n_455),
.Y(n_1131)
);

AOI222xp33_ASAP7_75t_L g1132 ( 
.A1(n_1123),
.A2(n_899),
.B1(n_454),
.B2(n_459),
.C1(n_455),
.C2(n_904),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1121),
.A2(n_904),
.B1(n_899),
.B2(n_917),
.Y(n_1133)
);

OAI211xp5_ASAP7_75t_L g1134 ( 
.A1(n_1117),
.A2(n_879),
.B(n_892),
.C(n_459),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1104),
.B(n_1120),
.C(n_1116),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_1124),
.A2(n_1106),
.B1(n_1105),
.B2(n_1114),
.C(n_1113),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1107),
.A2(n_925),
.B1(n_922),
.B2(n_919),
.Y(n_1137)
);

AOI211x1_ASAP7_75t_SL g1138 ( 
.A1(n_1111),
.A2(n_455),
.B(n_459),
.C(n_404),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1112),
.A2(n_922),
.B1(n_925),
.B2(n_919),
.Y(n_1139)
);

AOI222xp33_ASAP7_75t_L g1140 ( 
.A1(n_1103),
.A2(n_945),
.B1(n_919),
.B2(n_922),
.C1(n_914),
.C2(n_913),
.Y(n_1140)
);

AOI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1108),
.A2(n_53),
.B(n_54),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1115),
.B(n_924),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1110),
.A2(n_864),
.B(n_891),
.Y(n_1143)
);

OAI211xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1102),
.A2(n_886),
.B(n_404),
.C(n_59),
.Y(n_1144)
);

AOI222xp33_ASAP7_75t_L g1145 ( 
.A1(n_1102),
.A2(n_913),
.B1(n_914),
.B2(n_864),
.C1(n_902),
.C2(n_897),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1125),
.B(n_913),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1125),
.B(n_432),
.C(n_914),
.Y(n_1147)
);

NAND4xp25_ASAP7_75t_L g1148 ( 
.A(n_1102),
.B(n_902),
.C(n_927),
.D(n_60),
.Y(n_1148)
);

AOI221x1_ASAP7_75t_L g1149 ( 
.A1(n_1124),
.A2(n_432),
.B1(n_927),
.B2(n_906),
.C(n_920),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_1128),
.B(n_432),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1146),
.B(n_432),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1126),
.A2(n_902),
.B1(n_931),
.B2(n_918),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1135),
.B(n_918),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1127),
.B(n_57),
.Y(n_1154)
);

OAI31xp33_ASAP7_75t_L g1155 ( 
.A1(n_1134),
.A2(n_902),
.A3(n_927),
.B(n_62),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1129),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1147),
.Y(n_1157)
);

NAND4xp75_ASAP7_75t_L g1158 ( 
.A(n_1130),
.B(n_931),
.C(n_61),
.D(n_68),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1138),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1148),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1136),
.A2(n_1144),
.B1(n_1133),
.B2(n_1145),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1142),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1149),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1139),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_1131),
.B(n_432),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1132),
.B(n_58),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_L g1167 ( 
.A(n_1141),
.B(n_432),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1137),
.B(n_902),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1143),
.B(n_70),
.Y(n_1169)
);

NOR4xp75_ASAP7_75t_L g1170 ( 
.A(n_1140),
.B(n_71),
.C(n_72),
.D(n_74),
.Y(n_1170)
);

OA22x2_ASAP7_75t_L g1171 ( 
.A1(n_1129),
.A2(n_918),
.B1(n_897),
.B2(n_901),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1156),
.B(n_75),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1162),
.A2(n_902),
.B1(n_909),
.B2(n_911),
.C(n_920),
.Y(n_1173)
);

NAND4xp25_ASAP7_75t_L g1174 ( 
.A(n_1161),
.B(n_78),
.C(n_79),
.D(n_82),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1150),
.Y(n_1175)
);

NAND4xp75_ASAP7_75t_L g1176 ( 
.A(n_1167),
.B(n_83),
.C(n_95),
.D(n_97),
.Y(n_1176)
);

AOI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_1151),
.B1(n_1160),
.B2(n_1157),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1171),
.A2(n_900),
.B(n_918),
.Y(n_1178)
);

NOR2x1p5_ASAP7_75t_L g1179 ( 
.A(n_1164),
.B(n_101),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1154),
.A2(n_1169),
.B(n_1166),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1159),
.B(n_1153),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1165),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1153),
.A2(n_902),
.B1(n_918),
.B2(n_948),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1170),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1155),
.A2(n_102),
.B(n_103),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1158),
.Y(n_1186)
);

AOI322xp5_ASAP7_75t_L g1187 ( 
.A1(n_1152),
.A2(n_920),
.A3(n_901),
.B1(n_903),
.B2(n_906),
.C1(n_921),
.C2(n_928),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_1181),
.B(n_1168),
.C(n_106),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1176),
.B(n_1179),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1172),
.Y(n_1190)
);

AOI322xp5_ASAP7_75t_L g1191 ( 
.A1(n_1184),
.A2(n_920),
.A3(n_901),
.B1(n_903),
.B2(n_906),
.C1(n_928),
.C2(n_921),
.Y(n_1191)
);

OAI211xp5_ASAP7_75t_L g1192 ( 
.A1(n_1177),
.A2(n_104),
.B(n_108),
.C(n_111),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1175),
.B(n_1186),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1182),
.Y(n_1194)
);

NOR3x1_ASAP7_75t_L g1195 ( 
.A(n_1174),
.B(n_114),
.C(n_128),
.Y(n_1195)
);

OAI211xp5_ASAP7_75t_SL g1196 ( 
.A1(n_1180),
.A2(n_129),
.B(n_130),
.C(n_132),
.Y(n_1196)
);

OA22x2_ASAP7_75t_L g1197 ( 
.A1(n_1185),
.A2(n_1178),
.B1(n_1173),
.B2(n_1183),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1187),
.A2(n_918),
.B1(n_901),
.B2(n_903),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1179),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1175),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1181),
.A2(n_911),
.B1(n_909),
.B2(n_139),
.C(n_141),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1184),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1194),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1202),
.A2(n_918),
.B1(n_906),
.B2(n_903),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1200),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1200),
.Y(n_1206)
);

AOI31xp33_ASAP7_75t_L g1207 ( 
.A1(n_1189),
.A2(n_136),
.A3(n_137),
.B(n_144),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1199),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1190),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1188),
.A2(n_918),
.B1(n_921),
.B2(n_928),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1193),
.A2(n_928),
.B1(n_921),
.B2(n_911),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1197),
.A2(n_1201),
.B1(n_1196),
.B2(n_1198),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1205),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1208),
.A2(n_1192),
.B1(n_1195),
.B2(n_1191),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1203),
.A2(n_1206),
.B1(n_1212),
.B2(n_1209),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1210),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1207),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_911),
.B1(n_909),
.B2(n_846),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1217),
.A2(n_1204),
.B1(n_151),
.B2(n_153),
.Y(n_1219)
);

AOI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1213),
.A2(n_146),
.B1(n_154),
.B2(n_155),
.Y(n_1220)
);

OAI22x1_ASAP7_75t_L g1221 ( 
.A1(n_1214),
.A2(n_156),
.B1(n_160),
.B2(n_168),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1215),
.B(n_169),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1216),
.B1(n_1218),
.B2(n_911),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1223),
.B(n_1219),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1224),
.B(n_1221),
.Y(n_1225)
);

XNOR2xp5_ASAP7_75t_L g1226 ( 
.A(n_1225),
.B(n_1220),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_170),
.B1(n_174),
.B2(n_176),
.C(n_177),
.Y(n_1227)
);

AOI211xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_178),
.B(n_179),
.C(n_181),
.Y(n_1228)
);


endmodule