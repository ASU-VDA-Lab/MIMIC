module fake_netlist_1_8888_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_38;
wire n_20;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_8), .B(n_4), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_9), .B(n_12), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_3), .B(n_7), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_10), .B(n_3), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_17), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g25 ( .A(n_17), .B(n_5), .C(n_1), .Y(n_25) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_21), .B(n_0), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_24), .B(n_15), .Y(n_27) );
OAI21x1_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_19), .B(n_15), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_16), .B(n_22), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_31), .B(n_29), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_26), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
O2A1O1Ixp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_36), .B(n_34), .C(n_30), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
AOI31xp33_ASAP7_75t_R g39 ( .A1(n_36), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_39) );
CKINVDCx16_ASAP7_75t_R g40 ( .A(n_39), .Y(n_40) );
NOR2x1_ASAP7_75t_L g41 ( .A(n_37), .B(n_25), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_38), .Y(n_42) );
AOI21xp5_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_16), .B(n_20), .Y(n_43) );
HB1xp67_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_44), .Y(n_45) );
AOI22x1_ASAP7_75t_L g46 ( .A1(n_45), .A2(n_40), .B1(n_43), .B2(n_2), .Y(n_46) );
endmodule