module real_jpeg_21683_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_67;
wire n_58;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_61;
wire n_25;
wire n_71;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_39;
wire n_36;
wire n_40;
wire n_70;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_6),
.B1(n_15),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_6),
.B(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_20),
.B1(n_44),
.B2(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_2),
.A2(n_6),
.B1(n_15),
.B2(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_18),
.B1(n_30),
.B2(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_6),
.B1(n_15),
.B2(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_15),
.Y(n_14)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_5),
.A2(n_6),
.B1(n_15),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_8),
.B1(n_15),
.B2(n_28),
.Y(n_36)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_53),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_40),
.B(n_52),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_24),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_22),
.A2(n_45),
.B(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_26),
.B(n_32),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_36),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_30),
.A2(n_31),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_51),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_73),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);


endmodule