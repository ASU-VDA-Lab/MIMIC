module real_jpeg_27558_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_0),
.A2(n_32),
.B1(n_40),
.B2(n_41),
.Y(n_86)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_42),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_67),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_9),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_62),
.B(n_63),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_40),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_9),
.A2(n_40),
.B(n_44),
.C(n_179),
.D(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_72),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_25),
.B(n_192),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_9),
.A2(n_64),
.B(n_75),
.C(n_111),
.D(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_9),
.B(n_64),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_56),
.Y(n_199)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_80),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_80),
.Y(n_194)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_26),
.B1(n_33),
.B2(n_50),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_130)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_21),
.B(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_87),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_22),
.B(n_81),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_23),
.B(n_54),
.C(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_24),
.B(n_38),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_25),
.A2(n_34),
.B1(n_36),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_25),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_34),
.B(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_25),
.A2(n_34),
.B1(n_104),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_25),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_25),
.B(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_26),
.B(n_45),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_29),
.B(n_98),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_35),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g178 ( 
.A1(n_33),
.A2(n_41),
.A3(n_46),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_33),
.B(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_34),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_34),
.A2(n_199),
.B(n_207),
.Y(n_206)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_35),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_39),
.A2(n_51),
.B(n_145),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_45),
.Y(n_47)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_40),
.A2(n_63),
.A3(n_221),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_41),
.B(n_230),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_43),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_44),
.A2(n_48),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_44),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_44),
.A2(n_48),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_51),
.B(n_147),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_51),
.A2(n_145),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_51),
.B(n_98),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_61),
.B(n_98),
.C(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_59),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_60),
.B(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_66),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_74),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_71),
.B1(n_107),
.B2(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_79),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_71),
.A2(n_74),
.B(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_72),
.A2(n_75),
.B1(n_109),
.B2(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_87),
.A2(n_88),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.C(n_105),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_90),
.B1(n_105),
.B2(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_93),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_92),
.B(n_98),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_102),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_132),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_131),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_171),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_157),
.B(n_170),
.Y(n_136)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_137),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_154),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_142),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_151),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_144),
.B1(n_151),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_160),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_164),
.B(n_165),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_166),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_167),
.B(n_169),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_249),
.C(n_250),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_244),
.B(n_248),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_233),
.B(n_243),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_216),
.B(n_232),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_195),
.B(n_215),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_177),
.B(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_181),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_203),
.B(n_214),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_208),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_209),
.B(n_213),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.C(n_225),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_228),
.Y(n_239)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);


endmodule