module fake_netlist_6_3615_n_1911 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1911);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1911;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_14),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_36),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_39),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_7),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_68),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_95),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_16),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_81),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_94),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_80),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_64),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_147),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_0),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_164),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_132),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_117),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_8),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_91),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_99),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_30),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_98),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_158),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_152),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_39),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_88),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_93),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_30),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_46),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_57),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_38),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_71),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_162),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_62),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_21),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_35),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_150),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_160),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_59),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_89),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_27),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_11),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_115),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_63),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_122),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_62),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_107),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_124),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_112),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_3),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_177),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_109),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_46),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_114),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_47),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_135),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_79),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_66),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_108),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_14),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_21),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_22),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_100),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_33),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_103),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_144),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_87),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_44),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_163),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_137),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_179),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_16),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_26),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_82),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_70),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_37),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_170),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_58),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_37),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_136),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_0),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_63),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_41),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_102),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_8),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_51),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_138),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_42),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_118),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_73),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_60),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_18),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_123),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_174),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_52),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_17),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_140),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_13),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_49),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_104),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_53),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_86),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_165),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_56),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_33),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_181),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_47),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_120),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_64),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_55),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_41),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_29),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_119),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_111),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_74),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_146),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_2),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_175),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_19),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_154),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_166),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_51),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_11),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_131),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_105),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_72),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_50),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_19),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_189),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_9),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_44),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_34),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_101),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_31),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_153),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_130),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_141),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_43),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_157),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_67),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_52),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_182),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_23),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_106),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_6),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_186),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_43),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_205),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_255),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_332),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_234),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_255),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_247),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_247),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_238),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_239),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_280),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_203),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_209),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_240),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_230),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_254),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_199),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_199),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_193),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_242),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_256),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_262),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_219),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_261),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_263),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_268),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_274),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_266),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_244),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_276),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_279),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_288),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_230),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_270),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_377),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_306),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_196),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_219),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_314),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_199),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_192),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_230),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_322),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_272),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_329),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_340),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_192),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_194),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_345),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_282),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_284),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_287),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_363),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_372),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_246),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_260),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_257),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_257),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_195),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_210),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_220),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_248),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_222),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_250),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_227),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_297),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_230),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_230),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_245),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_253),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_211),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_211),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_215),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_271),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_215),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_298),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_217),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_230),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_258),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_217),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_251),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_267),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_310),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_265),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_251),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_391),
.B(n_294),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_251),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_401),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_438),
.B(n_294),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_267),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_437),
.A2(n_223),
.B1(n_194),
.B2(n_201),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_321),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_391),
.B(n_294),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_243),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_389),
.A2(n_300),
.B1(n_291),
.B2(n_346),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_482),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_402),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_410),
.A2(n_320),
.B1(n_317),
.B2(n_319),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_405),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_484),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_423),
.B(n_321),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_484),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_423),
.B(n_334),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_487),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_201),
.Y(n_526)
);

BUFx8_ASAP7_75t_L g527 ( 
.A(n_398),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_R g528 ( 
.A(n_414),
.B(n_197),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_409),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_406),
.B(n_334),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_416),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_435),
.B(n_465),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_419),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_468),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_415),
.B(n_307),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_470),
.B(n_383),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_392),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_420),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_472),
.B(n_383),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_476),
.B(n_273),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_424),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_R g556 ( 
.A(n_395),
.B(n_429),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_422),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_415),
.B(n_307),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_422),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_460),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_477),
.B(n_277),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_398),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_491),
.B(n_290),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_475),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_390),
.B(n_307),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_425),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_469),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_485),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_535),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_506),
.B(n_417),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_538),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_500),
.B(n_280),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_539),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_539),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_496),
.B(n_280),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_511),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_544),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_544),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_481),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_498),
.B(n_418),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_552),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_498),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_510),
.B(n_428),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_500),
.B(n_393),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_511),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_534),
.B(n_252),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_538),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_540),
.B(n_428),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_526),
.B(n_471),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_500),
.B(n_394),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_552),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_559),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_434),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_521),
.A2(n_304),
.B(n_292),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_500),
.A2(n_448),
.B1(n_449),
.B2(n_441),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_516),
.B(n_462),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_538),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_496),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_524),
.A2(n_315),
.B(n_309),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_557),
.B(n_463),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_496),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_538),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_494),
.B(n_486),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_538),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_543),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_560),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_560),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_496),
.A2(n_554),
.B1(n_502),
.B2(n_546),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_543),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_566),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_571),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_571),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_571),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_554),
.A2(n_431),
.B1(n_436),
.B2(n_432),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_574),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_511),
.Y(n_635)
);

AO21x2_ASAP7_75t_L g636 ( 
.A1(n_550),
.A2(n_335),
.B(n_328),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_527),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_557),
.B(n_434),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_512),
.A2(n_368),
.B1(n_339),
.B2(n_257),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_574),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_R g643 ( 
.A(n_556),
.B(n_445),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_SL g644 ( 
.A(n_528),
.B(n_445),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_545),
.B(n_451),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_505),
.A2(n_249),
.B1(n_324),
.B2(n_323),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_545),
.A2(n_382),
.B1(n_233),
.B2(n_229),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_451),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_568),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_507),
.A2(n_364),
.B1(n_302),
.B2(n_382),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_543),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_558),
.B(n_453),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_511),
.Y(n_655)
);

AO22x2_ASAP7_75t_L g656 ( 
.A1(n_558),
.A2(n_347),
.B1(n_381),
.B2(n_362),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_527),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_542),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_554),
.B(n_542),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_511),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_554),
.B(n_230),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_511),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_517),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_542),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_520),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_567),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_567),
.B(n_453),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_514),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_517),
.Y(n_671)
);

AND3x2_ASAP7_75t_L g672 ( 
.A(n_514),
.B(n_305),
.C(n_440),
.Y(n_672)
);

INVxp33_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_533),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_454),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_527),
.B(n_454),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_520),
.B(n_473),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_519),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_519),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_564),
.B(n_473),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_565),
.B(n_490),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_493),
.B(n_396),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_523),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_564),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_493),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_520),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_497),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_520),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_564),
.B(n_483),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_564),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_548),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_546),
.B(n_483),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_495),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_495),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_499),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_546),
.B(n_490),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_537),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_541),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_499),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_541),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_503),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_504),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_504),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_508),
.B(n_269),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_547),
.A2(n_360),
.B1(n_233),
.B2(n_229),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_546),
.B(n_293),
.Y(n_713)
);

AND3x2_ASAP7_75t_L g714 ( 
.A(n_547),
.B(n_361),
.C(n_341),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_508),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_551),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_509),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_555),
.A2(n_464),
.B1(n_439),
.B2(n_443),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_555),
.Y(n_720)
);

OAI21xp33_ASAP7_75t_SL g721 ( 
.A1(n_569),
.A2(n_427),
.B(n_426),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_569),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_509),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_570),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_611),
.B(n_513),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_592),
.B(n_570),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_611),
.A2(n_230),
.B1(n_380),
.B2(n_303),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_598),
.B(n_336),
.C(n_326),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_615),
.A2(n_518),
.B(n_513),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_615),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_675),
.B(n_515),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_690),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_690),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_581),
.B(n_518),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_674),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_592),
.B(n_531),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_639),
.B(n_573),
.C(n_549),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_301),
.B1(n_259),
.B2(n_264),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_576),
.B(n_562),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_581),
.B(n_522),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_593),
.B(n_197),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_581),
.B(n_522),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_650),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_620),
.A2(n_529),
.B(n_525),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_623),
.B(n_717),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_618),
.B(n_600),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_589),
.B(n_206),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_717),
.B(n_525),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_665),
.A2(n_280),
.B1(n_380),
.B2(n_303),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_706),
.B(n_529),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_699),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_667),
.B(n_280),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_658),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_706),
.B(n_665),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_659),
.A2(n_572),
.B(n_532),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_706),
.B(n_530),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_658),
.B(n_572),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_644),
.A2(n_275),
.B1(n_278),
.B2(n_281),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_532),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_594),
.A2(n_325),
.B1(n_283),
.B2(n_285),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_721),
.A2(n_450),
.B(n_444),
.C(n_446),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_687),
.B(n_286),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_658),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_697),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_702),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_643),
.B(n_198),
.Y(n_767)
);

INVx8_ASAP7_75t_L g768 ( 
.A(n_584),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_699),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_687),
.B(n_289),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_584),
.B(n_303),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_607),
.B(n_348),
.C(n_337),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_604),
.B(n_198),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_691),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_636),
.A2(n_303),
.B1(n_380),
.B2(n_447),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_703),
.B(n_295),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_704),
.B(n_705),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_704),
.B(n_296),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_L g779 ( 
.A(n_682),
.B(n_353),
.C(n_352),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_669),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_636),
.A2(n_380),
.B1(n_456),
.B2(n_455),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_699),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_670),
.B(n_380),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_594),
.A2(n_330),
.B1(n_299),
.B2(n_312),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_601),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_700),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_707),
.B(n_313),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_670),
.B(n_318),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_707),
.B(n_716),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_720),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_669),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_636),
.A2(n_452),
.B1(n_206),
.B2(n_360),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_670),
.B(n_331),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_700),
.Y(n_794)
);

BUFx6f_ASAP7_75t_SL g795 ( 
.A(n_596),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_661),
.B(n_338),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_700),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_722),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_601),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_722),
.B(n_724),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_636),
.A2(n_369),
.B1(n_216),
.B2(n_223),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_590),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_701),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_701),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_692),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_671),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_683),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_721),
.A2(n_459),
.B(n_458),
.C(n_457),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_708),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_711),
.B(n_343),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_708),
.B(n_710),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_708),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_589),
.B(n_426),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_710),
.B(n_344),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_710),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_683),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_664),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_715),
.B(n_349),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_715),
.Y(n_820)
);

NOR2x1p5_ASAP7_75t_L g821 ( 
.A(n_693),
.B(n_214),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_715),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_718),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_709),
.A2(n_459),
.B(n_458),
.C(n_457),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_718),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_614),
.B(n_430),
.C(n_427),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_661),
.B(n_355),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_673),
.B(n_339),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_584),
.A2(n_375),
.B1(n_214),
.B2(n_216),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_723),
.B(n_356),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_723),
.B(n_713),
.Y(n_831)
);

NAND2x1_ASAP7_75t_L g832 ( 
.A(n_692),
.B(n_397),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_SL g833 ( 
.A1(n_596),
.A2(n_237),
.B1(n_302),
.B2(n_364),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_612),
.B(n_430),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_647),
.B(n_357),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_692),
.B(n_359),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_577),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_671),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_577),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_577),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_578),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_694),
.B(n_200),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_578),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_578),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_200),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_648),
.B(n_339),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_678),
.B(n_202),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_671),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_580),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_580),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_694),
.B(n_202),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_580),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_596),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_638),
.B(n_358),
.C(n_237),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_680),
.B(n_204),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_663),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_663),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_663),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_653),
.B(n_207),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_653),
.B(n_207),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_596),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_645),
.B(n_208),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_579),
.B(n_212),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_654),
.B(n_212),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_677),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_579),
.B(n_213),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_579),
.B(n_213),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_579),
.B(n_218),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_583),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_596),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_677),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_656),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_668),
.B(n_218),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_583),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_698),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_684),
.B(n_221),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_652),
.B(n_369),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_684),
.B(n_221),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_583),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_684),
.B(n_224),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_656),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_791),
.B(n_696),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_754),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_732),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_806),
.B(n_656),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_754),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_881),
.A2(n_656),
.B1(n_584),
.B2(n_648),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_881),
.A2(n_656),
.B1(n_584),
.B2(n_712),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_823),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_823),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_846),
.A2(n_637),
.B1(n_657),
.B2(n_688),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_799),
.B(n_597),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_747),
.A2(n_608),
.B(n_631),
.C(n_712),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_732),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_758),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_780),
.B(n_828),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_744),
.B(n_676),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_873),
.B(n_652),
.C(n_672),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_766),
.A2(n_584),
.B1(n_681),
.B2(n_695),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_612),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_746),
.A2(n_875),
.B1(n_730),
.B2(n_758),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_733),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_735),
.A2(n_637),
.B1(n_657),
.B2(n_688),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_777),
.A2(n_373),
.B(n_375),
.C(n_719),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_734),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_754),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_742),
.B(n_597),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_764),
.B(n_714),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_SL g909 ( 
.A(n_731),
.B(n_373),
.C(n_225),
.Y(n_909)
);

AO22x1_ASAP7_75t_L g910 ( 
.A1(n_854),
.A2(n_367),
.B1(n_224),
.B2(n_225),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_734),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_773),
.B(n_610),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_736),
.B(n_610),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_774),
.B(n_610),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_765),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_814),
.B(n_397),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_752),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_764),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_790),
.B(n_610),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_798),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_831),
.B(n_616),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_741),
.B(n_616),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_765),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_789),
.B(n_616),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_768),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_802),
.B(n_686),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_752),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_818),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_769),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_737),
.B(n_399),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_800),
.B(n_616),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_811),
.B(n_619),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_807),
.A2(n_633),
.B(n_666),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_743),
.B(n_619),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_872),
.A2(n_584),
.B1(n_624),
.B2(n_575),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_769),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_756),
.B(n_619),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_749),
.B(n_619),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_725),
.B(n_625),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_808),
.B(n_399),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_782),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_817),
.B(n_625),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_775),
.A2(n_591),
.B1(n_642),
.B2(n_609),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_834),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_760),
.B(n_807),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_R g946 ( 
.A(n_740),
.B(n_606),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_782),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_877),
.B(n_726),
.Y(n_948)
);

AND2x4_ASAP7_75t_SL g949 ( 
.A(n_834),
.B(n_684),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_853),
.A2(n_641),
.B1(n_632),
.B2(n_625),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_853),
.B(n_606),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_807),
.B(n_632),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_755),
.B(n_632),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_861),
.B(n_786),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_812),
.A2(n_641),
.B(n_582),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_726),
.B(n_686),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_726),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_861),
.B(n_641),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_726),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_748),
.Y(n_960)
);

INVxp67_ASAP7_75t_SL g961 ( 
.A(n_838),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_834),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_824),
.A2(n_622),
.B(n_575),
.C(n_582),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_786),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_838),
.B(n_641),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_767),
.B(n_400),
.Y(n_966)
);

BUFx8_ASAP7_75t_L g967 ( 
.A(n_795),
.Y(n_967)
);

OR2x6_ASAP7_75t_SL g968 ( 
.A(n_772),
.B(n_226),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_870),
.B(n_686),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_862),
.B(n_633),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_794),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_768),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_797),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_797),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_803),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_834),
.B(n_400),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_803),
.Y(n_977)
);

INVx5_ASAP7_75t_L g978 ( 
.A(n_768),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_848),
.B(n_609),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_767),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_848),
.B(n_622),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_804),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_804),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_821),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_842),
.A2(n_689),
.B1(n_685),
.B2(n_679),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_832),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_805),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_845),
.B(n_624),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_805),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_810),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_851),
.B(n_629),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_810),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_809),
.A2(n_629),
.B(n_642),
.C(n_407),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_820),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_862),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_763),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_813),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_864),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_864),
.B(n_788),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_795),
.B(n_613),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_795),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_816),
.B(n_684),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_770),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_826),
.B(n_779),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_751),
.B(n_587),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_822),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_L g1007 ( 
.A1(n_753),
.A2(n_613),
.B(n_685),
.C(n_679),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_792),
.B(n_633),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_837),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_825),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_757),
.B(n_587),
.Y(n_1011)
);

BUFx8_ASAP7_75t_L g1012 ( 
.A(n_833),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_836),
.B(n_633),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_837),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_839),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_839),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_835),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_840),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_776),
.B(n_588),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_778),
.B(n_588),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_L g1021 ( 
.A(n_863),
.B(n_866),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_729),
.B(n_646),
.Y(n_1022)
);

OR2x4_ASAP7_75t_L g1023 ( 
.A(n_787),
.B(n_403),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_840),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_728),
.B(n_655),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_841),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_762),
.B(n_655),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_847),
.B(n_599),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_843),
.B(n_646),
.Y(n_1029)
);

NOR2x2_ASAP7_75t_L g1030 ( 
.A(n_801),
.B(n_835),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_843),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_847),
.B(n_599),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_781),
.A2(n_634),
.B1(n_599),
.B2(n_602),
.Y(n_1033)
);

BUFx8_ASAP7_75t_SL g1034 ( 
.A(n_738),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_844),
.B(n_849),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_844),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_829),
.B(n_403),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_796),
.B(n_602),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_859),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_849),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_867),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_850),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_759),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_852),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_856),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_852),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_869),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_739),
.B(n_677),
.Y(n_1048)
);

BUFx4f_ASAP7_75t_L g1049 ( 
.A(n_857),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_860),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_1043),
.B(n_762),
.C(n_824),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_920),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_961),
.B(n_874),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1013),
.A2(n_793),
.B(n_788),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_897),
.B(n_761),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_893),
.A2(n_796),
.B(n_827),
.C(n_793),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_928),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_896),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_1003),
.B(n_784),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_1013),
.A2(n_753),
.B(n_880),
.C(n_878),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_945),
.A2(n_771),
.B(n_783),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_893),
.A2(n_860),
.B(n_827),
.C(n_878),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_928),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_930),
.B(n_783),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_897),
.B(n_855),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1017),
.A2(n_880),
.B(n_876),
.C(n_868),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1003),
.B(n_815),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_926),
.B(n_819),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_926),
.B(n_830),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_948),
.A2(n_876),
.B1(n_745),
.B2(n_374),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_937),
.A2(n_871),
.B(n_865),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_909),
.A2(n_771),
.B(n_858),
.C(n_874),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_898),
.B(n_226),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1041),
.B(n_879),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_879),
.B(n_685),
.C(n_689),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_925),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_996),
.B(n_228),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1050),
.A2(n_727),
.B(n_750),
.C(n_689),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_SL g1080 ( 
.A1(n_923),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_998),
.B(n_231),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_948),
.A2(n_235),
.B1(n_232),
.B2(n_236),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_927),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1021),
.A2(n_666),
.B(n_586),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_956),
.B(n_235),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_956),
.B(n_236),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_883),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1050),
.A2(n_662),
.B(n_655),
.C(n_651),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_916),
.B(n_603),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_995),
.B(n_980),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_915),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_966),
.Y(n_1092)
);

OAI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_999),
.A2(n_308),
.B1(n_378),
.B2(n_365),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_SL g1094 ( 
.A(n_891),
.B(n_370),
.C(n_367),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_932),
.A2(n_666),
.B(n_586),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1039),
.B(n_603),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_1001),
.B(n_308),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1039),
.A2(n_662),
.B(n_649),
.C(n_651),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_968),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_999),
.A2(n_365),
.B1(n_387),
.B2(n_366),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_984),
.B(n_366),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_976),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_999),
.A2(n_370),
.B1(n_385),
.B2(n_374),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1004),
.B(n_376),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_887),
.A2(n_376),
.B1(n_378),
.B2(n_385),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_970),
.A2(n_662),
.B(n_627),
.C(n_605),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_957),
.A2(n_651),
.B(n_649),
.C(n_626),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_887),
.A2(n_387),
.B1(n_404),
.B2(n_407),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_929),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_901),
.B(n_617),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_R g1111 ( 
.A(n_946),
.B(n_75),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1034),
.Y(n_1112)
);

HAxp5_ASAP7_75t_L g1113 ( 
.A(n_1012),
.B(n_1034),
.CON(n_1113),
.SN(n_1113)
);

XOR2xp5_ASAP7_75t_L g1114 ( 
.A(n_899),
.B(n_76),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_940),
.B(n_404),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_918),
.B(n_621),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_957),
.A2(n_627),
.B(n_634),
.C(n_621),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_889),
.B(n_621),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_890),
.B(n_626),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_900),
.B(n_666),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_978),
.A2(n_586),
.B(n_585),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_903),
.A2(n_628),
.B(n_634),
.C(n_626),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_960),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_976),
.A2(n_413),
.B1(n_412),
.B2(n_5),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_910),
.B(n_412),
.C(n_413),
.Y(n_1125)
);

NOR3xp33_ASAP7_75t_SL g1126 ( 
.A(n_969),
.B(n_2),
.C(n_4),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_883),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1023),
.B(n_660),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_993),
.A2(n_640),
.B(n_630),
.C(n_628),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1023),
.B(n_660),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_888),
.A2(n_627),
.B1(n_640),
.B2(n_630),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_891),
.A2(n_5),
.B1(n_12),
.B2(n_15),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_941),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_886),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_978),
.A2(n_586),
.B(n_635),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_895),
.A2(n_630),
.B1(n_635),
.B2(n_660),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_959),
.B(n_660),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_944),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1048),
.A2(n_660),
.B(n_635),
.C(n_595),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_947),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_884),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_978),
.A2(n_635),
.B(n_595),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_993),
.A2(n_12),
.B(n_15),
.C(n_17),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_962),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_937),
.A2(n_991),
.B(n_988),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1030),
.Y(n_1146)
);

OR2x6_ASAP7_75t_SL g1147 ( 
.A(n_942),
.B(n_20),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_976),
.B(n_635),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_L g1149 ( 
.A1(n_907),
.A2(n_595),
.B(n_585),
.C(n_184),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_912),
.A2(n_595),
.B(n_585),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_882),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_921),
.B(n_595),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1045),
.B(n_585),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_924),
.B(n_585),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_908),
.Y(n_1155)
);

AO32x2_ASAP7_75t_L g1156 ( 
.A1(n_985),
.A2(n_20),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1008),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_964),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_885),
.A2(n_25),
.B(n_28),
.C(n_29),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_922),
.A2(n_77),
.B(n_178),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1045),
.A2(n_28),
.B(n_31),
.C(n_32),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1037),
.A2(n_32),
.B(n_34),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1049),
.B(n_156),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1019),
.A2(n_155),
.B(n_149),
.Y(n_1164)
);

AO22x2_ASAP7_75t_L g1165 ( 
.A1(n_1027),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1020),
.A2(n_145),
.B(n_128),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_922),
.A2(n_127),
.B(n_125),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1049),
.B(n_121),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1025),
.A2(n_116),
.B1(n_96),
.B2(n_84),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_967),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_946),
.B(n_40),
.Y(n_1171)
);

AO21x1_ASAP7_75t_L g1172 ( 
.A1(n_954),
.A2(n_934),
.B(n_1032),
.Y(n_1172)
);

INVx6_ASAP7_75t_L g1173 ( 
.A(n_886),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_906),
.B(n_45),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_973),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_906),
.B(n_48),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_906),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_974),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_975),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_994),
.B(n_1006),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1060),
.B(n_931),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1057),
.A2(n_1007),
.B(n_955),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1139),
.A2(n_1172),
.A3(n_1067),
.B(n_1088),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1053),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1058),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1072),
.A2(n_1007),
.B(n_1022),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1063),
.A2(n_972),
.B(n_925),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_SL g1188 ( 
.A1(n_1167),
.A2(n_1028),
.B(n_888),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1064),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1055),
.A2(n_1038),
.A3(n_939),
.B(n_938),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1051),
.A2(n_1008),
.B(n_1025),
.C(n_963),
.Y(n_1191)
);

NAND3x1_ASAP7_75t_L g1192 ( 
.A(n_1103),
.B(n_1012),
.C(n_950),
.Y(n_1192)
);

AND3x2_ASAP7_75t_L g1193 ( 
.A(n_1092),
.B(n_908),
.C(n_1027),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1146),
.A2(n_949),
.B1(n_958),
.B2(n_1006),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1138),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1150),
.A2(n_1022),
.B(n_953),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1145),
.A2(n_1005),
.B(n_1011),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1069),
.A2(n_1010),
.B(n_914),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1059),
.B(n_994),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1157),
.A2(n_935),
.B1(n_943),
.B2(n_949),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1115),
.B(n_905),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1141),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1112),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1066),
.B(n_1089),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1106),
.A2(n_1129),
.B(n_1142),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1077),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1075),
.B(n_935),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1098),
.A2(n_982),
.A3(n_997),
.B(n_990),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1068),
.B(n_911),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1180),
.B(n_971),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1076),
.A2(n_1002),
.B(n_952),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1061),
.A2(n_1035),
.B(n_981),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1121),
.A2(n_965),
.B(n_933),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1062),
.A2(n_979),
.B(n_1029),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1083),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1149),
.A2(n_1152),
.B(n_1154),
.Y(n_1217)
);

AOI211x1_ASAP7_75t_L g1218 ( 
.A1(n_1162),
.A2(n_892),
.B(n_913),
.C(n_919),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1109),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1077),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1087),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_1130),
.B(n_1128),
.C(n_1071),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1152),
.A2(n_943),
.B(n_1033),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1154),
.A2(n_1033),
.B(n_987),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1110),
.A2(n_1047),
.B(n_1015),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_1090),
.Y(n_1226)
);

AOI221x1_ASAP7_75t_L g1227 ( 
.A1(n_1165),
.A2(n_1044),
.B1(n_1018),
.B2(n_1014),
.C(n_1026),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1133),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1094),
.A2(n_1000),
.B1(n_986),
.B2(n_1009),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1126),
.B(n_1100),
.C(n_1082),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1114),
.A2(n_983),
.B1(n_977),
.B2(n_989),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1081),
.B(n_894),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1155),
.B(n_992),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1084),
.A2(n_1054),
.B(n_1095),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1165),
.A2(n_1046),
.B1(n_1009),
.B2(n_1036),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1144),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1123),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1159),
.A2(n_936),
.B(n_917),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1170),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1153),
.A2(n_1026),
.B(n_902),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1087),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1122),
.A2(n_1042),
.B(n_1040),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1104),
.B(n_1031),
.Y(n_1243)
);

AO32x2_ASAP7_75t_L g1244 ( 
.A1(n_1132),
.A2(n_951),
.A3(n_1000),
.B1(n_1024),
.B2(n_1016),
.Y(n_1244)
);

OA22x2_ASAP7_75t_L g1245 ( 
.A1(n_1080),
.A2(n_1046),
.B1(n_55),
.B2(n_57),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1135),
.A2(n_951),
.B(n_1026),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1171),
.B(n_61),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1165),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_1248)
);

OA22x2_ASAP7_75t_L g1249 ( 
.A1(n_1102),
.A2(n_60),
.B1(n_1078),
.B2(n_1105),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1096),
.A2(n_1164),
.B(n_1166),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1107),
.A2(n_1117),
.B(n_1160),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1087),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1140),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1073),
.A2(n_1079),
.B(n_1131),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1158),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1116),
.A2(n_1118),
.B(n_1119),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1175),
.B(n_1179),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1077),
.A2(n_1120),
.B(n_1163),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1091),
.B(n_1151),
.Y(n_1259)
);

AOI31xp67_ASAP7_75t_L g1260 ( 
.A1(n_1136),
.A2(n_1169),
.A3(n_1168),
.B(n_1137),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1085),
.B(n_1086),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1178),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1093),
.B(n_1148),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1097),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1077),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1127),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1147),
.Y(n_1267)
);

AO32x2_ASAP7_75t_L g1268 ( 
.A1(n_1108),
.A2(n_1105),
.A3(n_1156),
.B1(n_1052),
.B2(n_1177),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1162),
.B(n_1161),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1124),
.B(n_1113),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1143),
.A2(n_1174),
.B(n_1176),
.C(n_1125),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1101),
.B(n_1124),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1127),
.B(n_1134),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1099),
.B(n_1156),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1156),
.A2(n_1173),
.B(n_1134),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1127),
.Y(n_1276)
);

NOR4xp25_ASAP7_75t_L g1277 ( 
.A(n_1173),
.B(n_1159),
.C(n_1143),
.D(n_1162),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1134),
.B(n_1173),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1060),
.B(n_747),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1057),
.A2(n_1063),
.B(n_1145),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1145),
.A2(n_1055),
.B(n_1021),
.Y(n_1281)
);

NOR4xp25_ASAP7_75t_L g1282 ( 
.A(n_1159),
.B(n_1143),
.C(n_1162),
.D(n_1157),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1077),
.B(n_883),
.Y(n_1283)
);

O2A1O1Ixp5_ASAP7_75t_SL g1284 ( 
.A1(n_1162),
.A2(n_1066),
.B(n_1056),
.C(n_835),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1061),
.A2(n_1149),
.B(n_1139),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1057),
.A2(n_1063),
.B(n_1145),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1145),
.A2(n_1055),
.B(n_1021),
.Y(n_1287)
);

NOR4xp25_ASAP7_75t_L g1288 ( 
.A(n_1159),
.B(n_1143),
.C(n_1162),
.D(n_1157),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1060),
.B(n_747),
.Y(n_1289)
);

O2A1O1Ixp5_ASAP7_75t_L g1290 ( 
.A1(n_1056),
.A2(n_1066),
.B(n_1149),
.C(n_1055),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1291)
);

OAI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1114),
.A2(n_1146),
.B1(n_1103),
.B2(n_1056),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1060),
.B(n_737),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1157),
.A2(n_639),
.B(n_898),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1077),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1144),
.Y(n_1297)
);

NOR2x1_ASAP7_75t_R g1298 ( 
.A(n_1170),
.B(n_693),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1058),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1056),
.A2(n_1094),
.B1(n_1146),
.B2(n_1114),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1180),
.Y(n_1302)
);

AOI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1063),
.A2(n_1056),
.B(n_731),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1145),
.A2(n_1055),
.B(n_1021),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1146),
.B(n_896),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1058),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1060),
.B(n_747),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1060),
.B(n_737),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1058),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1056),
.A2(n_747),
.B(n_1063),
.C(n_1017),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1077),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1060),
.B(n_744),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1060),
.B(n_747),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1155),
.B(n_959),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1053),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1060),
.B(n_747),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_1111),
.B(n_697),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1072),
.A2(n_1150),
.B(n_1106),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1060),
.B(n_747),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1225),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1237),
.B(n_1236),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1299),
.A2(n_1316),
.B(n_1309),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1280),
.A2(n_1286),
.B(n_1182),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1221),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1221),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1280),
.A2(n_1286),
.B(n_1182),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1184),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1221),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1204),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1320),
.A2(n_1196),
.B(n_1206),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1281),
.A2(n_1304),
.B(n_1287),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1193),
.B(n_1216),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1305),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1234),
.A2(n_1186),
.B(n_1212),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1312),
.B(n_1207),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1294),
.A2(n_1308),
.B(n_1295),
.C(n_1303),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1254),
.A2(n_1227),
.B(n_1290),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1295),
.A2(n_1201),
.B(n_1303),
.C(n_1313),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1301),
.A2(n_1321),
.B1(n_1318),
.B2(n_1314),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1187),
.A2(n_1197),
.B(n_1311),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1230),
.A2(n_1269),
.B1(n_1248),
.B2(n_1249),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1189),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1235),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1181),
.B(n_1200),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1239),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1254),
.A2(n_1213),
.B(n_1197),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1199),
.B(n_1270),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1230),
.A2(n_1269),
.B1(n_1248),
.B2(n_1249),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1292),
.A2(n_1279),
.B1(n_1289),
.B2(n_1307),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1203),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1213),
.A2(n_1251),
.B(n_1215),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1317),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1200),
.B(n_1195),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1274),
.A2(n_1272),
.B1(n_1267),
.B2(n_1271),
.C(n_1247),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1274),
.A2(n_1245),
.B1(n_1201),
.B2(n_1231),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1257),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1284),
.A2(n_1222),
.B(n_1288),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1253),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1202),
.B(n_1302),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1215),
.A2(n_1256),
.B(n_1246),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1264),
.Y(n_1365)
);

INVxp67_ASAP7_75t_SL g1366 ( 
.A(n_1297),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1191),
.A2(n_1235),
.B(n_1223),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1262),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1245),
.A2(n_1231),
.B1(n_1263),
.B2(n_1319),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1282),
.A2(n_1288),
.B(n_1232),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1261),
.A2(n_1282),
.B(n_1259),
.C(n_1277),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1209),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1241),
.Y(n_1373)
);

AOI221xp5_ASAP7_75t_L g1374 ( 
.A1(n_1277),
.A2(n_1188),
.B1(n_1198),
.B2(n_1218),
.C(n_1238),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1198),
.A2(n_1242),
.B(n_1224),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1219),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1185),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1242),
.A2(n_1224),
.B(n_1223),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1194),
.A2(n_1229),
.B1(n_1192),
.B2(n_1208),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1300),
.A2(n_1306),
.B1(n_1310),
.B2(n_1243),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1209),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1238),
.A2(n_1205),
.B(n_1240),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1285),
.A2(n_1250),
.B(n_1217),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1285),
.A2(n_1250),
.B(n_1217),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1228),
.A2(n_1255),
.B1(n_1210),
.B2(n_1226),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1258),
.A2(n_1211),
.B(n_1233),
.C(n_1268),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1220),
.Y(n_1387)
);

BUFx12f_ASAP7_75t_L g1388 ( 
.A(n_1226),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1300),
.B(n_1315),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1278),
.B(n_1273),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1283),
.A2(n_1220),
.B(n_1296),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1260),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1209),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1275),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1275),
.A2(n_1244),
.B1(n_1296),
.B2(n_1268),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1283),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1276),
.B(n_1273),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1276),
.A2(n_1268),
.B(n_1244),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1190),
.A2(n_1183),
.B(n_1244),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1241),
.A2(n_1252),
.B1(n_1266),
.B2(n_1298),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1252),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1295),
.A2(n_1201),
.B(n_1303),
.C(n_1313),
.Y(n_1406)
);

BUFx2_ASAP7_75t_R g1407 ( 
.A(n_1239),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1184),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1187),
.B(n_1258),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1294),
.A2(n_747),
.B(n_1308),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1265),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1237),
.B(n_791),
.Y(n_1413)
);

AO22x1_ASAP7_75t_L g1414 ( 
.A1(n_1313),
.A2(n_731),
.B1(n_1248),
.B2(n_618),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1294),
.A2(n_747),
.B(n_1308),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1204),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1230),
.A2(n_1132),
.B1(n_1308),
.B2(n_1294),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1184),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1187),
.B(n_1258),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1313),
.B(n_1181),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1230),
.A2(n_1132),
.B1(n_1308),
.B2(n_1294),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1184),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1425)
);

NAND2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1221),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1313),
.B(n_1181),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1279),
.B(n_1146),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_SL g1432 ( 
.A1(n_1191),
.A2(n_1248),
.B(n_1057),
.C(n_1303),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1182),
.A2(n_1286),
.B(n_1280),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1235),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1184),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1184),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1182),
.A2(n_1286),
.B(n_1280),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1265),
.B(n_1312),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1280),
.A2(n_1286),
.B(n_1182),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1294),
.A2(n_747),
.B(n_1308),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1280),
.A2(n_1286),
.B(n_1182),
.Y(n_1443)
);

BUFx4f_ASAP7_75t_L g1444 ( 
.A(n_1204),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1294),
.B(n_731),
.C(n_747),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1214),
.A2(n_1293),
.B(n_1291),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1305),
.B(n_1146),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1225),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1184),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1184),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1193),
.B(n_1216),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1225),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1184),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1184),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1225),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1294),
.A2(n_1308),
.B(n_1295),
.C(n_1303),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1182),
.A2(n_1286),
.B(n_1280),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1204),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_L g1459 ( 
.A(n_1237),
.B(n_791),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1187),
.B(n_1258),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1184),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_SL g1462 ( 
.A(n_1298),
.B(n_693),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1313),
.A2(n_1301),
.B1(n_731),
.B2(n_747),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1184),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1225),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1225),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1346),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1421),
.B(n_1428),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1363),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1458),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1418),
.A2(n_1423),
.B1(n_1352),
.B2(n_1345),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1383),
.A2(n_1384),
.B(n_1361),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1344),
.A2(n_1335),
.B(n_1433),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1357),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1331),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1418),
.A2(n_1423),
.B1(n_1352),
.B2(n_1345),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1463),
.A2(n_1342),
.B(n_1406),
.C(n_1343),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1340),
.A2(n_1456),
.B(n_1342),
.C(n_1406),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1326),
.A2(n_1334),
.B(n_1322),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1445),
.A2(n_1415),
.B(n_1411),
.Y(n_1480)
);

BUFx2_ASAP7_75t_SL g1481 ( 
.A(n_1413),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1438),
.A2(n_1457),
.B(n_1367),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1369),
.B(n_1353),
.Y(n_1483)
);

OAI31xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1379),
.A2(n_1370),
.A3(n_1414),
.B(n_1442),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1371),
.A2(n_1369),
.B(n_1374),
.C(n_1358),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1432),
.A2(n_1348),
.B(n_1430),
.C(n_1337),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1458),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1360),
.B(n_1366),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1447),
.B(n_1390),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1385),
.B(n_1368),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1385),
.B(n_1362),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1359),
.A2(n_1327),
.B1(n_1443),
.B2(n_1440),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1386),
.A2(n_1359),
.B(n_1389),
.C(n_1420),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1389),
.A2(n_1460),
.B(n_1410),
.C(n_1420),
.Y(n_1494)
);

CKINVDCx16_ASAP7_75t_R g1495 ( 
.A(n_1462),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1334),
.A2(n_1322),
.B(n_1446),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1327),
.B(n_1330),
.Y(n_1497)
);

OA22x2_ASAP7_75t_L g1498 ( 
.A1(n_1380),
.A2(n_1401),
.B1(n_1399),
.B2(n_1461),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1330),
.A2(n_1440),
.B1(n_1443),
.B2(n_1395),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1440),
.A2(n_1443),
.B1(n_1434),
.B2(n_1347),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1347),
.A2(n_1434),
.B1(n_1464),
.B2(n_1449),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1410),
.A2(n_1460),
.B(n_1420),
.C(n_1377),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1459),
.A2(n_1325),
.B(n_1409),
.C(n_1424),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1410),
.A2(n_1460),
.B(n_1376),
.C(n_1356),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1403),
.A2(n_1429),
.B(n_1404),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1354),
.B(n_1419),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1436),
.A2(n_1454),
.B(n_1453),
.C(n_1450),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1437),
.A2(n_1341),
.B1(n_1350),
.B2(n_1378),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1341),
.A2(n_1350),
.B1(n_1378),
.B2(n_1407),
.Y(n_1509)
);

NOR2xp67_ASAP7_75t_L g1510 ( 
.A(n_1388),
.B(n_1365),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1416),
.A2(n_1388),
.B1(n_1365),
.B2(n_1349),
.Y(n_1511)
);

AND2x6_ASAP7_75t_L g1512 ( 
.A(n_1329),
.B(n_1332),
.Y(n_1512)
);

AOI221x1_ASAP7_75t_SL g1513 ( 
.A1(n_1394),
.A2(n_1393),
.B1(n_1381),
.B2(n_1372),
.C(n_1466),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1387),
.B(n_1350),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1396),
.B(n_1375),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1329),
.A2(n_1332),
.B(n_1328),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_R g1518 ( 
.A(n_1349),
.B(n_1416),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1375),
.B(n_1397),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1382),
.B(n_1375),
.C(n_1355),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1382),
.B(n_1323),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1333),
.B(n_1444),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1397),
.B(n_1373),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1373),
.B(n_1398),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1339),
.A2(n_1324),
.B(n_1417),
.C(n_1439),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1339),
.A2(n_1324),
.B(n_1417),
.C(n_1439),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1373),
.B(n_1398),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1373),
.B(n_1412),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1412),
.B(n_1332),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1427),
.B(n_1465),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1391),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1400),
.B(n_1455),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1364),
.B(n_1402),
.Y(n_1534)
);

AOI21x1_ASAP7_75t_SL g1535 ( 
.A1(n_1402),
.A2(n_1444),
.B(n_1392),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1435),
.B(n_1392),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1448),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1364),
.B(n_1452),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1405),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1408),
.B(n_1425),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1431),
.B(n_1441),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1338),
.A2(n_1344),
.B(n_1335),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1463),
.A2(n_1294),
.B(n_1308),
.C(n_1295),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1357),
.B(n_1363),
.Y(n_1544)
);

OA22x2_ASAP7_75t_L g1545 ( 
.A1(n_1353),
.A2(n_1295),
.B1(n_1274),
.B2(n_1248),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1336),
.B(n_1451),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1343),
.A2(n_1248),
.B(n_1201),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1331),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1344),
.A2(n_1335),
.B(n_1303),
.Y(n_1549)
);

AOI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1414),
.A2(n_1463),
.B(n_731),
.C(n_747),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1418),
.A2(n_1099),
.B1(n_1313),
.B2(n_1301),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1348),
.B(n_1370),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1421),
.B(n_1428),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1357),
.B(n_1363),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1368),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1418),
.A2(n_1423),
.B1(n_1165),
.B2(n_1157),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1344),
.A2(n_1335),
.B(n_1303),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1340),
.A2(n_747),
.B(n_1295),
.C(n_731),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1418),
.A2(n_1423),
.B1(n_1165),
.B2(n_1157),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1363),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1463),
.A2(n_1294),
.B(n_1308),
.C(n_1295),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1421),
.B(n_1428),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1463),
.A2(n_1294),
.B(n_1308),
.C(n_1295),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1348),
.B(n_1370),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1351),
.B(n_1146),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1562),
.A2(n_1478),
.B(n_1477),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1473),
.A2(n_1520),
.B(n_1482),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1475),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1521),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1521),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1502),
.A2(n_1563),
.B(n_1560),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1499),
.B(n_1515),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1539),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1518),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1549),
.A2(n_1561),
.B(n_1542),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1532),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1508),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1512),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1474),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1534),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1479),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1548),
.Y(n_1590)
);

BUFx4f_ASAP7_75t_SL g1591 ( 
.A(n_1467),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1492),
.B(n_1514),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1552),
.B(n_1569),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1470),
.Y(n_1595)
);

OAI31xp33_ASAP7_75t_L g1596 ( 
.A1(n_1560),
.A2(n_1563),
.A3(n_1471),
.B(n_1476),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1512),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1504),
.B(n_1494),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1509),
.A2(n_1492),
.B(n_1516),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1534),
.B(n_1547),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1534),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1531),
.B(n_1540),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1469),
.B(n_1552),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1505),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1513),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1500),
.B(n_1472),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1472),
.B(n_1536),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1507),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1496),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1537),
.B(n_1541),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1501),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1569),
.A2(n_1485),
.B(n_1530),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1506),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1564),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1490),
.A2(n_1491),
.B(n_1558),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1480),
.A2(n_1493),
.B(n_1471),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1476),
.B(n_1551),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1545),
.B(n_1553),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1543),
.A2(n_1565),
.B(n_1567),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1545),
.B(n_1484),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1488),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1544),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1556),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1484),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1498),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1576),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1468),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1498),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1483),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1572),
.B(n_1559),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1594),
.B(n_1554),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1580),
.B(n_1557),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1580),
.B(n_1555),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1595),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1574),
.B(n_1489),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1588),
.B(n_1546),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1574),
.B(n_1503),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1601),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1589),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1584),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1589),
.Y(n_1645)
);

OAI211xp5_ASAP7_75t_L g1646 ( 
.A1(n_1618),
.A2(n_1550),
.B(n_1486),
.C(n_1570),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1528),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1608),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1580),
.B(n_1571),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1588),
.B(n_1601),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1577),
.B(n_1529),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1617),
.A2(n_1526),
.B(n_1525),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1603),
.B(n_1533),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1578),
.B(n_1568),
.Y(n_1654)
);

NAND2x1_ASAP7_75t_L g1655 ( 
.A(n_1586),
.B(n_1512),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1592),
.B(n_1523),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1607),
.B(n_1527),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1524),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1584),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1575),
.A2(n_1535),
.B(n_1517),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1586),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_R g1662 ( 
.A(n_1638),
.B(n_1582),
.Y(n_1662)
);

OAI211xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1646),
.A2(n_1573),
.B(n_1596),
.C(n_1579),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1646),
.A2(n_1596),
.B(n_1618),
.C(n_1625),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1628),
.A2(n_1621),
.B1(n_1619),
.B2(n_1598),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1650),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1641),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1641),
.B(n_1621),
.C(n_1612),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1639),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1648),
.A2(n_1621),
.B1(n_1619),
.B2(n_1626),
.C(n_1617),
.Y(n_1671)
);

AO21x1_ASAP7_75t_SL g1672 ( 
.A1(n_1641),
.A2(n_1605),
.B(n_1613),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1652),
.A2(n_1619),
.B1(n_1598),
.B2(n_1626),
.C(n_1581),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1637),
.B(n_1653),
.Y(n_1675)
);

OAI211xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1648),
.A2(n_1608),
.B(n_1622),
.C(n_1587),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1587),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1632),
.B(n_1591),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1632),
.A2(n_1647),
.B(n_1605),
.C(n_1611),
.Y(n_1681)
);

AOI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1634),
.A2(n_1611),
.B1(n_1617),
.B2(n_1622),
.C1(n_1623),
.C2(n_1624),
.Y(n_1682)
);

O2A1O1Ixp5_ASAP7_75t_L g1683 ( 
.A1(n_1655),
.A2(n_1585),
.B(n_1597),
.C(n_1586),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1647),
.A2(n_1598),
.B(n_1612),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1639),
.B(n_1495),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1634),
.A2(n_1617),
.B1(n_1620),
.B2(n_1598),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1639),
.B(n_1581),
.Y(n_1688)
);

AOI33xp33_ASAP7_75t_L g1689 ( 
.A1(n_1634),
.A2(n_1593),
.A3(n_1624),
.B1(n_1623),
.B2(n_1606),
.B3(n_1590),
.Y(n_1689)
);

OAI31xp33_ASAP7_75t_L g1690 ( 
.A1(n_1633),
.A2(n_1581),
.A3(n_1617),
.B(n_1642),
.Y(n_1690)
);

NOR4xp25_ASAP7_75t_L g1691 ( 
.A(n_1629),
.B(n_1606),
.C(n_1585),
.D(n_1613),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1654),
.A2(n_1598),
.B1(n_1581),
.B2(n_1600),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1635),
.A2(n_1620),
.B1(n_1615),
.B2(n_1593),
.C(n_1614),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1655),
.B(n_1598),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1661),
.B(n_1598),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1654),
.B(n_1612),
.C(n_1616),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1610),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1649),
.A2(n_1600),
.B1(n_1606),
.B2(n_1593),
.C(n_1620),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1695),
.B(n_1659),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1685),
.A2(n_1604),
.B(n_1609),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1667),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1668),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1691),
.B(n_1640),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1664),
.B(n_1649),
.C(n_1655),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1694),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1697),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1697),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1697),
.Y(n_1710)
);

INVx5_ASAP7_75t_L g1711 ( 
.A(n_1666),
.Y(n_1711)
);

AOI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1681),
.A2(n_1645),
.B(n_1643),
.Y(n_1712)
);

OR2x2_ASAP7_75t_SL g1713 ( 
.A(n_1669),
.B(n_1612),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1698),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1663),
.A2(n_1620),
.B(n_1660),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1670),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1683),
.Y(n_1719)
);

INVx4_ASAP7_75t_SL g1720 ( 
.A(n_1684),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1684),
.Y(n_1722)
);

INVx4_ASAP7_75t_SL g1723 ( 
.A(n_1696),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1671),
.B(n_1640),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1693),
.B(n_1630),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1720),
.B(n_1677),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1721),
.B(n_1675),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1707),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1714),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1714),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1720),
.B(n_1696),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1720),
.B(n_1699),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1706),
.A2(n_1663),
.B1(n_1674),
.B2(n_1665),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1717),
.B(n_1690),
.C(n_1687),
.D(n_1682),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1704),
.B(n_1700),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1707),
.B(n_1661),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1704),
.Y(n_1738)
);

OAI332xp33_ASAP7_75t_L g1739 ( 
.A1(n_1721),
.A2(n_1511),
.A3(n_1692),
.B1(n_1673),
.B2(n_1678),
.B3(n_1686),
.C1(n_1688),
.C2(n_1680),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1717),
.A2(n_1676),
.B(n_1629),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_R g1741 ( 
.A(n_1706),
.B(n_1487),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1715),
.B(n_1718),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1720),
.B(n_1657),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1704),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1707),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1658),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1705),
.B(n_1676),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1705),
.A2(n_1724),
.B(n_1715),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1704),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1631),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1715),
.B(n_1656),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1725),
.A2(n_1599),
.B1(n_1600),
.B2(n_1660),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1711),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1633),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1703),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1636),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1714),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1703),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1713),
.B(n_1651),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1708),
.B(n_1522),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1723),
.B(n_1636),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1755),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1755),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1758),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1728),
.B(n_1725),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1747),
.A2(n_1724),
.B1(n_1710),
.B2(n_1708),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1729),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1726),
.B(n_1723),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.B(n_1723),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1758),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1709),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1738),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.B(n_1709),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1738),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1739),
.B(n_1716),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1732),
.B(n_1709),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1760),
.B(n_1591),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1744),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1713),
.Y(n_1779)
);

AOI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1748),
.A2(n_1716),
.B(n_1719),
.C(n_1710),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1730),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1730),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1729),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1732),
.B(n_1722),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1731),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1716),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1744),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1742),
.B(n_1701),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1747),
.B(n_1716),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_R g1792 ( 
.A(n_1741),
.B(n_1481),
.Y(n_1792)
);

NOR2xp67_ASAP7_75t_L g1793 ( 
.A(n_1753),
.B(n_1722),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1743),
.B(n_1746),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1743),
.B(n_1722),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_L g1796 ( 
.A(n_1734),
.B(n_1662),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1731),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_SL g1798 ( 
.A(n_1737),
.B(n_1661),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1794),
.B(n_1737),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1775),
.A2(n_1735),
.B1(n_1752),
.B2(n_1736),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1767),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1787),
.B(n_1757),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1783),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1762),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1762),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_R g1806 ( 
.A(n_1796),
.B(n_1737),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1797),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1767),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1768),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1791),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1776),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1790),
.B(n_1757),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1776),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1763),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1794),
.B(n_1754),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1766),
.A2(n_1753),
.B(n_1719),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1771),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1780),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.B(n_1749),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1764),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1768),
.B(n_1754),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1798),
.B(n_1740),
.Y(n_1822)
);

INVx3_ASAP7_75t_SL g1823 ( 
.A(n_1769),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1769),
.B(n_1754),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1796),
.A2(n_1735),
.B1(n_1702),
.B2(n_1583),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1771),
.B(n_1754),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1800),
.A2(n_1765),
.B1(n_1779),
.B2(n_1785),
.Y(n_1827)
);

OAI32xp33_ASAP7_75t_L g1828 ( 
.A1(n_1800),
.A2(n_1779),
.A3(n_1785),
.B1(n_1745),
.B2(n_1719),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1826),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1812),
.Y(n_1830)
);

OAI322xp33_ASAP7_75t_L g1831 ( 
.A1(n_1818),
.A2(n_1745),
.A3(n_1789),
.B1(n_1781),
.B2(n_1782),
.C1(n_1786),
.C2(n_1759),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1818),
.A2(n_1702),
.B1(n_1719),
.B2(n_1773),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1822),
.A2(n_1773),
.B1(n_1784),
.B2(n_1795),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1812),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1825),
.A2(n_1793),
.B(n_1784),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1812),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1801),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1801),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1817),
.A2(n_1712),
.B1(n_1702),
.B2(n_1789),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1821),
.B(n_1795),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1826),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1817),
.B(n_1770),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1809),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1803),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1825),
.B(n_1777),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1802),
.A2(n_1727),
.B1(n_1761),
.B2(n_1756),
.C(n_1759),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1845),
.B(n_1803),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1829),
.B(n_1811),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1842),
.B(n_1811),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1846),
.B(n_1823),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1830),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1840),
.B(n_1810),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1833),
.B(n_1823),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1845),
.B(n_1810),
.Y(n_1855)
);

NAND2x1_ASAP7_75t_L g1856 ( 
.A(n_1834),
.B(n_1799),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1836),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1837),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1843),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1827),
.B(n_1811),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1851),
.A2(n_1835),
.B1(n_1846),
.B2(n_1832),
.C(n_1802),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1855),
.A2(n_1828),
.B1(n_1831),
.B2(n_1839),
.C(n_1832),
.Y(n_1862)
);

AOI322xp5_ASAP7_75t_L g1863 ( 
.A1(n_1854),
.A2(n_1847),
.A3(n_1839),
.B1(n_1807),
.B2(n_1813),
.C1(n_1799),
.C2(n_1838),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1853),
.A2(n_1824),
.B1(n_1821),
.B2(n_1823),
.Y(n_1864)
);

AOI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1855),
.A2(n_1859),
.B1(n_1848),
.B2(n_1860),
.C(n_1806),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1856),
.B(n_1809),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1849),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1848),
.A2(n_1807),
.B1(n_1857),
.B2(n_1852),
.C(n_1813),
.Y(n_1868)
);

HAxp5_ASAP7_75t_SL g1869 ( 
.A(n_1858),
.B(n_1841),
.CON(n_1869),
.SN(n_1869)
);

OAI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1850),
.A2(n_1824),
.B(n_1821),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1849),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1851),
.B(n_1799),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1851),
.B(n_1813),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1867),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1869),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1861),
.A2(n_1809),
.B1(n_1824),
.B2(n_1826),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1862),
.A2(n_1844),
.B(n_1808),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1865),
.A2(n_1809),
.B1(n_1820),
.B2(n_1814),
.C(n_1808),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1870),
.B(n_1809),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1866),
.Y(n_1880)
);

XNOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1510),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1880),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1875),
.B(n_1871),
.Y(n_1883)
);

CKINVDCx14_ASAP7_75t_R g1884 ( 
.A(n_1874),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1876),
.B(n_1872),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1879),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1878),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1877),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1882),
.B(n_1868),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1883),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1884),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1886),
.B(n_1873),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1885),
.A2(n_1881),
.B1(n_1808),
.B2(n_1815),
.Y(n_1893)
);

NAND3x1_ASAP7_75t_L g1894 ( 
.A(n_1888),
.B(n_1820),
.C(n_1814),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1891),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1893),
.A2(n_1884),
.B1(n_1887),
.B2(n_1819),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1889),
.A2(n_1816),
.B(n_1805),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1895),
.B(n_1892),
.Y(n_1898)
);

AOI211xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1898),
.A2(n_1896),
.B(n_1890),
.C(n_1897),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1894),
.B(n_1863),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1899),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1900),
.A2(n_1805),
.B(n_1804),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1901),
.B(n_1804),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1903),
.Y(n_1904)
);

AO22x2_ASAP7_75t_L g1905 ( 
.A1(n_1902),
.A2(n_1819),
.B1(n_1815),
.B2(n_1774),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1904),
.B(n_1819),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1906),
.B(n_1905),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1907),
.B(n_1816),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1816),
.B1(n_1815),
.B2(n_1772),
.Y(n_1909)
);

AOI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1788),
.B1(n_1778),
.B2(n_1774),
.C(n_1772),
.Y(n_1910)
);

AOI211xp5_ASAP7_75t_L g1911 ( 
.A1(n_1910),
.A2(n_1792),
.B(n_1788),
.C(n_1778),
.Y(n_1911)
);


endmodule