module real_aes_16863_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_836, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_836;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g827 ( .A(n_0), .B(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_1), .A2(n_3), .B1(n_124), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_2), .A2(n_43), .B1(n_131), .B2(n_237), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_4), .A2(n_24), .B1(n_202), .B2(n_237), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_5), .A2(n_15), .B1(n_121), .B2(n_170), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_6), .A2(n_59), .B1(n_149), .B2(n_204), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_7), .A2(n_17), .B1(n_131), .B2(n_153), .Y(n_516) );
INVx1_ASAP7_75t_L g828 ( .A(n_8), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_9), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_10), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_11), .A2(n_19), .B1(n_148), .B2(n_151), .Y(n_147) );
OR2x2_ASAP7_75t_L g789 ( .A(n_12), .B(n_40), .Y(n_789) );
BUFx2_ASAP7_75t_L g832 ( .A(n_12), .Y(n_832) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_14), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_16), .A2(n_102), .B1(n_824), .B2(n_833), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g805 ( .A1(n_18), .A2(n_71), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_18), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_20), .A2(n_99), .B1(n_121), .B2(n_124), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_21), .A2(n_39), .B1(n_165), .B2(n_167), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_122), .Y(n_215) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_23), .A2(n_57), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_25), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_26), .Y(n_611) );
INVx4_ASAP7_75t_R g528 ( .A(n_27), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_28), .B(n_128), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_29), .A2(n_47), .B1(n_181), .B2(n_183), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_30), .A2(n_66), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_30), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_31), .A2(n_53), .B1(n_121), .B2(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_32), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_33), .B(n_165), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_34), .Y(n_228) );
INVx1_ASAP7_75t_L g541 ( .A(n_35), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_36), .B(n_237), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_37), .A2(n_127), .B(n_131), .C(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_38), .A2(n_54), .B1(n_131), .B2(n_183), .Y(n_609) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_40), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_41), .A2(n_86), .B1(n_131), .B2(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_42), .A2(n_46), .B1(n_131), .B2(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_44), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_45), .A2(n_58), .B1(n_121), .B2(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g563 ( .A(n_48), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_49), .B(n_131), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_50), .Y(n_503) );
INVx2_ASAP7_75t_L g799 ( .A(n_51), .Y(n_799) );
BUFx3_ASAP7_75t_L g788 ( .A(n_52), .Y(n_788) );
INVx1_ASAP7_75t_L g816 ( .A(n_52), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_55), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_56), .A2(n_87), .B1(n_131), .B2(n_183), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_60), .A2(n_74), .B1(n_130), .B2(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_61), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_62), .A2(n_76), .B1(n_131), .B2(n_153), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_63), .A2(n_98), .B1(n_121), .B2(n_151), .Y(n_225) );
AND2x4_ASAP7_75t_L g117 ( .A(n_64), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
INVx1_ASAP7_75t_L g783 ( .A(n_66), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_67), .A2(n_90), .B1(n_181), .B2(n_183), .Y(n_537) );
AO22x1_ASAP7_75t_L g494 ( .A1(n_68), .A2(n_75), .B1(n_167), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g118 ( .A(n_69), .Y(n_118) );
AND2x2_ASAP7_75t_L g481 ( .A(n_70), .B(n_221), .Y(n_481) );
INVx1_ASAP7_75t_L g806 ( .A(n_71), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_72), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_73), .B(n_204), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_77), .B(n_237), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_78), .Y(n_793) );
INVx2_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_80), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_81), .B(n_221), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_82), .A2(n_97), .B1(n_183), .B2(n_204), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_83), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_84), .B(n_138), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_85), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_88), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_89), .B(n_221), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_91), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_92), .B(n_221), .Y(n_500) );
INVx1_ASAP7_75t_L g461 ( .A(n_93), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_93), .B(n_815), .Y(n_814) );
NAND2xp33_ASAP7_75t_L g218 ( .A(n_94), .B(n_122), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_95), .A2(n_155), .B(n_204), .C(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g530 ( .A(n_96), .B(n_531), .Y(n_530) );
NAND2xp33_ASAP7_75t_L g508 ( .A(n_100), .B(n_166), .Y(n_508) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_795), .B(n_800), .Y(n_102) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_781), .B(n_790), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_104), .A2(n_791), .B1(n_792), .B2(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_458), .B1(n_462), .B2(n_779), .Y(n_105) );
INVx2_ASAP7_75t_L g808 ( .A(n_106), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_106), .B(n_810), .Y(n_809) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_367), .Y(n_106) );
NOR2x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_306), .Y(n_107) );
NAND4xp25_ASAP7_75t_L g108 ( .A(n_109), .B(n_257), .C(n_276), .D(n_287), .Y(n_108) );
O2A1O1Ixp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_188), .B(n_195), .C(n_229), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_160), .Y(n_110) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_111), .B(n_322), .C(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g403 ( .A(n_111), .B(n_285), .Y(n_403) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_144), .Y(n_111) );
AND2x2_ASAP7_75t_L g247 ( .A(n_112), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g265 ( .A(n_112), .B(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g282 ( .A(n_112), .Y(n_282) );
AND2x2_ASAP7_75t_L g327 ( .A(n_112), .B(n_162), .Y(n_327) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g192 ( .A(n_113), .Y(n_192) );
AND2x4_ASAP7_75t_L g275 ( .A(n_113), .B(n_266), .Y(n_275) );
AO31x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .A3(n_135), .B(n_141), .Y(n_113) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_114), .A2(n_156), .A3(n_224), .B(n_227), .Y(n_223) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_115), .A2(n_523), .B(n_526), .Y(n_522) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_116), .A2(n_146), .A3(n_156), .B(n_158), .Y(n_145) );
AO31x2_ASAP7_75t_L g162 ( .A1(n_116), .A2(n_163), .A3(n_172), .B(n_174), .Y(n_162) );
AO31x2_ASAP7_75t_L g234 ( .A1(n_116), .A2(n_235), .A3(n_239), .B(n_240), .Y(n_234) );
AO31x2_ASAP7_75t_L g514 ( .A1(n_116), .A2(n_143), .A3(n_515), .B(n_518), .Y(n_514) );
BUFx10_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g185 ( .A(n_117), .Y(n_185) );
INVx1_ASAP7_75t_L g480 ( .A(n_117), .Y(n_480) );
BUFx10_ASAP7_75t_L g512 ( .A(n_117), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B1(n_129), .B2(n_132), .Y(n_119) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_122), .Y(n_495) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g125 ( .A(n_123), .Y(n_125) );
INVx3_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
INVx1_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_123), .Y(n_168) );
INVx1_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_123), .Y(n_183) );
INVx2_ASAP7_75t_L g202 ( .A(n_123), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_123), .Y(n_204) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_123), .Y(n_237) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_125), .B(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_126), .A2(n_147), .B1(n_152), .B2(n_154), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_126), .A2(n_132), .B1(n_164), .B2(n_169), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_126), .A2(n_132), .B1(n_180), .B2(n_182), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_126), .A2(n_200), .B1(n_203), .B2(n_205), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_126), .A2(n_217), .B(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_126), .A2(n_154), .B1(n_225), .B2(n_226), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_126), .A2(n_132), .B1(n_236), .B2(n_238), .Y(n_235) );
OAI22x1_ASAP7_75t_L g515 ( .A1(n_126), .A2(n_205), .B1(n_516), .B2(n_517), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_126), .A2(n_205), .B1(n_537), .B2(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_126), .A2(n_490), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx6_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
O2A1O1Ixp5_ASAP7_75t_L g213 ( .A1(n_127), .A2(n_153), .B(n_214), .C(n_215), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_127), .B(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_127), .A2(n_508), .B(n_509), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_127), .A2(n_489), .B(n_494), .C(n_497), .Y(n_549) );
BUFx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
INVx1_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
INVx1_ASAP7_75t_L g476 ( .A(n_128), .Y(n_476) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
INVx4_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g490 ( .A(n_133), .Y(n_490) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g506 ( .A(n_134), .Y(n_506) );
AO31x2_ASAP7_75t_L g178 ( .A1(n_135), .A2(n_179), .A3(n_184), .B(n_186), .Y(n_178) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_135), .A2(n_522), .B(n_530), .Y(n_521) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g158 ( .A(n_137), .B(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_137), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g143 ( .A(n_138), .Y(n_143) );
INVx2_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_138), .A2(n_480), .B(n_492), .Y(n_497) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_143), .B(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g193 ( .A(n_144), .B(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g250 ( .A(n_144), .B(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_144), .Y(n_273) );
INVx1_ASAP7_75t_L g284 ( .A(n_144), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_144), .B(n_176), .Y(n_293) );
INVx2_ASAP7_75t_L g300 ( .A(n_144), .Y(n_300) );
INVx4_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g245 ( .A(n_145), .B(n_162), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_145), .B(n_252), .Y(n_318) );
AND2x2_ASAP7_75t_L g326 ( .A(n_145), .B(n_178), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_145), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g379 ( .A(n_145), .Y(n_379) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_150), .B(n_525), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_153), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
INVx1_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
AOI21x1_ASAP7_75t_L g468 ( .A1(n_156), .A2(n_469), .B(n_481), .Y(n_468) );
AO31x2_ASAP7_75t_L g535 ( .A1(n_156), .A2(n_184), .A3(n_536), .B(n_540), .Y(n_535) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_157), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g531 ( .A(n_157), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_157), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_157), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g395 ( .A(n_161), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_176), .Y(n_161) );
INVx1_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
INVx1_ASAP7_75t_L g252 ( .A(n_162), .Y(n_252) );
INVx2_ASAP7_75t_L g286 ( .A(n_162), .Y(n_286) );
OR2x2_ASAP7_75t_L g290 ( .A(n_162), .B(n_178), .Y(n_290) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_162), .Y(n_339) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_166), .A2(n_171), .B1(n_528), .B2(n_529), .Y(n_527) );
OAI21xp33_ASAP7_75t_SL g559 ( .A1(n_167), .A2(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_172), .A2(n_184), .A3(n_199), .B(n_206), .Y(n_198) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_173), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_SL g211 ( .A(n_173), .Y(n_211) );
INVx4_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_173), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_173), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g567 ( .A(n_173), .B(n_512), .Y(n_567) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x2_ASAP7_75t_L g312 ( .A(n_177), .B(n_192), .Y(n_312) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
INVx2_ASAP7_75t_L g266 ( .A(n_178), .Y(n_266) );
AND2x4_ASAP7_75t_L g285 ( .A(n_178), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g373 ( .A(n_178), .Y(n_373) );
INVx2_ASAP7_75t_L g539 ( .A(n_183), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_183), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g219 ( .A(n_185), .Y(n_219) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_193), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g291 ( .A(n_191), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_191), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g354 ( .A(n_192), .Y(n_354) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2x1_ASAP7_75t_L g196 ( .A(n_197), .B(n_208), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_197), .B(n_209), .Y(n_304) );
INVx1_ASAP7_75t_L g402 ( .A(n_197), .Y(n_402) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g242 ( .A(n_198), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g256 ( .A(n_198), .B(n_234), .Y(n_256) );
AND2x4_ASAP7_75t_L g279 ( .A(n_198), .B(n_222), .Y(n_279) );
INVx2_ASAP7_75t_L g296 ( .A(n_198), .Y(n_296) );
AND2x2_ASAP7_75t_L g322 ( .A(n_198), .B(n_223), .Y(n_322) );
INVx1_ASAP7_75t_L g387 ( .A(n_198), .Y(n_387) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_202), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_205), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g347 ( .A(n_208), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_222), .Y(n_208) );
AND2x2_ASAP7_75t_L g313 ( .A(n_209), .B(n_270), .Y(n_313) );
AND2x4_ASAP7_75t_L g329 ( .A(n_209), .B(n_296), .Y(n_329) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx2_ASAP7_75t_L g323 ( .A(n_210), .Y(n_323) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_210) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_244) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_219), .Y(n_212) );
INVx2_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_221), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
INVx3_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_222), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_222), .B(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g295 ( .A(n_223), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g419 ( .A(n_223), .Y(n_419) );
OAI33xp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_245), .A3(n_246), .B1(n_247), .B2(n_249), .B3(n_253), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2x1_ASAP7_75t_L g231 ( .A(n_232), .B(n_242), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g353 ( .A(n_233), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g262 ( .A(n_234), .B(n_244), .Y(n_262) );
INVx2_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
INVx1_ASAP7_75t_L g278 ( .A(n_234), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_237), .B(n_472), .Y(n_471) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_239), .A2(n_512), .A3(n_607), .B(n_610), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_242), .A2(n_298), .B1(n_301), .B2(n_305), .Y(n_297) );
OR2x2_ASAP7_75t_L g437 ( .A(n_242), .B(n_255), .Y(n_437) );
AND2x4_ASAP7_75t_L g341 ( .A(n_243), .B(n_303), .Y(n_341) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_244), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_245), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g305 ( .A(n_245), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_245), .B(n_281), .Y(n_383) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g356 ( .A(n_247), .Y(n_356) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g414 ( .A(n_250), .B(n_282), .Y(n_414) );
NAND2x1_ASAP7_75t_L g432 ( .A(n_250), .B(n_281), .Y(n_432) );
AND2x2_ASAP7_75t_L g456 ( .A(n_250), .B(n_275), .Y(n_456) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g446 ( .A(n_254), .B(n_323), .Y(n_446) );
NOR2x1p5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g380 ( .A(n_255), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g348 ( .A(n_256), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_263), .B1(n_267), .B2(n_271), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g355 ( .A(n_260), .B(n_323), .Y(n_355) );
AND2x2_ASAP7_75t_L g392 ( .A(n_260), .B(n_341), .Y(n_392) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g267 ( .A(n_261), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_261), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g433 ( .A(n_261), .B(n_262), .Y(n_433) );
AND2x2_ASAP7_75t_L g294 ( .A(n_262), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g413 ( .A(n_262), .B(n_279), .Y(n_413) );
AND2x2_ASAP7_75t_L g457 ( .A(n_262), .B(n_322), .Y(n_457) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_267), .A2(n_392), .B1(n_393), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_391) );
AND2x2_ASAP7_75t_L g314 ( .A(n_268), .B(n_282), .Y(n_314) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g345 ( .A(n_269), .Y(n_345) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_269), .Y(n_390) );
INVx2_ASAP7_75t_L g303 ( .A(n_270), .Y(n_303) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g360 ( .A(n_273), .Y(n_360) );
INVx2_ASAP7_75t_L g366 ( .A(n_274), .Y(n_366) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g350 ( .A(n_275), .B(n_339), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x4_ASAP7_75t_L g381 ( .A(n_278), .B(n_329), .Y(n_381) );
INVx2_ASAP7_75t_L g428 ( .A(n_278), .Y(n_428) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g371 ( .A(n_282), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g405 ( .A(n_282), .B(n_290), .Y(n_405) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g310 ( .A(n_284), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g417 ( .A(n_285), .B(n_333), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B(n_294), .C(n_297), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g298 ( .A(n_290), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_291), .B(n_326), .Y(n_430) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g406 ( .A(n_293), .B(n_375), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_295), .B(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_295), .A2(n_311), .B1(n_353), .B2(n_355), .Y(n_352) );
AND2x2_ASAP7_75t_L g358 ( .A(n_295), .B(n_323), .Y(n_358) );
AND2x2_ASAP7_75t_L g427 ( .A(n_295), .B(n_428), .Y(n_427) );
O2A1O1Ixp33_ASAP7_75t_L g420 ( .A1(n_298), .A2(n_400), .B(n_421), .C(n_424), .Y(n_420) );
INVx2_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g411 ( .A(n_303), .Y(n_411) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_305), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_351) );
NAND3xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_319), .C(n_342), .Y(n_306) );
AO22x1_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .B1(n_314), .B2(n_315), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_312), .Y(n_445) );
OR2x2_ASAP7_75t_L g452 ( .A(n_312), .B(n_333), .Y(n_452) );
AND2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_322), .Y(n_364) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g440 ( .A(n_318), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .C(n_330), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
AND2x4_ASAP7_75t_SL g398 ( .A(n_322), .B(n_341), .Y(n_398) );
INVx1_ASAP7_75t_SL g409 ( .A(n_322), .Y(n_409) );
OR2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x4_ASAP7_75t_L g338 ( .A(n_326), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g396 ( .A(n_327), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g418 ( .A(n_329), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_329), .B(n_423), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_337), .B2(n_340), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x4_ASAP7_75t_L g378 ( .A(n_334), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g400 ( .A(n_334), .Y(n_400) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g455 ( .A(n_338), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_351), .C(n_359), .Y(n_342) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g424 ( .A(n_345), .Y(n_424) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_350), .A2(n_448), .B1(n_451), .B2(n_453), .C1(n_455), .C2(n_457), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_353), .B(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B(n_363), .C(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_425), .Y(n_367) );
NAND4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_391), .C(n_401), .D(n_412), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_380), .B1(n_382), .B2(n_384), .Y(n_369) );
NAND3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .C(n_377), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_371), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_375), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g422 ( .A(n_387), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_389), .Y(n_454) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g449 ( .A(n_398), .Y(n_449) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .C(n_410), .Y(n_401) );
AOI21xp33_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_406), .B(n_407), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_405), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_415), .B2(n_418), .C(n_420), .Y(n_412) );
INVx1_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
AOI31xp33_ASAP7_75t_L g434 ( .A1(n_416), .A2(n_435), .A3(n_436), .B(n_437), .Y(n_434) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_419), .Y(n_423) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_438), .C(n_447), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_426) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g435 ( .A(n_433), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_444), .B2(n_446), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR3x1_ASAP7_75t_L g825 ( .A(n_460), .B(n_788), .C(n_826), .Y(n_825) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g780 ( .A(n_461), .Y(n_780) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_679), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_582), .C(n_641), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_482), .B1(n_569), .B2(n_575), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g638 ( .A(n_467), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_467), .B(n_556), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_467), .B(n_602), .Y(n_749) );
AND2x2_ASAP7_75t_L g755 ( .A(n_467), .B(n_581), .Y(n_755) );
INVxp67_ASAP7_75t_L g760 ( .A(n_467), .Y(n_760) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g573 ( .A(n_468), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_477), .B(n_480), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B(n_475), .Y(n_470) );
BUFx4f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_476), .B(n_563), .Y(n_562) );
OAI21xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_532), .B(n_542), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_513), .Y(n_484) );
INVx1_ASAP7_75t_L g676 ( .A(n_485), .Y(n_676) );
AND2x2_ASAP7_75t_L g705 ( .A(n_485), .B(n_667), .Y(n_705) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .Y(n_485) );
AND2x2_ASAP7_75t_L g599 ( .A(n_486), .B(n_521), .Y(n_599) );
INVx1_ASAP7_75t_L g654 ( .A(n_486), .Y(n_654) );
AND2x2_ASAP7_75t_L g704 ( .A(n_486), .B(n_520), .Y(n_704) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g579 ( .A(n_487), .B(n_520), .Y(n_579) );
AND2x4_ASAP7_75t_L g723 ( .A(n_487), .B(n_521), .Y(n_723) );
AOI21x1_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_493), .B(n_496), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI21x1_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_490), .A2(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g648 ( .A(n_498), .Y(n_648) );
AND2x2_ASAP7_75t_L g717 ( .A(n_498), .B(n_521), .Y(n_717) );
AND2x2_ASAP7_75t_L g724 ( .A(n_498), .B(n_550), .Y(n_724) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g546 ( .A(n_499), .Y(n_546) );
BUFx3_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
AND2x2_ASAP7_75t_L g592 ( .A(n_499), .B(n_578), .Y(n_592) );
AND2x2_ASAP7_75t_L g655 ( .A(n_499), .B(n_514), .Y(n_655) );
AND2x2_ASAP7_75t_L g660 ( .A(n_499), .B(n_521), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_507), .B(n_510), .Y(n_501) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_513), .B(n_666), .Y(n_768) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
INVx2_ASAP7_75t_L g550 ( .A(n_514), .Y(n_550) );
OR2x2_ASAP7_75t_L g553 ( .A(n_514), .B(n_521), .Y(n_553) );
INVx2_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_514), .B(n_548), .Y(n_594) );
AND2x2_ASAP7_75t_L g667 ( .A(n_514), .B(n_521), .Y(n_667) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_533), .B(n_630), .Y(n_776) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g588 ( .A(n_534), .Y(n_588) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g568 ( .A(n_535), .Y(n_568) );
AND2x2_ASAP7_75t_L g574 ( .A(n_535), .B(n_556), .Y(n_574) );
INVx1_ASAP7_75t_L g622 ( .A(n_535), .Y(n_622) );
OR2x2_ASAP7_75t_L g627 ( .A(n_535), .B(n_606), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_535), .B(n_606), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_535), .B(n_605), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_535), .B(n_573), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_551), .B(n_554), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
OR2x2_ASAP7_75t_L g552 ( .A(n_545), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g703 ( .A(n_545), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g733 ( .A(n_545), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_546), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g701 ( .A(n_546), .Y(n_701) );
OR2x2_ASAP7_75t_L g614 ( .A(n_547), .B(n_615), .Y(n_614) );
INVxp33_ASAP7_75t_L g732 ( .A(n_547), .Y(n_732) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx2_ASAP7_75t_L g636 ( .A(n_548), .Y(n_636) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g590 ( .A(n_550), .Y(n_590) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_552), .A2(n_623), .B1(n_628), .B2(n_699), .C(n_702), .Y(n_698) );
OR2x2_ASAP7_75t_L g685 ( .A(n_553), .B(n_636), .Y(n_685) );
INVx2_ASAP7_75t_L g734 ( .A(n_553), .Y(n_734) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g634 ( .A(n_555), .Y(n_634) );
OR2x2_ASAP7_75t_L g637 ( .A(n_555), .B(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_555), .Y(n_678) );
OR2x2_ASAP7_75t_L g691 ( .A(n_555), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_568), .Y(n_555) );
NAND2x1p5_ASAP7_75t_SL g587 ( .A(n_556), .B(n_572), .Y(n_587) );
INVx3_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_556), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_556), .Y(n_625) );
AND2x2_ASAP7_75t_L g706 ( .A(n_556), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_556), .B(n_620), .Y(n_713) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B(n_567), .Y(n_558) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_574), .Y(n_569) );
AND2x2_ASAP7_75t_L g765 ( .A(n_570), .B(n_624), .Y(n_765) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g669 ( .A(n_572), .B(n_639), .Y(n_669) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g604 ( .A(n_573), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g630 ( .A(n_573), .B(n_606), .Y(n_630) );
AND2x4_ASAP7_75t_L g727 ( .A(n_574), .B(n_697), .Y(n_727) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g646 ( .A(n_579), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_580), .B(n_667), .Y(n_751) );
AND2x2_ASAP7_75t_L g758 ( .A(n_580), .B(n_718), .Y(n_758) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g683 ( .A(n_581), .Y(n_683) );
AOI321xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_596), .A3(n_612), .B1(n_613), .B2(n_616), .C(n_631), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_584), .B(n_593), .Y(n_583) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_589), .B(n_591), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_586), .A2(n_597), .B(n_600), .Y(n_596) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g695 ( .A(n_587), .B(n_627), .Y(n_695) );
INVx1_ASAP7_75t_L g687 ( .A(n_588), .Y(n_687) );
INVx2_ASAP7_75t_L g672 ( .A(n_589), .Y(n_672) );
OAI32xp33_ASAP7_75t_L g775 ( .A1(n_589), .A2(n_737), .A3(n_748), .B1(n_776), .B2(n_777), .Y(n_775) );
INVx1_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
INVx1_ASAP7_75t_L g640 ( .A(n_591), .Y(n_640) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_SL g728 ( .A(n_592), .B(n_635), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_593), .B(n_597), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_593), .A2(n_669), .B1(n_730), .B2(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g718 ( .A(n_594), .Y(n_718) );
INVx1_ASAP7_75t_L g615 ( .A(n_595), .Y(n_615) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g700 ( .A(n_599), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_600), .B(n_617), .C(n_623), .D(n_628), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVxp67_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
AND2x2_ASAP7_75t_L g721 ( .A(n_601), .B(n_630), .Y(n_721) );
OR2x2_ASAP7_75t_L g730 ( .A(n_601), .B(n_604), .Y(n_730) );
AND2x2_ASAP7_75t_L g754 ( .A(n_601), .B(n_626), .Y(n_754) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g668 ( .A(n_602), .B(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g675 ( .A(n_602), .B(n_622), .Y(n_675) );
INVx1_ASAP7_75t_L g739 ( .A(n_603), .Y(n_739) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g647 ( .A(n_604), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g697 ( .A(n_604), .Y(n_697) );
INVx1_ASAP7_75t_L g639 ( .A(n_605), .Y(n_639) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g620 ( .A(n_606), .Y(n_620) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x4_ASAP7_75t_L g633 ( .A(n_619), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g674 ( .A(n_619), .Y(n_674) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_621), .Y(n_738) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g629 ( .A(n_625), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g715 ( .A(n_627), .Y(n_715) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g692 ( .A(n_630), .Y(n_692) );
AND2x2_ASAP7_75t_L g735 ( .A(n_630), .B(n_675), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_635), .B(n_637), .C(n_640), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g746 ( .A(n_635), .B(n_724), .Y(n_746) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g650 ( .A(n_638), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B(n_656), .C(n_670), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_645), .A2(n_753), .B(n_756), .Y(n_752) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g666 ( .A(n_648), .Y(n_666) );
AND2x2_ASAP7_75t_L g726 ( .A(n_648), .B(n_723), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g745 ( .A(n_653), .Y(n_745) );
AND2x2_ASAP7_75t_L g771 ( .A(n_653), .B(n_734), .Y(n_771) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_654), .Y(n_659) );
INVx2_ASAP7_75t_L g710 ( .A(n_655), .Y(n_710) );
NAND2x1_ASAP7_75t_L g744 ( .A(n_655), .B(n_745), .Y(n_744) );
AOI33xp33_ASAP7_75t_L g762 ( .A1(n_655), .A2(n_675), .A3(n_713), .B1(n_723), .B2(n_755), .B3(n_836), .Y(n_762) );
OAI22xp33_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_661), .B1(n_664), .B2(n_668), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g689 ( .A(n_660), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_661), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
OR2x2_ASAP7_75t_L g774 ( .A(n_663), .B(n_708), .Y(n_774) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
OAI22xp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B1(n_676), .B2(n_677), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_674), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_674), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g696 ( .A(n_675), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g761 ( .A(n_675), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_740), .Y(n_679) );
NOR4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_698), .C(n_719), .D(n_736), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B1(n_688), .B2(n_691), .C(n_693), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_SL g736 ( .A1(n_682), .A2(n_737), .B(n_738), .C(n_739), .Y(n_736) );
NAND2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g769 ( .A(n_685), .Y(n_769) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_689), .A2(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x6_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_706), .C(n_709), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g748 ( .A(n_708), .B(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_708), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_714), .B2(n_716), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_722), .B(n_725), .C(n_731), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_723), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_775), .Y(n_770) );
INVx3_ASAP7_75t_L g778 ( .A(n_723), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_725) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g737 ( .A(n_734), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_763), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_752), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B(n_747), .C(n_750), .Y(n_742) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_746), .B(n_767), .C(n_769), .Y(n_766) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B(n_762), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_770), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g794 ( .A(n_780), .B(n_787), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_782), .B(n_786), .Y(n_791) );
INVxp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2x1_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g817 ( .A(n_789), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g802 ( .A(n_799), .Y(n_802) );
OAI21x1_ASAP7_75t_SL g800 ( .A1(n_801), .A2(n_803), .B(n_818), .Y(n_800) );
BUFx3_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_811), .Y(n_803) );
AOI21x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_808), .B(n_809), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_805), .Y(n_810) );
INVx5_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx8_ASAP7_75t_R g822 ( .A(n_813), .Y(n_822) );
AND2x6_ASAP7_75t_SL g813 ( .A(n_814), .B(n_817), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .Y(n_819) );
INVx4_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AND2x4_ASAP7_75t_L g824 ( .A(n_825), .B(n_829), .Y(n_824) );
AND2x2_ASAP7_75t_SL g834 ( .A(n_825), .B(n_829), .Y(n_834) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
NOR2x1p5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx6_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
endmodule