module real_jpeg_22218_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_0),
.A2(n_27),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_67),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_67),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_55),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_4),
.A2(n_16),
.B(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_4),
.B(n_153),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_31),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_60),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_27),
.B1(n_53),
.B2(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_177)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_10),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_90),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_27),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_63),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_63),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_13),
.A2(n_38),
.B1(n_50),
.B2(n_51),
.Y(n_82)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_31),
.A3(n_51),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_16),
.A2(n_50),
.B1(n_51),
.B2(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_16),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_80),
.Y(n_81)
);

BUFx3_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_99),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_68),
.B1(n_69),
.B2(n_98),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.C(n_56),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_24),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_25),
.B(n_34),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_26),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.CON(n_26),
.SN(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_30),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_30),
.B(n_33),
.C(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_28),
.A2(n_51),
.B(n_80),
.C(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_28),
.B(n_81),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_43),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_28),
.B(n_32),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_35),
.A2(n_39),
.B1(n_40),
.B2(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_36),
.B(n_143),
.Y(n_142)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_43),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_39),
.A2(n_40),
.B1(n_124),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_39),
.A2(n_127),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_39),
.A2(n_40),
.B1(n_159),
.B2(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_44),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_49),
.B1(n_54),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_46),
.A2(n_49),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_46),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_47),
.B(n_50),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_49),
.Y(n_153)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_65),
.B1(n_66),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_81),
.B1(n_89),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_81),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_78),
.A2(n_81),
.B1(n_135),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_78),
.A2(n_81),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_78),
.A2(n_81),
.B1(n_106),
.B2(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.C(n_103),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_100),
.B(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_102),
.B(n_103),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_110),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_218),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_214),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_203),
.B(n_213),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_182),
.B(n_202),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_161),
.B(n_181),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_147),
.B(n_160),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_136),
.B(n_146),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_141),
.B(n_145),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_157),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_170),
.B1(n_179),
.B2(n_180),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_167),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_171),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_184),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_196),
.B2(n_197),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_199),
.C(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_193),
.C(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_198),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);


endmodule