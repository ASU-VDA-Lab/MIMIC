module real_jpeg_5585_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_1),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_50),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_2),
.A2(n_50),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_2),
.A2(n_50),
.B1(n_152),
.B2(n_269),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_82),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_82),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_27),
.B1(n_82),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_4),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_6),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_6),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_22),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_36),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_22),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_22),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_71),
.B(n_223),
.C(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_10),
.B(n_256),
.C(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_10),
.B(n_93),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_176),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_107),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_212),
.B1(n_321),
.B2(n_322),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_211),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_177),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_177),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.C(n_160),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_18),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_51),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_19),
.B(n_52),
.C(n_95),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_47),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_25),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_22),
.A2(n_224),
.B(n_227),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_25),
.Y(n_132)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_28),
.B(n_48),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_35),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_36),
.B(n_197),
.Y(n_196)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_42),
.Y(n_207)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_44),
.Y(n_135)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_94),
.B1(n_95),
.B2(n_124),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_87),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_79),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_55),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_62),
.B2(n_66),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_58),
.Y(n_226)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_60),
.A2(n_128),
.A3(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_70),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_77),
.Y(n_70)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_72),
.Y(n_242)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_74),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_74),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_80),
.B(n_93),
.Y(n_162)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_87),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_88),
.B(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_118),
.B(n_119),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_97),
.B(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_97),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_97),
.B(n_186),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_103),
.B2(n_106),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_108),
.B1(n_110),
.B2(n_114),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_107),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_118),
.B(n_119),
.Y(n_239)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_125),
.A2(n_126),
.B1(n_160),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_139),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_127),
.B(n_139),
.Y(n_193)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_147),
.B(n_150),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_174),
.B(n_182),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_150),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_151),
.A2(n_169),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_151),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_164),
.B(n_205),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_168),
.B(n_282),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_172),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_174),
.B(n_267),
.Y(n_296)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_185),
.B(n_240),
.Y(n_272)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_212),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_246),
.B(n_320),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_214),
.B(n_217),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.C(n_236),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_218),
.B(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_221),
.A2(n_236),
.B1(n_237),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_222),
.A2(n_233),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_314),
.B(n_319),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_301),
.B(n_313),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_276),
.B(n_300),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_261),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_261),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_259),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_252),
.B1(n_259),
.B2(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_274),
.C(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_286),
.B(n_299),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_295),
.B(n_298),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_318),
.Y(n_319)
);


endmodule