module fake_jpeg_19708_n_206 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_50)
);

OR2x6_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_26),
.B1(n_12),
.B2(n_22),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_55),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_14),
.B1(n_11),
.B2(n_18),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_34),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_38),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_73),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_52),
.C(n_53),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_77),
.C(n_73),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_44),
.B(n_55),
.C(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_52),
.C(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_52),
.B1(n_47),
.B2(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_88),
.B1(n_58),
.B2(n_72),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_47),
.B1(n_50),
.B2(n_40),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_95),
.B1(n_48),
.B2(n_66),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_69),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_58),
.B1(n_64),
.B2(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_99),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_104),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_64),
.B1(n_42),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_66),
.B1(n_71),
.B2(n_48),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_64),
.B1(n_42),
.B2(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_74),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_105),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_64),
.A3(n_25),
.B1(n_70),
.B2(n_48),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_71),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_77),
.C(n_75),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_116),
.C(n_120),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_87),
.B(n_82),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_113),
.B(n_124),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_127),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_64),
.B1(n_84),
.B2(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_83),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_18),
.C(n_7),
.Y(n_114)
);

NOR2xp67_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_8),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_91),
.C(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_126),
.B1(n_35),
.B2(n_60),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_31),
.C(n_37),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_25),
.B(n_11),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_39),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_60),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_132),
.B1(n_140),
.B2(n_122),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_60),
.B1(n_23),
.B2(n_11),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_129),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_9),
.C(n_7),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_20),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_37),
.C(n_31),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_141),
.C(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_23),
.B1(n_31),
.B2(n_2),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_37),
.C(n_39),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_20),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_107),
.B1(n_123),
.B2(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_109),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_139),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_124),
.B1(n_111),
.B2(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_159),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_113),
.B(n_121),
.C(n_117),
.D(n_20),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_140),
.B(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_113),
.B1(n_9),
.B2(n_7),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_148),
.B1(n_158),
.B2(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_164),
.C(n_153),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_174),
.B(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_135),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_151),
.C(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_135),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_168),
.B(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_164),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_194),
.A3(n_0),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_144),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_160),
.B(n_1),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_194),
.B(n_2),
.C(n_3),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_37),
.C(n_54),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_198),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_54),
.A3(n_37),
.B1(n_13),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_54),
.A3(n_37),
.B1(n_13),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_0),
.B(n_3),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_196),
.C(n_13),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_200),
.C(n_5),
.Y(n_206)
);


endmodule