module fake_jpeg_28020_n_295 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_282;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_18),
.B(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_38),
.CON(n_72),
.SN(n_72)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_48),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_0),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_67),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_34),
.B1(n_29),
.B2(n_26),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_34),
.B1(n_26),
.B2(n_19),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_80),
.B(n_47),
.C(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_38),
.B1(n_19),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_82),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_31),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_36),
.B1(n_23),
.B2(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_37),
.B1(n_30),
.B2(n_23),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_35),
.B(n_22),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_20),
.C(n_44),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_43),
.B1(n_44),
.B2(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_96),
.B1(n_104),
.B2(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_109),
.B(n_112),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_20),
.B1(n_44),
.B2(n_35),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_73),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_113),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_43),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_115),
.Y(n_123)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_82),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_47),
.B(n_2),
.Y(n_109)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_65),
.B1(n_74),
.B2(n_58),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_3),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_65),
.B1(n_58),
.B2(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_135),
.B1(n_86),
.B2(n_108),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_85),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_64),
.B1(n_70),
.B2(n_54),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_144),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_56),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_114),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_118),
.B1(n_121),
.B2(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_7),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_11),
.C(n_12),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_101),
.C(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_85),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_166),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_158),
.B(n_171),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_154),
.B(n_162),
.Y(n_206)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_102),
.B1(n_103),
.B2(n_89),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_135),
.B1(n_124),
.B2(n_123),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_163),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_88),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_91),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_97),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_113),
.C(n_116),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_115),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_176),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_120),
.C(n_105),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_112),
.B(n_92),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_86),
.B1(n_138),
.B2(n_143),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_112),
.B(n_92),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_167),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_198),
.C(n_169),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_126),
.B1(n_134),
.B2(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_146),
.B1(n_136),
.B2(n_137),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_200),
.B1(n_167),
.B2(n_148),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_149),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_106),
.B1(n_148),
.B2(n_122),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_127),
.B(n_142),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_173),
.B(n_172),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_170),
.A2(n_124),
.B1(n_142),
.B2(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_157),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_90),
.B1(n_143),
.B2(n_13),
.C(n_14),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_156),
.Y(n_209)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_216),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_225),
.B1(n_189),
.B2(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_184),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_222),
.B(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_223),
.B1(n_228),
.B2(n_187),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_171),
.C(n_173),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_198),
.C(n_206),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_166),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_177),
.B1(n_174),
.B2(n_205),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_179),
.B(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_151),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_202),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_240),
.C(n_241),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_239),
.B(n_210),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_237),
.B1(n_243),
.B2(n_217),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_183),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_192),
.B1(n_151),
.B2(n_193),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_186),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_190),
.C(n_189),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_190),
.C(n_159),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_223),
.C(n_213),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_197),
.B1(n_187),
.B2(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_185),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_220),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_255),
.B1(n_219),
.B2(n_230),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_11),
.B(n_12),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_215),
.B(n_228),
.C(n_210),
.D(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_225),
.B1(n_226),
.B2(n_209),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_219),
.B1(n_147),
.B2(n_145),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_242),
.C(n_234),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_207),
.B1(n_212),
.B2(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.C(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_240),
.C(n_231),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_265),
.B1(n_269),
.B2(n_251),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_250),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_106),
.B1(n_105),
.B2(n_110),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_255),
.B1(n_246),
.B2(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_259),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_274),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_278),
.C(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_249),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_264),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_276),
.B1(n_262),
.B2(n_258),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_282),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_258),
.B1(n_106),
.B2(n_13),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_280),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_280),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_12),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_13),
.Y(n_295)
);


endmodule