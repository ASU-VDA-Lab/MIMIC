module real_jpeg_23257_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_1),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_28),
.B(n_43),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_94),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_1),
.A2(n_25),
.B1(n_182),
.B2(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_62),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_81),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_2),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_155),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_77),
.B1(n_78),
.B2(n_155),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_164),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_164),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_4),
.A2(n_67),
.B1(n_77),
.B2(n_164),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_7),
.A2(n_35),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_7),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_52),
.B1(n_77),
.B2(n_80),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_152),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_13),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_88),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_73),
.B1(n_74),
.B2(n_88),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_88),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_69),
.B1(n_77),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_14),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_116),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_116),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_116),
.Y(n_261)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_20),
.B(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_103),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_21),
.A2(n_83),
.B1(n_84),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_21),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_53),
.B2(n_82),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_54),
.B(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_24),
.A2(n_36),
.B1(n_54),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_25),
.A2(n_109),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_25),
.A2(n_172),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_33),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_25),
.A2(n_211),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_26),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_26),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_26),
.A2(n_248),
.B1(n_249),
.B2(n_252),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_27),
.B(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_31),
.B(n_152),
.Y(n_189)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_32),
.A2(n_107),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_34),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_47),
.B(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_37),
.A2(n_46),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_37),
.A2(n_97),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_38),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_38),
.A2(n_98),
.B(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_38),
.A2(n_99),
.B1(n_154),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_38),
.A2(n_99),
.B1(n_163),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_38),
.A2(n_50),
.B(n_98),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_41),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_40),
.B(n_92),
.Y(n_209)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_41),
.A2(n_45),
.B(n_152),
.C(n_157),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_41),
.A2(n_62),
.A3(n_91),
.B1(n_200),
.B2(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_46),
.B(n_152),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_46),
.A2(n_100),
.B(n_113),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_70),
.B(n_75),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_115),
.B(n_117),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_57),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_57),
.A2(n_58),
.B1(n_115),
.B2(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_58),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_59),
.A2(n_63),
.A3(n_73),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_60),
.B(n_62),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_63),
.B1(n_91),
.B2(n_92),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_63),
.B(n_152),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_81),
.Y(n_117)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_128),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_77),
.A2(n_152),
.B(n_245),
.Y(n_264)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_81),
.A2(n_128),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_81),
.A2(n_128),
.B1(n_265),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_96),
.B(n_102),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_96),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_90),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_95),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_89),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_89),
.A2(n_94),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_89),
.A2(n_94),
.B1(n_224),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_89),
.A2(n_261),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_90),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_90),
.B(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_120),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_123),
.B1(n_137),
.B2(n_138),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_103),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.C(n_118),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_104),
.A2(n_105),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_106),
.B(n_112),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_108),
.B(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_114),
.B(n_118),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_139),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_136),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_134),
.A2(n_201),
.B(n_276),
.Y(n_291)
);

AOI311xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_300),
.A3(n_312),
.B(n_316),
.C(n_317),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_267),
.C(n_295),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_239),
.B(n_266),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_217),
.B(n_238),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_193),
.B(n_216),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_168),
.B(n_192),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_158),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_150),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_165),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_165),
.C(n_166),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_178),
.B(n_191),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_176),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_185),
.B(n_190),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_207),
.B1(n_214),
.B2(n_215),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_206),
.C(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_231),
.B2(n_232),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_234),
.C(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_241),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_258),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_257),
.C(n_258),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_253),
.B2(n_254),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_253),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_268),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_285),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_269),
.B(n_285),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_280),
.C(n_281),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_271),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_281),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_284),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_285),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_293),
.CI(n_294),
.CON(n_285),
.SN(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_313),
.B(n_318),
.C(n_321),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_309),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_308),
.Y(n_302)
);

FAx1_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_306),
.CI(n_308),
.CON(n_315),
.SN(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_315),
.Y(n_322)
);


endmodule