module fake_jpeg_30390_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_23),
.B1(n_43),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_63),
.B1(n_65),
.B2(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_48),
.B1(n_65),
.B2(n_63),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_107),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_61),
.B(n_49),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_105),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_87),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_66),
.B1(n_61),
.B2(n_49),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_89),
.B1(n_84),
.B2(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_66),
.B1(n_54),
.B2(n_57),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_47),
.B(n_64),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_56),
.B(n_79),
.C(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_70),
.B(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_59),
.B1(n_53),
.B2(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_62),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_100),
.A3(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_2),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_5),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_5),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_128),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_28),
.A3(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_19),
.C(n_24),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_17),
.C(n_18),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_127),
.B(n_34),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_144),
.C(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_143),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_155),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_137),
.C(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_159),
.A3(n_138),
.B1(n_145),
.B2(n_141),
.C1(n_156),
.C2(n_150),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_155),
.B(n_152),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_139),
.B(n_136),
.C(n_36),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_32),
.Y(n_168)
);


endmodule