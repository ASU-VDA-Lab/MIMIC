module fake_ariane_907_n_1829 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1829);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1829;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1803;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_21),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_61),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_1),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_72),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_59),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_76),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

INVx4_ASAP7_75t_R g179 ( 
.A(n_54),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_71),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_53),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_40),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_15),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_31),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_42),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_17),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_80),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_81),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_6),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_147),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_69),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_7),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_100),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_95),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_28),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_79),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_113),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_93),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_132),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_90),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_21),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_17),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_20),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_110),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_29),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_60),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_57),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_151),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_0),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_32),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_2),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_116),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_32),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_13),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_135),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_130),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_49),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_46),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_26),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_29),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_45),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_115),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_84),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_51),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_31),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_142),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_73),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_37),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_70),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_101),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_62),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_124),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_19),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_48),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_112),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_77),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_96),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_127),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_105),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_25),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_114),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_11),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_45),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_50),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_117),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_62),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_41),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_44),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_98),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_104),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_128),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_12),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_51),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_74),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_49),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_33),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_107),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_43),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_123),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_121),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_94),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_86),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_24),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_28),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_108),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_14),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_1),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_38),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_7),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_66),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_41),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_30),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_173),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_173),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_173),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_281),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_173),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_251),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_244),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_242),
.B(n_0),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_281),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_166),
.Y(n_351)
);

BUFx6f_ASAP7_75t_SL g352 ( 
.A(n_267),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_337),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_253),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_259),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_239),
.B(n_2),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_186),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_264),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_286),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_203),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_169),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_207),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_207),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_242),
.B(n_3),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_218),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_168),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_292),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_292),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_167),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_220),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_188),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_227),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_182),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_273),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_230),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_185),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_193),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_198),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_236),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_237),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_258),
.B(n_3),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_221),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_221),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_187),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_238),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_243),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_245),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_277),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_250),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_255),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_271),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_246),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_247),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_278),
.B(n_5),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_285),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_287),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_291),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_302),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_310),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_307),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_168),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_249),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_189),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_254),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_195),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_318),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_196),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_256),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_364),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_377),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_373),
.B(n_233),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_232),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_360),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_380),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g446 ( 
.A(n_369),
.B(n_336),
.C(n_191),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_205),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_351),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_354),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_299),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_362),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_356),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_363),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_366),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_346),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_371),
.B(n_175),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_357),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_370),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_371),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_205),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_399),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_352),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_376),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_420),
.B(n_210),
.Y(n_470)
);

CKINVDCx8_ASAP7_75t_R g471 ( 
.A(n_355),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_352),
.B(n_210),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_422),
.Y(n_485)
);

AND3x2_ASAP7_75t_L g486 ( 
.A(n_382),
.B(n_202),
.C(n_197),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_359),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_359),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_365),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_378),
.B(n_267),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_412),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_421),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_365),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_383),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_386),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_368),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_438),
.B(n_352),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_428),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_480),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_361),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_428),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_472),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

INVx4_ASAP7_75t_SL g510 ( 
.A(n_470),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_480),
.B(n_414),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_438),
.B(n_342),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_435),
.B(n_388),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_389),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_427),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_472),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_397),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_403),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_456),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_485),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_446),
.B(n_404),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_433),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_466),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_446),
.A2(n_358),
.B1(n_348),
.B2(n_405),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_415),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_466),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_453),
.B(n_447),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_458),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_447),
.B(n_419),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_470),
.A2(n_447),
.B1(n_465),
.B2(n_405),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_181),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_488),
.B(n_423),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_447),
.A2(n_390),
.B1(n_172),
.B2(n_309),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_488),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_472),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_484),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_451),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_350),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_464),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_484),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_457),
.A2(n_178),
.B1(n_191),
.B2(n_252),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_208),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_448),
.Y(n_560)
);

OAI21xp33_ASAP7_75t_SL g561 ( 
.A1(n_473),
.A2(n_398),
.B(n_396),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_443),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_473),
.Y(n_565)
);

INVx4_ASAP7_75t_SL g566 ( 
.A(n_426),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_465),
.B(n_374),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_469),
.A2(n_334),
.B1(n_290),
.B2(n_294),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_498),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_465),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_426),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_468),
.B(n_170),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_465),
.B(n_375),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_468),
.B(n_170),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_452),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_379),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_429),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_426),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_381),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_496),
.B(n_178),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_439),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_460),
.A2(n_490),
.B1(n_494),
.B2(n_489),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_429),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_471),
.B(n_171),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_460),
.B(n_290),
.C(n_252),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_471),
.B(n_171),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_454),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_479),
.A2(n_260),
.B1(n_262),
.B2(n_265),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_479),
.B(n_396),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_475),
.B(n_398),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_477),
.B(n_181),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_467),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_489),
.A2(n_384),
.B1(n_385),
.B2(n_299),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_430),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_477),
.B(n_400),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_500),
.B(n_400),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_401),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_492),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_430),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_444),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_444),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_481),
.B(n_401),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_445),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_481),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_483),
.B(n_402),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_490),
.B(n_402),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_445),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_449),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_434),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_494),
.B(n_418),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_434),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_483),
.B(n_174),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_495),
.A2(n_293),
.B1(n_267),
.B2(n_413),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_476),
.B(n_406),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_434),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_495),
.B(n_406),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_493),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_486),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_459),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_497),
.B(n_174),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_497),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_450),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_476),
.B(n_407),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_437),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_499),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_499),
.B(n_407),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_459),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_500),
.B(n_418),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_476),
.B(n_408),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_450),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_487),
.A2(n_293),
.B1(n_413),
.B2(n_411),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_426),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_487),
.B(n_408),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_437),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_461),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_461),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_487),
.B(n_211),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_462),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_462),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_486),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_437),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_426),
.Y(n_649)
);

CKINVDCx14_ASAP7_75t_R g650 ( 
.A(n_426),
.Y(n_650)
);

AND2x2_ASAP7_75t_SL g651 ( 
.A(n_431),
.B(n_214),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_209),
.Y(n_652)
);

NOR3x1_ASAP7_75t_L g653 ( 
.A(n_557),
.B(n_410),
.C(n_409),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_539),
.B(n_241),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_536),
.B(n_268),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_501),
.B(n_303),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_513),
.B(n_269),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_506),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_634),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_634),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_544),
.B(n_322),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_504),
.Y(n_664)
);

O2A1O1Ixp5_ASAP7_75t_L g665 ( 
.A1(n_571),
.A2(n_225),
.B(n_275),
.C(n_263),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_514),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_572),
.B(n_176),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_571),
.B(n_176),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_504),
.B(n_409),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_513),
.B(n_270),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_572),
.B(n_177),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_529),
.A2(n_311),
.B1(n_320),
.B2(n_317),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_571),
.B(n_177),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_515),
.B(n_521),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_570),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_541),
.B(n_519),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_528),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_535),
.A2(n_305),
.B(n_304),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_548),
.B(n_180),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_567),
.B(n_272),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_592),
.B(n_283),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_503),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_511),
.B(n_410),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_556),
.B(n_180),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_601),
.B(n_190),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_579),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_592),
.B(n_321),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_560),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_570),
.B(n_411),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_527),
.B(n_549),
.Y(n_692)
);

OAI221xp5_ASAP7_75t_L g693 ( 
.A1(n_619),
.A2(n_306),
.B1(n_317),
.B2(n_336),
.C(n_311),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_644),
.A2(n_293),
.B1(n_441),
.B2(n_455),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_510),
.B(n_416),
.Y(n_695)
);

NOR2x1p5_ASAP7_75t_L g696 ( 
.A(n_505),
.B(n_316),
.Y(n_696)
);

BUFx2_ASAP7_75t_SL g697 ( 
.A(n_523),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_533),
.A2(n_455),
.B(n_441),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_509),
.B(n_316),
.C(n_332),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_644),
.A2(n_455),
.B1(n_441),
.B2(n_332),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_542),
.A2(n_333),
.B1(n_334),
.B2(n_179),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_530),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_510),
.A2(n_416),
.B1(n_216),
.B2(n_219),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_601),
.B(n_190),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_510),
.B(n_192),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_602),
.A2(n_616),
.B1(n_632),
.B2(n_610),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_511),
.B(n_333),
.C(n_288),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_523),
.B(n_431),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_558),
.B(n_192),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_533),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_523),
.B(n_199),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_610),
.B(n_199),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_564),
.B(n_431),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_632),
.B(n_288),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_538),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_592),
.B(n_301),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_585),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_651),
.A2(n_279),
.B1(n_248),
.B2(n_231),
.Y(n_718)
);

BUFx4_ASAP7_75t_L g719 ( 
.A(n_517),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_558),
.B(n_301),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_651),
.B(n_308),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_549),
.B(n_308),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_538),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_562),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_585),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_312),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_518),
.B(n_312),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_553),
.B(n_313),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_553),
.B(n_313),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_583),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_518),
.B(n_314),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_584),
.B(n_314),
.Y(n_732)
);

AND2x4_ASAP7_75t_SL g733 ( 
.A(n_564),
.B(n_215),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_597),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_564),
.B(n_431),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_503),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_518),
.B(n_315),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_607),
.Y(n_741)
);

OAI221xp5_ASAP7_75t_L g742 ( 
.A1(n_545),
.A2(n_224),
.B1(n_226),
.B2(n_297),
.C(n_228),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_602),
.B(n_315),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_602),
.B(n_335),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_602),
.B(n_335),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_542),
.A2(n_229),
.B1(n_295),
.B2(n_325),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_607),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_518),
.B(n_296),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_609),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_609),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_612),
.B(n_200),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_577),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_590),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_518),
.B(n_552),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_616),
.B(n_298),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_505),
.B(n_591),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_616),
.B(n_5),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_577),
.B(n_436),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_552),
.B(n_184),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_612),
.B(n_201),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_613),
.A2(n_436),
.B(n_431),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_542),
.A2(n_436),
.B1(n_431),
.B2(n_181),
.Y(n_762)
);

INVx8_ASAP7_75t_L g763 ( 
.A(n_616),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_622),
.B(n_204),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_8),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_613),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_568),
.B(n_206),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_561),
.A2(n_436),
.B(n_330),
.C(n_327),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_590),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_599),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_633),
.B(n_212),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_588),
.B(n_436),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_635),
.B(n_213),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_507),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_599),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_542),
.A2(n_261),
.B1(n_324),
.B2(n_319),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_532),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_605),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_614),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_578),
.A2(n_257),
.B1(n_284),
.B2(n_282),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_605),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_586),
.B(n_14),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_502),
.B(n_184),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_581),
.A2(n_234),
.B1(n_280),
.B2(n_222),
.Y(n_785)
);

BUFx6f_ASAP7_75t_SL g786 ( 
.A(n_624),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_589),
.B(n_15),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_633),
.B(n_274),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_552),
.B(n_563),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_625),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_625),
.Y(n_791)
);

O2A1O1Ixp5_ASAP7_75t_L g792 ( 
.A1(n_618),
.A2(n_436),
.B(n_266),
.C(n_240),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_627),
.B(n_16),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_615),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_629),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_524),
.B(n_223),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_647),
.B(n_194),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_647),
.B(n_604),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_507),
.B(n_16),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_623),
.B(n_18),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_525),
.B(n_276),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_SL g802 ( 
.A(n_626),
.B(n_194),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_600),
.A2(n_276),
.B1(n_184),
.B2(n_194),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_531),
.B(n_19),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_624),
.B(n_22),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_531),
.B(n_532),
.Y(n_806)
);

NAND2x1_ASAP7_75t_L g807 ( 
.A(n_639),
.B(n_194),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_615),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_629),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_637),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_617),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_546),
.B(n_276),
.Y(n_812)
);

NOR2x1p5_ASAP7_75t_L g813 ( 
.A(n_635),
.B(n_181),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_552),
.B(n_276),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_637),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_531),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_677),
.A2(n_574),
.B1(n_576),
.B2(n_650),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_677),
.B(n_626),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_675),
.B(n_551),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_675),
.B(n_554),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_654),
.B(n_565),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_763),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_663),
.B(n_582),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_652),
.A2(n_563),
.B1(n_628),
.B2(n_569),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_660),
.B(n_662),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_789),
.A2(n_502),
.B(n_559),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_587),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_706),
.B(n_624),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_659),
.B(n_563),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_709),
.A2(n_646),
.B(n_645),
.C(n_611),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_789),
.A2(n_559),
.B(n_550),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_661),
.B(n_645),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_676),
.B(n_537),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_666),
.B(n_646),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_664),
.B(n_598),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_754),
.A2(n_526),
.B(n_520),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_678),
.B(n_520),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_754),
.A2(n_522),
.B(n_550),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_669),
.A2(n_522),
.B(n_526),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_688),
.B(n_582),
.Y(n_842)
);

BUFx5_ASAP7_75t_L g843 ( 
.A(n_695),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_761),
.A2(n_540),
.B(n_642),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_669),
.A2(n_674),
.B(n_806),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_736),
.B(n_537),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_684),
.B(n_593),
.Y(n_847)
);

OAI21xp33_ASAP7_75t_L g848 ( 
.A1(n_656),
.A2(n_643),
.B(n_595),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_658),
.B(n_534),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_587),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_658),
.B(n_640),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_756),
.B(n_638),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_710),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_698),
.A2(n_540),
.B(n_512),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_763),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_674),
.A2(n_555),
.B(n_508),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_752),
.B(n_603),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_806),
.A2(n_508),
.B(n_547),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_671),
.B(n_608),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_763),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_759),
.A2(n_631),
.B(n_648),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_671),
.B(n_594),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_673),
.B(n_630),
.C(n_636),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_716),
.A2(n_547),
.B(n_555),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_715),
.A2(n_508),
.B1(n_555),
.B2(n_547),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_695),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_723),
.B(n_617),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_730),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_665),
.A2(n_512),
.B(n_648),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_691),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_690),
.B(n_639),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_734),
.B(n_621),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_735),
.B(n_621),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_692),
.B(n_691),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_724),
.B(n_620),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_716),
.A2(n_512),
.B(n_639),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_682),
.A2(n_552),
.B(n_641),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_739),
.A2(n_741),
.B1(n_815),
.B2(n_810),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_719),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_747),
.B(n_641),
.Y(n_880)
);

AOI21x1_ASAP7_75t_L g881 ( 
.A1(n_759),
.A2(n_631),
.B(n_566),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_749),
.B(n_543),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_682),
.A2(n_649),
.B(n_573),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_656),
.B(n_649),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_750),
.B(n_543),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_743),
.A2(n_543),
.B1(n_649),
.B2(n_580),
.Y(n_886)
);

CKINVDCx10_ASAP7_75t_R g887 ( 
.A(n_786),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_782),
.A2(n_649),
.B(n_580),
.C(n_573),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_766),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_689),
.A2(n_649),
.B(n_573),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_743),
.B(n_580),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_689),
.A2(n_580),
.B(n_573),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_695),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_773),
.B(n_566),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_680),
.A2(n_580),
.B(n_573),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_779),
.A2(n_795),
.B1(n_791),
.B2(n_790),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_670),
.B(n_543),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_685),
.A2(n_194),
.B(n_181),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_777),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_784),
.B(n_543),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_809),
.A2(n_566),
.B(n_596),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_765),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_814),
.A2(n_596),
.B(n_276),
.Y(n_903)
);

AO32x1_ASAP7_75t_L g904 ( 
.A1(n_687),
.A2(n_596),
.A3(n_276),
.B1(n_184),
.B2(n_35),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_755),
.B(n_596),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_801),
.A2(n_276),
.B(n_184),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_777),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_812),
.A2(n_184),
.B(n_78),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_755),
.B(n_184),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_657),
.B(n_27),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_802),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_814),
.A2(n_184),
.B(n_82),
.Y(n_912)
);

AO22x1_ASAP7_75t_L g913 ( 
.A1(n_757),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_765),
.B(n_36),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_738),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_733),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_697),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_744),
.B(n_36),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_798),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_765),
.A2(n_718),
.B1(n_757),
.B2(n_744),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_774),
.A2(n_91),
.B(n_163),
.Y(n_921)
);

O2A1O1Ixp5_ASAP7_75t_L g922 ( 
.A1(n_709),
.A2(n_38),
.B(n_39),
.C(n_42),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_774),
.A2(n_119),
.B(n_158),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_717),
.B(n_43),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_753),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_725),
.B(n_753),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_745),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_745),
.B(n_48),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_769),
.B(n_52),
.Y(n_929)
);

AND2x6_ASAP7_75t_SL g930 ( 
.A(n_782),
.B(n_53),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_786),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_707),
.B(n_54),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_733),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_681),
.B(n_55),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_681),
.B(n_55),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_655),
.B(n_56),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_769),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_758),
.B(n_57),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_58),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_729),
.B(n_58),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_679),
.B(n_65),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_738),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_751),
.B(n_122),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_787),
.A2(n_125),
.B(n_126),
.C(n_131),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_787),
.B(n_133),
.C(n_134),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_770),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_760),
.B(n_139),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_777),
.B(n_722),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_800),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_767),
.B(n_165),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_805),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_738),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_770),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_764),
.B(n_788),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_720),
.A2(n_704),
.B(n_714),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_771),
.B(n_726),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_727),
.A2(n_740),
.B(n_731),
.C(n_792),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_686),
.A2(n_712),
.B(n_668),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_672),
.A2(n_796),
.B(n_727),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_777),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_775),
.B(n_808),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_797),
.B(n_693),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_793),
.A2(n_721),
.B(n_699),
.C(n_711),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_721),
.A2(n_701),
.B1(n_793),
.B2(n_776),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_778),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_762),
.A2(n_746),
.B1(n_816),
.B2(n_683),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_696),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_742),
.B(n_740),
.C(n_731),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_683),
.A2(n_799),
.B1(n_804),
.B2(n_694),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_732),
.B(n_785),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_781),
.A2(n_808),
.B(n_811),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_708),
.A2(n_737),
.B1(n_713),
.B2(n_703),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_703),
.A2(n_780),
.B1(n_813),
.B2(n_705),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_781),
.A2(n_811),
.B(n_794),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_799),
.A2(n_804),
.B(n_705),
.C(n_807),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_794),
.A2(n_783),
.B(n_738),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_748),
.A2(n_772),
.B(n_700),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_703),
.B(n_653),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_748),
.B(n_803),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_789),
.A2(n_754),
.B(n_674),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_677),
.B(n_570),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_654),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_654),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_789),
.A2(n_754),
.B(n_674),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_677),
.B(n_570),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_677),
.B(n_570),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_654),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_789),
.A2(n_754),
.B(n_674),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_763),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_677),
.B(n_360),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_971),
.A2(n_974),
.B(n_890),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_989),
.B(n_823),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_908),
.A2(n_888),
.B(n_844),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_883),
.A2(n_892),
.B(n_877),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_931),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_820),
.A2(n_821),
.B(n_859),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_836),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_838),
.A2(n_840),
.B(n_980),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_853),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_989),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_990),
.A2(n_970),
.B(n_819),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_823),
.B(n_860),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_931),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_831),
.A2(n_956),
.B(n_954),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_868),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_847),
.B(n_824),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_887),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_849),
.A2(n_845),
.B(n_862),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_981),
.B(n_985),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_866),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_918),
.A2(n_928),
.B(n_910),
.C(n_964),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_958),
.A2(n_884),
.B(n_969),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_984),
.A2(n_988),
.B(n_832),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_959),
.A2(n_975),
.B(n_947),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_827),
.A2(n_854),
.B(n_841),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_895),
.A2(n_976),
.B(n_864),
.Y(n_1017)
);

AOI21x1_ASAP7_75t_L g1018 ( 
.A1(n_909),
.A2(n_977),
.B(n_891),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_957),
.A2(n_935),
.B(n_934),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_889),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_823),
.B(n_860),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_901),
.A2(n_869),
.B(n_903),
.Y(n_1022)
);

AO31x2_ASAP7_75t_L g1023 ( 
.A1(n_941),
.A2(n_896),
.A3(n_878),
.B(n_979),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_963),
.A2(n_920),
.B(n_932),
.C(n_950),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_830),
.A2(n_835),
.B(n_833),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_856),
.A2(n_858),
.B(n_876),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_962),
.A2(n_842),
.B1(n_874),
.B2(n_846),
.Y(n_1027)
);

AO21x1_ASAP7_75t_L g1028 ( 
.A1(n_909),
.A2(n_912),
.B(n_968),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_986),
.B(n_852),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_911),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_982),
.B(n_987),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_830),
.A2(n_825),
.B(n_936),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_943),
.A2(n_848),
.B(n_822),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_983),
.B(n_897),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_870),
.B(n_978),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_822),
.A2(n_872),
.B(n_880),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_914),
.A2(n_940),
.B1(n_939),
.B2(n_972),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_850),
.B(n_951),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_817),
.B(n_875),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_924),
.A2(n_929),
.A3(n_966),
.B(n_898),
.Y(n_1041)
);

OA22x2_ASAP7_75t_L g1042 ( 
.A1(n_973),
.A2(n_879),
.B1(n_916),
.B2(n_837),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_867),
.A2(n_880),
.B(n_873),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_850),
.B(n_828),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_866),
.B(n_893),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_925),
.A2(n_961),
.B(n_926),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_924),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_867),
.A2(n_873),
.B(n_872),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_857),
.B(n_843),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_914),
.A2(n_839),
.B1(n_871),
.B2(n_893),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_SL g1051 ( 
.A1(n_927),
.A2(n_902),
.B(n_826),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_949),
.B(n_933),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_839),
.A2(n_865),
.B(n_882),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_944),
.A2(n_863),
.B(n_922),
.C(n_945),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_929),
.A2(n_923),
.B(n_921),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_SL g1056 ( 
.A1(n_882),
.A2(n_885),
.B(n_900),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_919),
.B(n_967),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_885),
.A2(n_900),
.B(n_938),
.Y(n_1058)
);

AND2x2_ASAP7_75t_SL g1059 ( 
.A(n_978),
.B(n_894),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_828),
.A2(n_886),
.B1(n_829),
.B2(n_905),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_894),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_937),
.A2(n_953),
.B(n_965),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_SL g1063 ( 
.A(n_915),
.B(n_952),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_855),
.B(n_960),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_843),
.B(n_855),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_915),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_946),
.A2(n_948),
.B(n_834),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_843),
.B(n_952),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_915),
.A2(n_952),
.B(n_942),
.C(n_913),
.Y(n_1069)
);

OAI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_930),
.A2(n_960),
.B1(n_899),
.B2(n_907),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_904),
.A2(n_942),
.B(n_899),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_904),
.A2(n_907),
.B(n_843),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_990),
.B(n_820),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_851),
.A2(n_831),
.B(n_821),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_819),
.B(n_530),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_990),
.B(n_820),
.Y(n_1076)
);

AOI21xp33_ASAP7_75t_L g1077 ( 
.A1(n_990),
.A2(n_663),
.B(n_970),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_990),
.B(n_820),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_836),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_990),
.B(n_820),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_819),
.B(n_664),
.Y(n_1083)
);

AOI221x1_ASAP7_75t_L g1084 ( 
.A1(n_918),
.A2(n_928),
.B1(n_920),
.B2(n_968),
.C(n_969),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_851),
.A2(n_831),
.B(n_821),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_906),
.A2(n_861),
.B(n_881),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_990),
.B(n_820),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_990),
.B(n_820),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_990),
.B(n_820),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_990),
.A2(n_928),
.B(n_918),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_817),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_887),
.Y(n_1097)
);

OAI222xp33_ASAP7_75t_L g1098 ( 
.A1(n_920),
.A2(n_964),
.B1(n_701),
.B2(n_746),
.C1(n_973),
.C2(n_776),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_819),
.B(n_664),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_990),
.A2(n_819),
.B1(n_928),
.B2(n_918),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_851),
.A2(n_831),
.B(n_821),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_836),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_879),
.B(n_763),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_970),
.A2(n_918),
.B(n_928),
.C(n_824),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_845),
.A2(n_861),
.B(n_883),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_836),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_990),
.B(n_660),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_906),
.A2(n_908),
.B(n_888),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_817),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_820),
.A2(n_821),
.B(n_851),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_990),
.B(n_820),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_823),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_990),
.B(n_820),
.Y(n_1115)
);

NAND2x1p5_ASAP7_75t_L g1116 ( 
.A(n_866),
.B(n_893),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_851),
.A2(n_831),
.B(n_821),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_989),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_970),
.A2(n_918),
.B(n_928),
.C(n_824),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_888),
.A2(n_969),
.A3(n_768),
.B(n_955),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_990),
.B(n_820),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_SL g1122 ( 
.A1(n_955),
.A2(n_706),
.B(n_833),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_990),
.A2(n_663),
.B(n_970),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_817),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_990),
.B(n_820),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_990),
.B(n_820),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_918),
.A2(n_928),
.B(n_969),
.C(n_935),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_845),
.A2(n_861),
.B(n_883),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_931),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_906),
.A2(n_861),
.B(n_881),
.Y(n_1130)
);

CKINVDCx8_ASAP7_75t_R g1131 ( 
.A(n_887),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_851),
.A2(n_820),
.B1(n_821),
.B2(n_920),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_998),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1035),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1100),
.B(n_1002),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1013),
.A2(n_1012),
.B(n_1127),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_1098),
.B(n_1024),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_1008),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1000),
.Y(n_1140)
);

AND2x6_ASAP7_75t_L g1141 ( 
.A(n_1011),
.B(n_993),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_993),
.B(n_1003),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1077),
.B(n_1123),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1083),
.B(n_1099),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1013),
.A2(n_1127),
.B(n_997),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1020),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_SL g1148 ( 
.A1(n_1042),
.A2(n_1007),
.B1(n_1081),
.B2(n_1078),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1003),
.B(n_1021),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_997),
.A2(n_1079),
.B(n_992),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1080),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1087),
.A2(n_1088),
.B1(n_1126),
.B2(n_1125),
.C(n_1090),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1113),
.A2(n_1121),
.B(n_1115),
.C(n_1132),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1068),
.B(n_1066),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1124),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1040),
.B(n_1110),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1035),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_992),
.B(n_1079),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1021),
.B(n_1045),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_996),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1102),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1114),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1082),
.B(n_1089),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1106),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1027),
.B(n_1082),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1061),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1089),
.A2(n_1096),
.B(n_1091),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1045),
.B(n_1044),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1038),
.A2(n_1042),
.B(n_1028),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1091),
.A2(n_1095),
.B(n_1094),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1075),
.A2(n_1029),
.B1(n_1036),
.B2(n_1059),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1110),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1045),
.B(n_1103),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1039),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1031),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1093),
.B(n_1030),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1084),
.A2(n_1095),
.B(n_1111),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1103),
.B(n_1001),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1093),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1052),
.B(n_1057),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1094),
.B(n_1096),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1051),
.A2(n_1111),
.B1(n_1109),
.B2(n_1112),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1009),
.A2(n_1033),
.B(n_1037),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1033),
.A2(n_1037),
.B(n_1015),
.Y(n_1186)
);

INVx3_ASAP7_75t_SL g1187 ( 
.A(n_1097),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_1059),
.B1(n_1098),
.B2(n_1047),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1107),
.B(n_1010),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1103),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1010),
.B(n_1025),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1114),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1060),
.A2(n_1034),
.B1(n_1050),
.B2(n_1070),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1005),
.A2(n_1019),
.B(n_1032),
.C(n_1054),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1070),
.B(n_1011),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1131),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1074),
.A2(n_1117),
.B(n_1101),
.C(n_1085),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1001),
.B(n_1118),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_L g1199 ( 
.A(n_1116),
.B(n_1118),
.Y(n_1199)
);

OAI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_1015),
.A2(n_1069),
.B(n_1053),
.Y(n_1200)
);

OAI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1058),
.A2(n_1049),
.B1(n_1053),
.B2(n_1129),
.C(n_1004),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1066),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_994),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_R g1204 ( 
.A(n_1065),
.B(n_1018),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_994),
.Y(n_1205)
);

BUFx4_ASAP7_75t_SL g1206 ( 
.A(n_1063),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1116),
.B(n_1023),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1064),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1058),
.A2(n_1072),
.B(n_1071),
.C(n_1067),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1023),
.B(n_1064),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1062),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1055),
.A2(n_1122),
.B(n_1017),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1023),
.B(n_1046),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1056),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1072),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1026),
.A2(n_1108),
.B(n_995),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1071),
.B(n_1041),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1108),
.A2(n_999),
.B(n_1016),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1120),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1014),
.A2(n_991),
.B(n_1130),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1022),
.A2(n_1086),
.B1(n_1041),
.B2(n_1120),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_1128),
.B(n_1105),
.Y(n_1222)
);

CKINVDCx6p67_ASAP7_75t_R g1223 ( 
.A(n_996),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_1104),
.B(n_1119),
.C(n_1012),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1083),
.B(n_819),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_993),
.B(n_989),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1110),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1100),
.B(n_1002),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1035),
.B(n_989),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_998),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_998),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1002),
.A2(n_1119),
.B(n_1104),
.C(n_1092),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_993),
.B(n_989),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_998),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_993),
.B(n_989),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1035),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_998),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1092),
.A2(n_1104),
.B(n_1119),
.C(n_1012),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1103),
.B(n_763),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1100),
.B(n_1002),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_998),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_998),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1008),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1100),
.B(n_1002),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1100),
.A2(n_1104),
.B1(n_1119),
.B2(n_1092),
.Y(n_1249)
);

INVx3_ASAP7_75t_SL g1250 ( 
.A(n_1008),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1019),
.A2(n_675),
.B(n_516),
.C(n_1100),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_998),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1008),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_1119),
.B(n_1092),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1092),
.A2(n_1100),
.B1(n_819),
.B2(n_920),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1008),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1100),
.A2(n_990),
.B1(n_1076),
.B2(n_1073),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1035),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_996),
.Y(n_1260)
);

AND2x6_ASAP7_75t_L g1261 ( 
.A(n_1011),
.B(n_823),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1035),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1131),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1083),
.B(n_819),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1266)
);

OAI21xp33_ASAP7_75t_L g1267 ( 
.A1(n_1092),
.A2(n_1100),
.B(n_1104),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1035),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_998),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1068),
.B(n_899),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1045),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1035),
.B(n_989),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1092),
.A2(n_990),
.B1(n_819),
.B2(n_920),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1008),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1092),
.A2(n_990),
.B1(n_819),
.B2(n_920),
.Y(n_1275)
);

BUFx4_ASAP7_75t_SL g1276 ( 
.A(n_1008),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_998),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1093),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1092),
.A2(n_1100),
.B1(n_819),
.B2(n_920),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_998),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1207),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1258),
.B1(n_1229),
.B2(n_1136),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1271),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1212),
.A2(n_1216),
.B(n_1220),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1241),
.A2(n_1248),
.B(n_1273),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1271),
.B(n_1166),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1133),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1140),
.Y(n_1289)
);

CKINVDCx11_ASAP7_75t_R g1290 ( 
.A(n_1263),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1157),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1218),
.A2(n_1186),
.B(n_1146),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1145),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1147),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1138),
.A2(n_1258),
.B1(n_1148),
.B2(n_1275),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1153),
.B(n_1151),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1173),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1141),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1267),
.A2(n_1188),
.B1(n_1256),
.B2(n_1279),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1191),
.B(n_1225),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1224),
.B(n_1264),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1144),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1152),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1256),
.A2(n_1279),
.B1(n_1249),
.B2(n_1239),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1185),
.A2(n_1205),
.B(n_1203),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1162),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1249),
.B(n_1176),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1210),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1141),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1165),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1231),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1232),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1180),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1163),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1174),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1141),
.Y(n_1316)
);

INVx8_ASAP7_75t_L g1317 ( 
.A(n_1141),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1219),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1168),
.A2(n_1171),
.B(n_1150),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1134),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1211),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1143),
.A2(n_1252),
.B1(n_1135),
.B2(n_1242),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1213),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1193),
.A2(n_1266),
.B1(n_1177),
.B2(n_1244),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1235),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1238),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1243),
.Y(n_1327)
);

INVx4_ASAP7_75t_SL g1328 ( 
.A(n_1261),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1156),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1154),
.B(n_1226),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1267),
.B(n_1245),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1253),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1228),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1170),
.A2(n_1172),
.B1(n_1265),
.B2(n_1247),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1217),
.B(n_1183),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1163),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1278),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1193),
.A2(n_1169),
.B1(n_1167),
.B2(n_1195),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1269),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1196),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1277),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1163),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1182),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1280),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1214),
.B(n_1222),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_1254),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1137),
.A2(n_1200),
.B(n_1178),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1178),
.B(n_1255),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1233),
.A2(n_1189),
.B1(n_1197),
.B2(n_1201),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1222),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1170),
.B(n_1181),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1276),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1159),
.A2(n_1164),
.B(n_1184),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1192),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1175),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1139),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1246),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1215),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1160),
.B(n_1240),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1222),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1209),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1204),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1175),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1190),
.A2(n_1142),
.B1(n_1240),
.B2(n_1149),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1192),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1187),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1134),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1257),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1142),
.A2(n_1240),
.B1(n_1149),
.B2(n_1160),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1155),
.A2(n_1179),
.B1(n_1227),
.B2(n_1236),
.Y(n_1371)
);

INVx5_ASAP7_75t_L g1372 ( 
.A(n_1261),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1202),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1250),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1270),
.A2(n_1198),
.B(n_1251),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1227),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1199),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1206),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1237),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1237),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1158),
.A2(n_1259),
.B1(n_1272),
.B2(n_1230),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1221),
.A2(n_1208),
.B(n_1234),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1262),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1268),
.B(n_1260),
.Y(n_1384)
);

INVx8_ASAP7_75t_L g1385 ( 
.A(n_1161),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1223),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1139),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1274),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1157),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1207),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1157),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1138),
.A2(n_1092),
.B1(n_1002),
.B2(n_1042),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1138),
.A2(n_1092),
.B1(n_1002),
.B2(n_1042),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1138),
.A2(n_1100),
.B1(n_1279),
.B2(n_1256),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1138),
.A2(n_1092),
.B1(n_1002),
.B2(n_1042),
.Y(n_1395)
);

AO21x1_ASAP7_75t_L g1396 ( 
.A1(n_1138),
.A2(n_1249),
.B(n_1242),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1138),
.B(n_1157),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1153),
.B(n_1151),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1218),
.A2(n_1216),
.B(n_1220),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1321),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1359),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1318),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1362),
.A2(n_1394),
.B(n_1396),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1348),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1359),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1363),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1361),
.B(n_1349),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1354),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1286),
.A2(n_1283),
.B(n_1304),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1363),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1343),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1361),
.B(n_1323),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1313),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1351),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1351),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1285),
.A2(n_1292),
.B(n_1399),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1331),
.B(n_1324),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1305),
.A2(n_1319),
.B(n_1345),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1335),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1345),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1347),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1319),
.A2(n_1305),
.B(n_1350),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1347),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1308),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1372),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1352),
.B(n_1305),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1288),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1390),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1289),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1293),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1294),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1372),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1303),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1352),
.B(n_1282),
.Y(n_1437)
);

AND2x4_ASAP7_75t_SL g1438 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1337),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1322),
.B(n_1296),
.Y(n_1440)
);

OAI321xp33_ASAP7_75t_L g1441 ( 
.A1(n_1295),
.A2(n_1392),
.A3(n_1395),
.B1(n_1393),
.B2(n_1299),
.C(n_1398),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1306),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1310),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1375),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1301),
.B(n_1330),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1397),
.B(n_1311),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1338),
.B(n_1397),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1312),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1325),
.A2(n_1332),
.B(n_1326),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1334),
.A2(n_1302),
.B1(n_1391),
.B2(n_1389),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1327),
.A2(n_1339),
.B(n_1341),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1390),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1344),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1382),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1287),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1291),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1287),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1356),
.B(n_1364),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1377),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1333),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1297),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1329),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1290),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1372),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1298),
.A2(n_1309),
.B(n_1316),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1403),
.B(n_1355),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1403),
.B(n_1355),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1410),
.B(n_1328),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1439),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1400),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1416),
.B(n_1367),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1403),
.B(n_1355),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1456),
.B(n_1373),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1406),
.B(n_1315),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1406),
.B(n_1315),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1400),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1400),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1456),
.B(n_1387),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1439),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1406),
.B(n_1355),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1409),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1461),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1409),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1387),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1437),
.B(n_1336),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1402),
.B(n_1360),
.Y(n_1487)
);

OAI222xp33_ASAP7_75t_L g1488 ( 
.A1(n_1440),
.A2(n_1376),
.B1(n_1309),
.B2(n_1365),
.C1(n_1371),
.C2(n_1370),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1402),
.B(n_1360),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1424),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1404),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1437),
.B(n_1336),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1429),
.B(n_1336),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1314),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1409),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1408),
.B(n_1314),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_SL g1497 ( 
.A(n_1412),
.B(n_1372),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1411),
.A2(n_1384),
.B(n_1381),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1404),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1452),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1429),
.B(n_1314),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1408),
.B(n_1386),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1412),
.A2(n_1372),
.B1(n_1386),
.B2(n_1378),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1429),
.B(n_1342),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1422),
.B(n_1366),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1422),
.B(n_1366),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1440),
.B(n_1316),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1452),
.B(n_1431),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1423),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1431),
.B(n_1284),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1460),
.B(n_1281),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1461),
.Y(n_1512)
);

BUFx4f_ASAP7_75t_SL g1513 ( 
.A(n_1463),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1435),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1485),
.B(n_1460),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1512),
.B(n_1462),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1483),
.B(n_1450),
.C(n_1420),
.D(n_1416),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1494),
.B(n_1462),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1503),
.A2(n_1441),
.B1(n_1420),
.B2(n_1447),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1469),
.A2(n_1413),
.B(n_1447),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1413),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1493),
.B(n_1431),
.Y(n_1522)
);

OAI221xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1487),
.A2(n_1450),
.B1(n_1489),
.B2(n_1502),
.C(n_1475),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1473),
.A2(n_1446),
.B1(n_1458),
.B2(n_1380),
.C(n_1454),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1468),
.B(n_1417),
.Y(n_1525)
);

OAI221xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1487),
.A2(n_1446),
.B1(n_1459),
.B2(n_1441),
.C(n_1426),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1470),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1479),
.B(n_1401),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1459),
.C(n_1427),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1493),
.B(n_1431),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1496),
.A2(n_1425),
.B(n_1427),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1501),
.B(n_1417),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1479),
.B(n_1401),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1407),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1497),
.A2(n_1405),
.B1(n_1454),
.B2(n_1415),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1407),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_L g1537 ( 
.A1(n_1505),
.A2(n_1425),
.B(n_1426),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1497),
.A2(n_1405),
.B1(n_1454),
.B2(n_1415),
.Y(n_1539)
);

NAND4xp25_ASAP7_75t_L g1540 ( 
.A(n_1508),
.B(n_1436),
.C(n_1443),
.D(n_1448),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1501),
.B(n_1417),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1480),
.B(n_1449),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1511),
.B(n_1453),
.C(n_1448),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1480),
.B(n_1449),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1504),
.B(n_1418),
.Y(n_1545)
);

OAI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1505),
.A2(n_1425),
.B(n_1414),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1468),
.B(n_1463),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1504),
.B(n_1449),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1490),
.A2(n_1421),
.B(n_1419),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1486),
.B(n_1418),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_R g1553 ( 
.A(n_1513),
.B(n_1353),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1466),
.B(n_1467),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1468),
.B(n_1463),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1466),
.B(n_1449),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1471),
.B(n_1357),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1472),
.B(n_1489),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1506),
.B(n_1357),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1506),
.A2(n_1438),
.B1(n_1455),
.B2(n_1457),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1488),
.A2(n_1442),
.B1(n_1443),
.B2(n_1453),
.C(n_1430),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1510),
.A2(n_1438),
.B1(n_1484),
.B2(n_1455),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1542),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1527),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1527),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1556),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1532),
.B(n_1486),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1491),
.Y(n_1571)
);

AOI33xp33_ASAP7_75t_L g1572 ( 
.A1(n_1519),
.A2(n_1430),
.A3(n_1432),
.B1(n_1433),
.B2(n_1434),
.B3(n_1436),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1557),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1508),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1548),
.B(n_1484),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1545),
.B(n_1509),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1543),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1525),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1534),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1529),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1525),
.B(n_1514),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1525),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1558),
.B(n_1346),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1521),
.B(n_1514),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1536),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1515),
.B(n_1510),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1518),
.B(n_1470),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1516),
.B(n_1476),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1476),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1529),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1545),
.B(n_1492),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1531),
.B(n_1491),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1522),
.B(n_1509),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1522),
.B(n_1492),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1530),
.B(n_1481),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1530),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1549),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1549),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1477),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1581),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1594),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1573),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1550),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1540),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1583),
.B(n_1531),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1517),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1579),
.A2(n_1563),
.B1(n_1517),
.B2(n_1535),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1567),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1567),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1588),
.B(n_1581),
.Y(n_1618)
);

AOI32xp33_ASAP7_75t_L g1619 ( 
.A1(n_1579),
.A2(n_1546),
.A3(n_1537),
.B1(n_1524),
.B2(n_1539),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1596),
.A2(n_1526),
.B1(n_1523),
.B2(n_1564),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1546),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1573),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1585),
.B(n_1481),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1568),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1578),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1582),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1555),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1585),
.B(n_1481),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1568),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1590),
.A2(n_1405),
.B1(n_1507),
.B2(n_1498),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1594),
.Y(n_1634)
);

NAND2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1584),
.B(n_1585),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1603),
.A2(n_1482),
.B1(n_1562),
.B2(n_1495),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1594),
.B(n_1435),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1592),
.Y(n_1638)
);

NAND2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1589),
.B(n_1435),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1573),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1482),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1603),
.B(n_1577),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1599),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1577),
.B(n_1482),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1578),
.B(n_1499),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1614),
.A2(n_1571),
.B(n_1604),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1590),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1616),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1616),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1609),
.B(n_1580),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1634),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1617),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1634),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1613),
.A2(n_1604),
.B(n_1537),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1571),
.Y(n_1657)
);

AOI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1612),
.A2(n_1566),
.B(n_1565),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1629),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.B(n_1597),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1607),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1607),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1627),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1611),
.B(n_1597),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1623),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1610),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1618),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1674)
);

OAI211xp5_ASAP7_75t_L g1675 ( 
.A1(n_1608),
.A2(n_1290),
.B(n_1553),
.C(n_1576),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1610),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1632),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1646),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1638),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1620),
.A2(n_1577),
.B1(n_1600),
.B2(n_1591),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1591),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1618),
.A2(n_1576),
.B(n_1575),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1633),
.A2(n_1605),
.B(n_1598),
.C(n_1575),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1607),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1644),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1595),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1650),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1655),
.Y(n_1692)
);

AND3x1_ASAP7_75t_L g1693 ( 
.A(n_1663),
.B(n_1631),
.C(n_1626),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1642),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1353),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1659),
.A2(n_1405),
.B1(n_1630),
.B2(n_1636),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1650),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1660),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1660),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1671),
.B(n_1670),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1676),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1655),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1662),
.B(n_1630),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1662),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1661),
.B(n_1642),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1665),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1653),
.B(n_1374),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1676),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1651),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1674),
.A2(n_1630),
.B1(n_1635),
.B2(n_1642),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1668),
.B(n_1608),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1374),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1654),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1648),
.A2(n_1635),
.B(n_1637),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1656),
.A2(n_1405),
.B1(n_1454),
.B2(n_1624),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1687),
.A2(n_1647),
.B1(n_1658),
.B2(n_1657),
.C(n_1682),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1649),
.B(n_1625),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

CKINVDCx16_ASAP7_75t_R g1719 ( 
.A(n_1688),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1647),
.A2(n_1688),
.B1(n_1684),
.B2(n_1652),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1664),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1673),
.B(n_1625),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1672),
.A2(n_1624),
.B1(n_1640),
.B2(n_1566),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1666),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1667),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1715),
.A2(n_1685),
.B1(n_1689),
.B2(n_1686),
.C(n_1683),
.Y(n_1726)
);

NOR2xp67_ASAP7_75t_SL g1727 ( 
.A(n_1719),
.B(n_1369),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1669),
.B(n_1689),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1702),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1700),
.A2(n_1605),
.B1(n_1598),
.B2(n_1681),
.C(n_1679),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1693),
.A2(n_1676),
.B(n_1678),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1691),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1706),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1694),
.B(n_1680),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1711),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1690),
.B(n_1595),
.Y(n_1738)
);

OAI32xp33_ASAP7_75t_L g1739 ( 
.A1(n_1710),
.A2(n_1635),
.A3(n_1637),
.B1(n_1598),
.B2(n_1605),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1714),
.A2(n_1631),
.B(n_1626),
.C(n_1385),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1695),
.B(n_1707),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1720),
.B(n_1569),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1718),
.B(n_1569),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1711),
.B(n_1574),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1690),
.B(n_1574),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1565),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1701),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1696),
.A2(n_1637),
.B(n_1639),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1727),
.B(n_1717),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1737),
.B(n_1724),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1722),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1734),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1743),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1735),
.B(n_1694),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1737),
.B(n_1708),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1751),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1735),
.B(n_1705),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1736),
.B(n_1705),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1708),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1741),
.B(n_1340),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1731),
.B(n_1713),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1741),
.B(n_1340),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1730),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1749),
.B(n_1713),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1748),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1721),
.Y(n_1771)
);

AOI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1726),
.B1(n_1732),
.B2(n_1750),
.C(n_1742),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1764),
.A2(n_1369),
.B(n_1733),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1755),
.A2(n_1740),
.B1(n_1746),
.B2(n_1744),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1767),
.A2(n_1739),
.B1(n_1747),
.B2(n_1697),
.C(n_1699),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1766),
.A2(n_1745),
.B(n_1699),
.Y(n_1776)
);

O2A1O1Ixp33_ASAP7_75t_SL g1777 ( 
.A1(n_1768),
.A2(n_1358),
.B(n_1725),
.C(n_1721),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1758),
.B(n_1738),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1760),
.A2(n_1698),
.B(n_1723),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1760),
.B(n_1725),
.C(n_1698),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_SL g1781 ( 
.A(n_1759),
.B(n_1388),
.C(n_1358),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1753),
.B(n_1738),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1758),
.A2(n_1385),
.B(n_1672),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1778),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1772),
.A2(n_1761),
.B1(n_1762),
.B2(n_1763),
.Y(n_1785)
);

NOR2xp67_ASAP7_75t_L g1786 ( 
.A(n_1782),
.B(n_1761),
.Y(n_1786)
);

AND4x1_ASAP7_75t_L g1787 ( 
.A(n_1781),
.B(n_1762),
.C(n_1770),
.D(n_1763),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1780),
.B(n_1756),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1779),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1775),
.B(n_1765),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1776),
.Y(n_1792)
);

OAI211xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1774),
.A2(n_1757),
.B(n_1754),
.C(n_1752),
.Y(n_1793)
);

NOR4xp25_ASAP7_75t_SL g1794 ( 
.A(n_1777),
.B(n_1770),
.C(n_1757),
.D(n_1769),
.Y(n_1794)
);

AND5x1_ASAP7_75t_L g1795 ( 
.A(n_1787),
.B(n_1783),
.C(n_1773),
.D(n_1769),
.E(n_1385),
.Y(n_1795)
);

AOI21xp33_ASAP7_75t_L g1796 ( 
.A1(n_1789),
.A2(n_1677),
.B(n_1385),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1786),
.B(n_1677),
.Y(n_1797)
);

NAND4xp75_ASAP7_75t_L g1798 ( 
.A(n_1791),
.B(n_1641),
.C(n_1645),
.D(n_1640),
.Y(n_1798)
);

NOR4xp25_ASAP7_75t_L g1799 ( 
.A(n_1793),
.B(n_1641),
.C(n_1645),
.D(n_1606),
.Y(n_1799)
);

NOR3xp33_ASAP7_75t_L g1800 ( 
.A(n_1790),
.B(n_1792),
.C(n_1785),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1788),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1784),
.A2(n_1794),
.B1(n_1639),
.B2(n_1606),
.C(n_1432),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1800),
.A2(n_1639),
.B1(n_1498),
.B2(n_1451),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1799),
.B(n_1570),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1801),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1798),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1797),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1802),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1796),
.B(n_1570),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1806),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1805),
.Y(n_1811)
);

NAND4xp75_ASAP7_75t_L g1812 ( 
.A(n_1808),
.B(n_1795),
.C(n_1602),
.D(n_1464),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1433),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1804),
.B(n_1601),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1811),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1810),
.B(n_1813),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1812),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1815),
.A2(n_1810),
.B1(n_1809),
.B2(n_1814),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1818),
.B(n_1816),
.C(n_1817),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1803),
.B1(n_1601),
.B2(n_1597),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1819),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1821),
.A2(n_1451),
.B1(n_1368),
.B2(n_1379),
.Y(n_1822)
);

XNOR2xp5_ASAP7_75t_L g1823 ( 
.A(n_1820),
.B(n_1281),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1823),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1822),
.A2(n_1317),
.B(n_1428),
.Y(n_1825)
);

OR2x6_ASAP7_75t_L g1826 ( 
.A(n_1824),
.B(n_1320),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1825),
.B1(n_1383),
.B2(n_1320),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1368),
.B1(n_1379),
.B2(n_1383),
.C(n_1442),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1465),
.B(n_1514),
.C(n_1444),
.Y(n_1829)
);


endmodule