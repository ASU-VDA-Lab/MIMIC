module fake_jpeg_1751_n_99 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_38),
.C(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_33),
.B1(n_29),
.B2(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_47),
.B1(n_42),
.B2(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_49),
.B1(n_28),
.B2(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_56),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_26),
.B(n_20),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_72),
.B(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_18),
.B1(n_17),
.B2(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_83),
.C(n_85),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_1),
.C(n_4),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_4),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.C(n_86),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_6),
.C(n_7),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_80),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_82),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_6),
.C(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_8),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_8),
.B(n_9),
.Y(n_99)
);


endmodule