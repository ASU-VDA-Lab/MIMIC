module fake_jpeg_11352_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_88),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_63),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_66),
.Y(n_180)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_68),
.B(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_77),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_1),
.CON(n_85),
.SN(n_85)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_47),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_15),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_10),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_65),
.Y(n_127)
);

CKINVDCx9p33_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_35),
.B(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_95),
.B(n_102),
.Y(n_185)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_35),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_110),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_101),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_107),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_39),
.B(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_111),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_27),
.B(n_9),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_30),
.A2(n_1),
.B(n_3),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_47),
.B(n_24),
.C(n_49),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_3),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_56),
.B1(n_37),
.B2(n_55),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_122),
.A2(n_125),
.B1(n_134),
.B2(n_138),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_124),
.A2(n_179),
.A3(n_129),
.B1(n_145),
.B2(n_162),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_30),
.B1(n_37),
.B2(n_55),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_51),
.B1(n_46),
.B2(n_33),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_172),
.C(n_161),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_28),
.B1(n_53),
.B2(n_38),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_173),
.B1(n_175),
.B2(n_178),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_40),
.B(n_38),
.C(n_20),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_132),
.A2(n_140),
.B(n_128),
.C(n_134),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_33),
.B1(n_53),
.B2(n_28),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_136),
.B(n_167),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_28),
.B1(n_53),
.B2(n_40),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_33),
.B1(n_45),
.B2(n_43),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_140),
.A2(n_155),
.B1(n_162),
.B2(n_169),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_45),
.B1(n_43),
.B2(n_27),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_47),
.B1(n_49),
.B2(n_24),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_194),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_67),
.B(n_4),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_47),
.B1(n_49),
.B2(n_7),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_170),
.B(n_139),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_78),
.B(n_6),
.C(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_69),
.A2(n_8),
.B1(n_9),
.B2(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_87),
.A2(n_113),
.B1(n_106),
.B2(n_104),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_74),
.A2(n_8),
.B1(n_85),
.B2(n_115),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_176),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_92),
.A2(n_8),
.B1(n_96),
.B2(n_72),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_75),
.A2(n_80),
.B1(n_114),
.B2(n_99),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_185),
.B(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_105),
.A2(n_64),
.B1(n_117),
.B2(n_79),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_176),
.B1(n_146),
.B2(n_137),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_64),
.B(n_117),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_88),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_202),
.B(n_209),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_204),
.B(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_124),
.A2(n_172),
.B1(n_150),
.B2(n_132),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVx5_ASAP7_75t_SL g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_216),
.Y(n_276)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_210),
.A2(n_214),
.B1(n_254),
.B2(n_259),
.Y(n_275)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_131),
.Y(n_211)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_146),
.A2(n_184),
.B1(n_168),
.B2(n_177),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_138),
.A2(n_198),
.B1(n_186),
.B2(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_147),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_151),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_247),
.C(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

OR2x4_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_148),
.B(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_223),
.B(n_229),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_184),
.A2(n_168),
.B1(n_177),
.B2(n_180),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_240),
.Y(n_287)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_153),
.B(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_171),
.B(n_144),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_144),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_231),
.B(n_234),
.Y(n_309)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_121),
.Y(n_234)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_121),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_122),
.B1(n_159),
.B2(n_195),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_237),
.A2(n_245),
.B1(n_206),
.B2(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_159),
.B(n_123),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_239),
.B(n_241),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_123),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_149),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_248),
.Y(n_288)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_252),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_186),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_152),
.A2(n_187),
.B1(n_189),
.B2(n_181),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_253),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_152),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_255),
.Y(n_292)
);

INVx4_ASAP7_75t_SL g251 ( 
.A(n_157),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_189),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_157),
.C(n_197),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_197),
.A2(n_130),
.B1(n_178),
.B2(n_124),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_185),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_264),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_150),
.B(n_139),
.CI(n_170),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_243),
.C(n_203),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_130),
.A2(n_93),
.B1(n_89),
.B2(n_84),
.Y(n_259)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_129),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_262),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_150),
.B(n_194),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_176),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_263),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_132),
.B(n_185),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_205),
.A2(n_254),
.B1(n_264),
.B2(n_256),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_279),
.B(n_295),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_199),
.A2(n_204),
.B1(n_249),
.B2(n_238),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_203),
.B1(n_199),
.B2(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_285),
.A2(n_294),
.B1(n_261),
.B2(n_251),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_200),
.B(n_228),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_291),
.B(n_307),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_247),
.B1(n_203),
.B2(n_252),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_216),
.B(n_226),
.Y(n_295)
);

FAx1_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_282),
.CI(n_271),
.CON(n_343),
.SN(n_343)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_257),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_210),
.A2(n_201),
.B1(n_232),
.B2(n_244),
.Y(n_299)
);

INVx11_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_225),
.B(n_217),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_217),
.B(n_230),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_208),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_316),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_265),
.A2(n_227),
.B1(n_219),
.B2(n_246),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_317),
.B1(n_320),
.B2(n_335),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_287),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_265),
.A2(n_219),
.B1(n_245),
.B2(n_220),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_215),
.B1(n_218),
.B2(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_276),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_273),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_273),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_329),
.Y(n_368)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_236),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_331),
.B(n_341),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_255),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_272),
.A2(n_297),
.B(n_271),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_343),
.B(n_307),
.Y(n_379)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_280),
.B(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_280),
.B(n_291),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_310),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_272),
.A2(n_284),
.B1(n_296),
.B2(n_290),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_284),
.B1(n_286),
.B2(n_293),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_348),
.B(n_278),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_341),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_353),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_369),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_362),
.B1(n_364),
.B2(n_335),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_283),
.C(n_279),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_266),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_361),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_306),
.C(n_281),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_318),
.A2(n_275),
.B1(n_289),
.B2(n_286),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_303),
.B1(n_289),
.B2(n_275),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_303),
.C(n_299),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_370),
.B(n_376),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_375),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_374),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_322),
.B(n_278),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_342),
.B(n_343),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_400),
.B(n_379),
.Y(n_416)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_325),
.B1(n_327),
.B2(n_318),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_391),
.B1(n_361),
.B2(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_316),
.Y(n_385)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_348),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_389),
.Y(n_405)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_342),
.B1(n_332),
.B2(n_343),
.Y(n_391)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_392),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_398),
.Y(n_409)
);

BUFx12_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_396),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_331),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_401),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_320),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_399),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_370),
.B(n_343),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_368),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_317),
.B1(n_314),
.B2(n_330),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_363),
.B1(n_330),
.B2(n_366),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_345),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_403),
.B(n_315),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_353),
.C(n_349),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_415),
.C(n_420),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_419),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_404),
.C(n_387),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_393),
.C(n_383),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_354),
.C(n_326),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_398),
.A2(n_330),
.B1(n_363),
.B2(n_350),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_426),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_400),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_372),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_424),
.B(n_425),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_350),
.B1(n_367),
.B2(n_366),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_391),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_428),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_393),
.B(n_401),
.C(n_383),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_435),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_382),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_433),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_416),
.A2(n_392),
.B(n_384),
.Y(n_433)
);

AOI221xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_315),
.B1(n_337),
.B2(n_395),
.C(n_357),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_434),
.B(n_390),
.Y(n_456)
);

AO221x1_ASAP7_75t_L g435 ( 
.A1(n_411),
.A2(n_357),
.B1(n_372),
.B2(n_367),
.C(n_365),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_402),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_418),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_438),
.B(n_439),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_423),
.C(n_413),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_424),
.C(n_409),
.Y(n_444)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_442),
.Y(n_452)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_399),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_407),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_444),
.B(n_446),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_430),
.A2(n_408),
.B1(n_421),
.B2(n_426),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_409),
.B1(n_418),
.B2(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_417),
.C(n_419),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_453),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_437),
.Y(n_463)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_433),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_456),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_436),
.C(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_461),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_452),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_428),
.B(n_429),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_462),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_427),
.C(n_439),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_451),
.A2(n_431),
.B(n_430),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_453),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_465),
.A2(n_445),
.B1(n_432),
.B2(n_455),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_462),
.C(n_466),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_458),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_471),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_448),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_467),
.B1(n_469),
.B2(n_464),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_460),
.B(n_443),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_474),
.B(n_463),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_472),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_478),
.A2(n_480),
.B1(n_414),
.B2(n_419),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g479 ( 
.A1(n_467),
.A2(n_455),
.B(n_381),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_479),
.A2(n_419),
.B1(n_414),
.B2(n_365),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_473),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_477),
.C(n_476),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_482),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g487 ( 
.A1(n_483),
.A2(n_389),
.A3(n_396),
.B1(n_359),
.B2(n_484),
.C1(n_300),
.C2(n_274),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_486),
.B(n_487),
.Y(n_488)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_484),
.C(n_359),
.Y(n_489)
);

AOI322xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_274),
.A3(n_396),
.B1(n_300),
.B2(n_333),
.C1(n_328),
.C2(n_323),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_488),
.Y(n_491)
);


endmodule