module fake_jpeg_1136_n_123 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_31),
.B(n_18),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_22),
.B1(n_16),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_36)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_3),
.Y(n_37)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_7),
.B1(n_27),
.B2(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_15),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_57),
.B1(n_52),
.B2(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_13),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_18),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_43),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_64),
.B(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_32),
.B(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_18),
.B1(n_43),
.B2(n_67),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_51),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_55),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_81),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_72),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_71),
.B1(n_83),
.B2(n_78),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_74),
.C(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.C(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_89),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_93),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_103),
.B(n_92),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_100),
.Y(n_113)
);

AO221x1_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_106),
.B1(n_102),
.B2(n_97),
.C(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_105),
.B(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_115),
.B1(n_114),
.B2(n_116),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);


endmodule