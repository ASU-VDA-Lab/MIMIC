module real_jpeg_24849_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_21),
.B1(n_25),
.B2(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_21),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_9),
.B1(n_53),
.B2(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_25),
.B(n_43),
.C(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_24),
.B(n_77),
.C(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_36),
.B1(n_79),
.B2(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_31),
.C(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_7),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_7),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_7),
.B(n_63),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_110),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_72),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_16),
.B(n_72),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_54),
.C(n_58),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_17),
.B(n_178),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_75),
.Y(n_74)
);

FAx1_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.CI(n_39),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_20),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_21),
.A2(n_25),
.B1(n_43),
.B2(n_47),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_23),
.A2(n_25),
.B(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_23),
.A2(n_24),
.B1(n_79),
.B2(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_27),
.B(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_28),
.A2(n_35),
.B(n_37),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_37),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_30),
.A2(n_31),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_31),
.B(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_34),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_44),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_37),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_48),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_41),
.B(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_45),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_45),
.B(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_49),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_54),
.B(n_58),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_55),
.A2(n_57),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_55),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_57),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_62),
.B(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_61),
.B(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_63),
.B(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_63),
.B(n_127),
.Y(n_126)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_68),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_70),
.B(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_86),
.B2(n_87),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B1(n_98),
.B2(n_108),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_105),
.B2(n_106),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_175),
.B(n_179),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_161),
.B(n_174),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_140),
.B(n_160),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_130),
.B2(n_139),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_129),
.C(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_148),
.B(n_159),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_155),
.B(n_158),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_163),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_169),
.C(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_177),
.Y(n_179)
);


endmodule