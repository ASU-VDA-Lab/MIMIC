module fake_jpeg_28966_n_360 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_14),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_15),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_21),
.B(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_55),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_28),
.B1(n_29),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_72),
.B1(n_49),
.B2(n_32),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_34),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_60),
.B(n_62),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_29),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_31),
.B(n_26),
.C(n_25),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_84),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_21),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_28),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_18),
.C(n_22),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_SL g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_17),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_17),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_40),
.B1(n_46),
.B2(n_36),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_94),
.A2(n_99),
.B1(n_116),
.B2(n_121),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_28),
.B1(n_54),
.B2(n_17),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_59),
.A2(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_105),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_126),
.B(n_22),
.Y(n_160)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_78),
.Y(n_143)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_120),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_39),
.B1(n_44),
.B2(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_122),
.B1(n_55),
.B2(n_65),
.Y(n_138)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_44),
.B1(n_42),
.B2(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_125),
.Y(n_131)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_42),
.B1(n_44),
.B2(n_34),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_18),
.A3(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_127),
.Y(n_139)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_20),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_91),
.B1(n_61),
.B2(n_63),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_138),
.B1(n_147),
.B2(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_78),
.C(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_15),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_153),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_92),
.A2(n_77),
.B1(n_67),
.B2(n_73),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_85),
.CON(n_148),
.SN(n_148)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_58),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_92),
.A2(n_67),
.B1(n_58),
.B2(n_57),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_112),
.B(n_68),
.C(n_87),
.Y(n_153)
);

AND2x4_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_77),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_160),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_57),
.C(n_73),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_35),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_77),
.A3(n_81),
.B1(n_90),
.B2(n_63),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_22),
.Y(n_184)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_116),
.B1(n_126),
.B2(n_99),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_174),
.B1(n_176),
.B2(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_128),
.B1(n_102),
.B2(n_118),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_180),
.B1(n_186),
.B2(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_118),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_102),
.B1(n_129),
.B2(n_106),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_113),
.B(n_111),
.C(n_120),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_115),
.B1(n_107),
.B2(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_181),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_98),
.B1(n_97),
.B2(n_93),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_81),
.B1(n_93),
.B2(n_104),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_187),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_160),
.B(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_189),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_131),
.B(n_13),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_196),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_138),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_141),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_35),
.B1(n_16),
.B2(n_11),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_11),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_173),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_137),
.B(n_143),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_211),
.B(n_170),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_186),
.B1(n_172),
.B2(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_221),
.B1(n_225),
.B2(n_182),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_133),
.C(n_131),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_210),
.C(n_213),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_133),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_230),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_132),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_153),
.B(n_144),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_153),
.A3(n_132),
.B1(n_154),
.B2(n_147),
.C1(n_142),
.C2(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_154),
.C(n_141),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_193),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_188),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_154),
.C(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_154),
.B1(n_155),
.B2(n_130),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_176),
.A2(n_155),
.B1(n_130),
.B2(n_35),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_170),
.A2(n_130),
.B(n_35),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_227),
.B(n_211),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_172),
.B(n_0),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_233),
.A2(n_5),
.B(n_6),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_167),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_242),
.B(n_247),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_224),
.B1(n_205),
.B2(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_180),
.B1(n_194),
.B2(n_177),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_258),
.B1(n_223),
.B2(n_230),
.Y(n_275)
);

XNOR2x2_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_169),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_206),
.B(n_187),
.Y(n_245)
);

NOR4xp25_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_2),
.C(n_4),
.D(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_165),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_197),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_208),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_196),
.C(n_181),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_220),
.C(n_203),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_214),
.B1(n_210),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_213),
.B1(n_209),
.B2(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_190),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_185),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_202),
.B(n_178),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_259),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_175),
.B1(n_195),
.B2(n_164),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_175),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_164),
.B(n_16),
.C(n_3),
.D(n_4),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_274),
.C(n_240),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_263),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_266),
.B1(n_277),
.B2(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_205),
.B(n_224),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_233),
.B(n_270),
.Y(n_286)
);

XOR2x1_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_231),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_238),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_231),
.C(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_279),
.B1(n_249),
.B2(n_253),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_244),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_247),
.A3(n_255),
.B1(n_257),
.B2(n_254),
.C1(n_259),
.C2(n_237),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_296),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_289),
.B(n_299),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_294),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_243),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_300),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_265),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_302),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_267),
.B1(n_272),
.B2(n_278),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_251),
.C(n_256),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_235),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_278),
.B(n_245),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g304 ( 
.A(n_265),
.B(n_263),
.C(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_306),
.A2(n_312),
.B1(n_320),
.B2(n_275),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_271),
.B1(n_276),
.B2(n_250),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_318),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_304),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_269),
.B1(n_277),
.B2(n_268),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_286),
.B(n_292),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_297),
.C(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_328),
.Y(n_334)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_293),
.B(n_288),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_323),
.A2(n_326),
.B1(n_319),
.B2(n_239),
.Y(n_341)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_291),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_327),
.A2(n_256),
.B1(n_7),
.B2(n_16),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_273),
.Y(n_328)
);

NAND4xp25_ASAP7_75t_SL g329 ( 
.A(n_310),
.B(n_289),
.C(n_279),
.D(n_239),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_282),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_320),
.A2(n_280),
.B(n_273),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_319),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_317),
.A2(n_299),
.B(n_246),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_307),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_316),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_337),
.Y(n_351)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_341),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_322),
.B(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_325),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_348),
.Y(n_353)
);

OAI211xp5_ASAP7_75t_L g348 ( 
.A1(n_342),
.A2(n_321),
.B(n_333),
.C(n_329),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_339),
.B(n_323),
.CI(n_330),
.CON(n_349),
.SN(n_349)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_344),
.C(n_351),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_334),
.A2(n_7),
.B(n_16),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_350),
.A2(n_342),
.B(n_338),
.C(n_341),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_352),
.Y(n_357)
);

NAND4xp25_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_355),
.C(n_356),
.D(n_349),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_16),
.C(n_346),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_353),
.B(n_356),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_357),
.Y(n_360)
);


endmodule