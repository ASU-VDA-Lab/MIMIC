module fake_jpeg_26416_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_50),
.Y(n_87)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_55),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_52),
.C(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_52),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_53),
.B1(n_58),
.B2(n_57),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_103),
.B1(n_106),
.B2(n_67),
.Y(n_117)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_104),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_102),
.B1(n_61),
.B2(n_50),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_53),
.B1(n_58),
.B2(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_49),
.B1(n_62),
.B2(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_0),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_84),
.B(n_89),
.C(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_61),
.B1(n_89),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_114),
.B1(n_116),
.B2(n_92),
.Y(n_120)
);

OAI22x1_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_61),
.B1(n_79),
.B2(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_121),
.B1(n_110),
.B2(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_99),
.B1(n_101),
.B2(n_92),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_118),
.B1(n_124),
.B2(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_65),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_97),
.C(n_60),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_79),
.C(n_96),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_68),
.B(n_63),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_54),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_66),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_17),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_138),
.B(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_132),
.B1(n_139),
.B2(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_3),
.C(n_4),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_15),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_19),
.C(n_43),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_16),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_3),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_1),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_149),
.C(n_150),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_21),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_45),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_145),
.B1(n_148),
.B2(n_137),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_143),
.CI(n_128),
.CON(n_155),
.SN(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_153),
.B1(n_152),
.B2(n_149),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_155),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_147),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_36),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_31),
.B(n_30),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_34),
.B(n_29),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_26),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_25),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_4),
.Y(n_164)
);


endmodule