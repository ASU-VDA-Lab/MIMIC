module fake_jpeg_27635_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_45),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_18),
.B(n_17),
.C(n_30),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_44),
.B(n_16),
.C(n_34),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_58),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_41),
.B1(n_42),
.B2(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_36),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_65),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_95),
.B1(n_97),
.B2(n_103),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_39),
.B1(n_24),
.B2(n_20),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_76),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_22),
.B1(n_16),
.B2(n_34),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_21),
.B(n_29),
.C(n_10),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_36),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_90),
.C(n_35),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_37),
.B(n_45),
.C(n_36),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_99),
.B1(n_39),
.B2(n_35),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_22),
.B1(n_40),
.B2(n_41),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_80),
.B1(n_88),
.B2(n_91),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_79),
.Y(n_129)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_92),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_58),
.B(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_23),
.B1(n_42),
.B2(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_53),
.B(n_49),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_51),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_116),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_42),
.A3(n_36),
.B1(n_21),
.B2(n_37),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_63),
.B1(n_26),
.B2(n_35),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_134),
.B1(n_98),
.B2(n_96),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_72),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_21),
.C(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_29),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_66),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_128),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_24),
.C(n_20),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_81),
.B1(n_83),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_24),
.B1(n_20),
.B2(n_39),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_137),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_139),
.A2(n_102),
.B1(n_80),
.B2(n_91),
.Y(n_195)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_64),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_81),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_142),
.B(n_148),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_145),
.B1(n_113),
.B2(n_122),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_73),
.B1(n_104),
.B2(n_74),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_151),
.B(n_163),
.Y(n_194)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_162),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_73),
.B1(n_74),
.B2(n_68),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_125),
.B1(n_107),
.B2(n_119),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_68),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_68),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_165),
.B(n_136),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_108),
.C(n_116),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_187),
.C(n_136),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_110),
.B1(n_106),
.B2(n_115),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_157),
.A2(n_106),
.B1(n_111),
.B2(n_110),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_185),
.B1(n_195),
.B2(n_197),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_120),
.B(n_124),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_182),
.B(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_179),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_120),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_177),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_124),
.A3(n_112),
.B1(n_128),
.B2(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_151),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_159),
.B1(n_154),
.B2(n_162),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_122),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_163),
.C(n_153),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_152),
.B1(n_163),
.B2(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_191),
.B1(n_187),
.B2(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_71),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_118),
.B1(n_117),
.B2(n_132),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_132),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_85),
.B1(n_75),
.B2(n_99),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_219),
.B1(n_226),
.B2(n_172),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_146),
.B(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_202),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_189),
.B(n_191),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_165),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_204),
.B(n_214),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_212),
.Y(n_233)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_222),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_179),
.A2(n_148),
.B1(n_136),
.B2(n_88),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_84),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_87),
.C(n_78),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_227),
.C(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_39),
.C(n_14),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_200),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_192),
.B1(n_183),
.B2(n_190),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_236),
.B1(n_251),
.B2(n_210),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_186),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_182),
.B1(n_181),
.B2(n_172),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_173),
.C(n_178),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_249),
.C(n_250),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_170),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_14),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_11),
.C(n_10),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_10),
.C(n_9),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_242),
.C(n_228),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_229),
.B(n_234),
.Y(n_255)
);

OAI322xp33_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_270),
.A3(n_245),
.B1(n_250),
.B2(n_249),
.C1(n_239),
.C2(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_210),
.B(n_211),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_198),
.B1(n_225),
.B2(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_227),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_220),
.B(n_202),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_230),
.B(n_203),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_201),
.B(n_224),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_219),
.B(n_223),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_206),
.B1(n_208),
.B2(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_206),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_9),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_278),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_233),
.B(n_232),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_266),
.B(n_261),
.Y(n_289)
);

OAI322xp33_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_240),
.A3(n_251),
.B1(n_9),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_0),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_0),
.C(n_1),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_271),
.C(n_268),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_281),
.B(n_288),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_299),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_253),
.B1(n_258),
.B2(n_252),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_295),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_285),
.B1(n_275),
.B2(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_284),
.B1(n_285),
.B2(n_282),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_255),
.B1(n_262),
.B2(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_3),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.C(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_8),
.C(n_5),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_305),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_273),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_309),
.C(n_292),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_273),
.B(n_276),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_275),
.B(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_312),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_301),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_288),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_291),
.B1(n_304),
.B2(n_303),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_301),
.C(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_304),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_314),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_323),
.B1(n_322),
.B2(n_318),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_318),
.A3(n_290),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_329)
);

OAI311xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.C1(n_8),
.Y(n_330)
);


endmodule