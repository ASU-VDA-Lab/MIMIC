module fake_jpeg_25423_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_31),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_21),
.B(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_26),
.C(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_31),
.C(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_22),
.B1(n_42),
.B2(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_71),
.B1(n_74),
.B2(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_69),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_42),
.B1(n_36),
.B2(n_34),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_42),
.B1(n_30),
.B2(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_32),
.B1(n_33),
.B2(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_21),
.B1(n_17),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_77),
.B1(n_33),
.B2(n_17),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_18),
.B1(n_23),
.B2(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_39),
.B1(n_40),
.B2(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_20),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_21),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_40),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_99),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_58),
.B1(n_55),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_66),
.B1(n_61),
.B2(n_64),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_80),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_84),
.Y(n_104)
);

FAx1_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_106),
.CI(n_80),
.CON(n_129),
.SN(n_129)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_79),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_27),
.B1(n_19),
.B2(n_69),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_62),
.C(n_65),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_133),
.Y(n_182)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_108),
.B(n_100),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_136),
.B1(n_115),
.B2(n_118),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_83),
.C(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_61),
.B1(n_73),
.B2(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_93),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_110),
.B1(n_119),
.B2(n_102),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_142),
.B1(n_143),
.B2(n_148),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_89),
.B1(n_66),
.B2(n_88),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_109),
.B1(n_94),
.B2(n_116),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_119),
.B1(n_103),
.B2(n_99),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_90),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_60),
.C(n_29),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_115),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_64),
.B1(n_29),
.B2(n_23),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_158),
.B1(n_160),
.B2(n_143),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_152),
.A2(n_172),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_161),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_106),
.CI(n_96),
.CON(n_157),
.SN(n_157)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_18),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_93),
.B1(n_117),
.B2(n_100),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_165),
.B(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_116),
.B1(n_117),
.B2(n_115),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_112),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_122),
.B1(n_148),
.B2(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_150),
.B1(n_162),
.B2(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_108),
.B(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_101),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_171),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_24),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_11),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_24),
.B(n_1),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_9),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_180),
.B1(n_176),
.B2(n_174),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_24),
.B(n_1),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_121),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_181),
.A2(n_3),
.B(n_4),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_195),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_122),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_202),
.B(n_207),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_120),
.C(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_190),
.C(n_194),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_189),
.B1(n_205),
.B2(n_160),
.Y(n_224)
);

AOI22x1_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_126),
.B1(n_138),
.B2(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_199),
.B1(n_166),
.B2(n_183),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_124),
.B1(n_134),
.B2(n_29),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_149),
.C(n_23),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_209),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_23),
.B1(n_18),
.B2(n_8),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_181),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_8),
.B(n_15),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_150),
.A2(n_18),
.B1(n_1),
.B2(n_3),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_0),
.B(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_152),
.A2(n_4),
.B(n_5),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_169),
.C(n_163),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_216),
.C(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_164),
.C(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_157),
.B1(n_158),
.B2(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_199),
.B1(n_209),
.B2(n_192),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_157),
.C(n_156),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_180),
.B1(n_177),
.B2(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_174),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_4),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_207),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_200),
.C(n_185),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_9),
.C(n_14),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_185),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_247),
.B1(n_217),
.B2(n_213),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_201),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_240),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_226),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_191),
.B1(n_210),
.B2(n_205),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_208),
.B(n_207),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_233),
.B1(n_211),
.B2(n_184),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_251),
.B1(n_222),
.B2(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_214),
.C(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_253),
.B(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_220),
.C(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_265),
.C(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_262),
.B1(n_246),
.B2(n_235),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_232),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_263),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_223),
.B1(n_221),
.B2(n_211),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_233),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_13),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_8),
.C(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_271),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_235),
.B(n_248),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_272),
.B(n_279),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_247),
.B1(n_252),
.B2(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.C(n_280),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_265),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_277),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_13),
.C(n_15),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_255),
.B(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_288),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_256),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_13),
.B(n_15),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_R g290 ( 
.A(n_280),
.B(n_7),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_269),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_276),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_6),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_5),
.C(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_287),
.C(n_282),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_300),
.B(n_291),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_303),
.B(n_300),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_301),
.C(n_296),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_292),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_297),
.B(n_7),
.Y(n_309)
);


endmodule