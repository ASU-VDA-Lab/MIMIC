module fake_netlist_6_59_n_2084 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2084);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2084;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_153),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_52),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_70),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_4),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_64),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_112),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_41),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_114),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_171),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_30),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_16),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_21),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_170),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_158),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_99),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_88),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_34),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_77),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_204),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_79),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_118),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_55),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_7),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_135),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_102),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_115),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_75),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_189),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_85),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_205),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_66),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_91),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_78),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_199),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_188),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_134),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_164),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_68),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_156),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_86),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_84),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_0),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_174),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_163),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_106),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_178),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_132),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_201),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_53),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_62),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_172),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_28),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_206),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_33),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_187),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_33),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_125),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_175),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_29),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_35),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_61),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_90),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_121),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_81),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_179),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_35),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_51),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_60),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_122),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_147),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_137),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_9),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_26),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_34),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_23),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_11),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_40),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_109),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_57),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_180),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_74),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_82),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_72),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_29),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_13),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_131),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_14),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_6),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_87),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_200),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_8),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_93),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_126),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_49),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_133),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_161),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_119),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_44),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_177),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_64),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_32),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_113),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_6),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_185),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_136),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_50),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_14),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_39),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_148),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_25),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_58),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_63),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_23),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_32),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_38),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_142),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_111),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_101),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_53),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_169),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_49),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_94),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_48),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_155),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_139),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_76),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_69),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_61),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_15),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_65),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_117),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_19),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_60),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_110),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_2),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_203),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_37),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_37),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_166),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_13),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_63),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_128),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_182),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_59),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_22),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_173),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_80),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_143),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_123),
.Y(n_406)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_57),
.Y(n_407)
);

INVx4_ASAP7_75t_R g408 ( 
.A(n_89),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_27),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_48),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_50),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_55),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_18),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_145),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_233),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_222),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_282),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_231),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_208),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_216),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_1),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_293),
.B(n_73),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_285),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_287),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_244),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_320),
.B(n_2),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_292),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_286),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_321),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_347),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_249),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_249),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_299),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_262),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_262),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_317),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_391),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_317),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_303),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_309),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_404),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_311),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_248),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_252),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_254),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_333),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_216),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_295),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_241),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_333),
.B(n_3),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_255),
.B(n_83),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_217),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_313),
.B(n_3),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_316),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_256),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_313),
.B(n_7),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_275),
.B(n_10),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_278),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_275),
.B(n_10),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_278),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_R g474 ( 
.A(n_257),
.B(n_92),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_318),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_324),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_246),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_213),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_219),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_261),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_11),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_327),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_329),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_265),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_217),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_266),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_229),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_267),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_276),
.B(n_12),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_230),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_330),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_247),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_251),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_253),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_276),
.B(n_18),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_268),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_269),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_271),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_280),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_331),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_246),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_281),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_300),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_310),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_270),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_272),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_218),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_273),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_259),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_274),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_323),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_325),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_277),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_340),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_343),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_349),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_355),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_246),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_334),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_361),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_218),
.Y(n_521)
);

BUFx6f_ASAP7_75t_SL g522 ( 
.A(n_260),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_486),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_477),
.B(n_260),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_348),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_506),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_462),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_466),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_468),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_419),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_452),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_416),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_L g545 ( 
.A(n_426),
.B(n_396),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_518),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_432),
.B(n_226),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_435),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_453),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_417),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_459),
.B(n_348),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_436),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_454),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_431),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_437),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_445),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_467),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_480),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_438),
.B(n_209),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_458),
.B(n_373),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_479),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_490),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_449),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_473),
.B(n_385),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_484),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_492),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_488),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_423),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_493),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_498),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_481),
.B(n_373),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_470),
.A2(n_221),
.B(n_215),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_471),
.B(n_284),
.Y(n_582)
);

BUFx2_ASAP7_75t_SL g583 ( 
.A(n_496),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_497),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_499),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_464),
.B(n_259),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_481),
.A2(n_228),
.B(n_224),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_503),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_504),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_439),
.B(n_234),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_505),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_441),
.B(n_284),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_511),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_508),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_R g597 ( 
.A(n_418),
.B(n_210),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_512),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_442),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_510),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_513),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_444),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_R g604 ( 
.A(n_425),
.B(n_279),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_425),
.B(n_260),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_446),
.B(n_235),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_455),
.B(n_236),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_539),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_527),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_527),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_576),
.B(n_421),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_546),
.B(n_430),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_576),
.B(n_489),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_586),
.B(n_469),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_SL g622 ( 
.A(n_608),
.B(n_424),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_586),
.A2(n_433),
.B1(n_491),
.B2(n_520),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_586),
.B(n_259),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_540),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_576),
.B(n_495),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_608),
.B(n_422),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_549),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_608),
.A2(n_305),
.B1(n_326),
.B2(n_356),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_548),
.A2(n_482),
.B1(n_430),
.B2(n_520),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_569),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_422),
.Y(n_635)
);

INVx4_ASAP7_75t_SL g636 ( 
.A(n_580),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_549),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_569),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_554),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_597),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_554),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_541),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_580),
.B(n_259),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_527),
.B(n_245),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_531),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_531),
.B(n_456),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_531),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_580),
.B(n_259),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_541),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_605),
.A2(n_456),
.B1(n_521),
.B2(n_485),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_580),
.B(n_434),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_541),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_529),
.B(n_434),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_582),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_529),
.B(n_440),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_440),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_546),
.B(n_485),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_552),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_561),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_529),
.B(n_447),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_447),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_604),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_572),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_526),
.A2(n_491),
.B1(n_451),
.B2(n_517),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_553),
.A2(n_581),
.B1(n_326),
.B2(n_356),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_553),
.B(n_448),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_553),
.B(n_448),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_524),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_572),
.B(n_465),
.C(n_451),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_581),
.B(n_305),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_541),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_523),
.A2(n_353),
.B1(n_342),
.B2(n_457),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_603),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_603),
.B(n_521),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_545),
.B(n_465),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_530),
.A2(n_369),
.B1(n_374),
.B2(n_362),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_550),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_582),
.B(n_475),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_603),
.B(n_475),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_545),
.B(n_476),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_552),
.B(n_463),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_525),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_562),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_543),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_587),
.B(n_476),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_568),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_603),
.B(n_482),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_603),
.B(n_483),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_525),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_568),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_578),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_603),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_528),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_483),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_555),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_536),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_551),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_592),
.B(n_500),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_592),
.B(n_500),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_581),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_581),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_592),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_579),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_570),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_591),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_532),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_532),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_535),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_592),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_606),
.B(n_514),
.Y(n_726)
);

AND2x6_ASAP7_75t_L g727 ( 
.A(n_606),
.B(n_250),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_535),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_606),
.B(n_515),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_535),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_591),
.Y(n_732)
);

INVx4_ASAP7_75t_SL g733 ( 
.A(n_559),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_595),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_589),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_595),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_606),
.A2(n_517),
.B1(n_516),
.B2(n_515),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_537),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_589),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_607),
.B(n_516),
.C(n_507),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_563),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_607),
.B(n_258),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_607),
.B(n_501),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_564),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_589),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_560),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_537),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_559),
.B(n_589),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_594),
.A2(n_522),
.B1(n_501),
.B2(n_405),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_537),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_573),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_598),
.B(n_522),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_588),
.A2(n_367),
.B1(n_397),
.B2(n_366),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_571),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_588),
.B(n_263),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_598),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_538),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_594),
.B(n_264),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_635),
.B(n_630),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_649),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_666),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_635),
.B(n_538),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_757),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_642),
.B(n_557),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_630),
.B(n_557),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_625),
.A2(n_367),
.B1(n_398),
.B2(n_411),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_757),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_636),
.B(n_557),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_657),
.B(n_210),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_708),
.B(n_538),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_708),
.B(n_565),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_649),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_688),
.Y(n_775)
);

INVxp33_ASAP7_75t_L g776 ( 
.A(n_664),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_624),
.B(n_622),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_670),
.B(n_677),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_625),
.A2(n_394),
.B1(n_401),
.B2(n_339),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_679),
.B(n_211),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_211),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_622),
.B(n_557),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_680),
.B(n_288),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_668),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_685),
.B(n_575),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_675),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_687),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_678),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_661),
.B(n_212),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_620),
.A2(n_368),
.B(n_298),
.C(n_590),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_672),
.B(n_294),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_678),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_693),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_672),
.B(n_297),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_672),
.B(n_301),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_659),
.B(n_212),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_636),
.B(n_364),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_680),
.A2(n_237),
.B1(n_346),
.B2(n_296),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_720),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_692),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_659),
.B(n_214),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_672),
.B(n_306),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_672),
.B(n_307),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_671),
.B(n_584),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_692),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_620),
.A2(n_599),
.B(n_590),
.C(n_585),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_618),
.B(n_308),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_627),
.B(n_312),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_609),
.B(n_322),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_684),
.B(n_593),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_701),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_684),
.A2(n_315),
.B1(n_283),
.B2(n_289),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_615),
.B(n_335),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_701),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_633),
.B(n_596),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_715),
.A2(n_336),
.B(n_382),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_674),
.A2(n_359),
.B(n_403),
.C(n_406),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_694),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_697),
.B(n_583),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_698),
.Y(n_820)
);

AND2x6_ASAP7_75t_SL g821 ( 
.A(n_617),
.B(n_360),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_662),
.B(n_669),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_706),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_616),
.B(n_626),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_628),
.B(n_372),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_702),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_629),
.B(n_375),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_704),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_718),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_712),
.B(n_214),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_662),
.B(n_220),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_707),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_631),
.B(n_637),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_674),
.A2(n_377),
.B(n_400),
.C(n_414),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_695),
.B(n_583),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_667),
.B(n_574),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_714),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_710),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_682),
.B(n_574),
.C(n_577),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_641),
.B(n_379),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_650),
.B(n_363),
.C(n_365),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_725),
.A2(n_599),
.B(n_590),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_746),
.Y(n_844)
);

NOR2x1p5_ASAP7_75t_L g845 ( 
.A(n_691),
.B(n_223),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_636),
.B(n_364),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_643),
.B(n_585),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_647),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_651),
.B(n_585),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_720),
.B(n_364),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_669),
.B(n_220),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_676),
.B(n_225),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_634),
.B(n_640),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_660),
.B(n_599),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_623),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_729),
.B(n_225),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_L g857 ( 
.A(n_740),
.B(n_223),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_719),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_746),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_743),
.A2(n_328),
.B1(n_358),
.B2(n_413),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_737),
.B(n_232),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_689),
.B(n_700),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_721),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_650),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_732),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_690),
.B(n_232),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_676),
.B(n_238),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_689),
.B(n_577),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_756),
.A2(n_408),
.B(n_601),
.C(n_602),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_700),
.B(n_290),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_735),
.B(n_364),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_713),
.B(n_227),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_734),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

INVx8_ASAP7_75t_L g875 ( 
.A(n_759),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_713),
.A2(n_354),
.B1(n_357),
.B2(n_351),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_611),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_759),
.B(n_727),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_690),
.B(n_238),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_726),
.A2(n_371),
.B1(n_350),
.B2(n_345),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_665),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_623),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_726),
.B(n_239),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_699),
.B(n_227),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_722),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_722),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_686),
.B(n_239),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_656),
.B(n_370),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_735),
.B(n_291),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_723),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_612),
.B(n_648),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_723),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_696),
.B(n_302),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_754),
.A2(n_344),
.B(n_341),
.C(n_338),
.Y(n_894)
);

BUFx6f_ASAP7_75t_SL g895 ( 
.A(n_656),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_739),
.B(n_304),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_647),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_623),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_699),
.A2(n_337),
.B1(n_332),
.B2(n_314),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_656),
.B(n_240),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_614),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_655),
.B(n_242),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_632),
.A2(n_364),
.B1(n_240),
.B2(n_413),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_739),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_745),
.B(n_319),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_358),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_619),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_652),
.B(n_242),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_745),
.B(n_243),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_647),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_614),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_754),
.B(n_243),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_619),
.B(n_381),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_621),
.B(n_646),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_638),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_621),
.B(n_381),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_638),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_639),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_646),
.B(n_383),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_639),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_653),
.B(n_383),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_653),
.B(n_384),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_759),
.B(n_384),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_759),
.B(n_388),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_742),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_759),
.B(n_388),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_828),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_762),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_762),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_761),
.B(n_715),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_778),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_798),
.A2(n_750),
.B(n_753),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_823),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_816),
.A2(n_756),
.B(n_717),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_862),
.A2(n_717),
.B(n_749),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_864),
.B(n_741),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_SL g937 ( 
.A1(n_817),
.A2(n_835),
.B(n_894),
.C(n_791),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_842),
.B(n_744),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_868),
.A2(n_634),
.B(n_640),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_777),
.A2(n_742),
.B(n_632),
.C(n_644),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_822),
.A2(n_644),
.B(n_758),
.C(n_730),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_819),
.B(n_711),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_822),
.A2(n_758),
.B(n_724),
.C(n_728),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_778),
.B(n_752),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_877),
.Y(n_945)
);

BUFx4f_ASAP7_75t_L g946 ( 
.A(n_836),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_783),
.A2(n_683),
.B(n_705),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_783),
.A2(n_751),
.B(n_748),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_828),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_895),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_774),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_823),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_789),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_781),
.B(n_727),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_781),
.B(n_727),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_914),
.A2(n_610),
.B(n_658),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_787),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_878),
.A2(n_772),
.B(n_794),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_764),
.B(n_727),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_774),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_891),
.B(n_727),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_795),
.A2(n_610),
.B(n_658),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_797),
.A2(n_730),
.B(n_751),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_891),
.B(n_705),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_788),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_828),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_790),
.A2(n_738),
.B(n_703),
.C(n_654),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_912),
.A2(n_738),
.B(n_703),
.C(n_654),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_773),
.A2(n_681),
.B(n_658),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_807),
.A2(n_681),
.B(n_747),
.C(n_709),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_802),
.A2(n_610),
.B(n_716),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_803),
.A2(n_610),
.B(n_716),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_808),
.B(n_716),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_925),
.A2(n_405),
.B1(n_399),
.B2(n_393),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_806),
.A2(n_716),
.B(n_645),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_824),
.A2(n_645),
.B(n_393),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_870),
.A2(n_733),
.B(n_364),
.C(n_474),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_771),
.B(n_733),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_834),
.A2(n_645),
.B(n_399),
.Y(n_980)
);

NOR2x1p5_ASAP7_75t_SL g981 ( 
.A(n_792),
.B(n_364),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_771),
.B(n_733),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_810),
.B(n_687),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_847),
.A2(n_645),
.B(n_376),
.Y(n_984)
);

O2A1O1Ixp5_ASAP7_75t_L g985 ( 
.A1(n_846),
.A2(n_364),
.B(n_461),
.C(n_352),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_775),
.B(n_755),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_830),
.A2(n_755),
.B1(n_709),
.B2(n_392),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_881),
.B(n_731),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_849),
.A2(n_392),
.B(n_412),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_850),
.A2(n_352),
.B(n_387),
.C(n_21),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_900),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_887),
.A2(n_919),
.B(n_922),
.C(n_921),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_883),
.A2(n_352),
.B(n_387),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_837),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_765),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_854),
.A2(n_376),
.B(n_412),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_830),
.B(n_390),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_844),
.B(n_390),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_796),
.A2(n_395),
.B(n_410),
.C(n_409),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_799),
.A2(n_378),
.B(n_410),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_792),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_905),
.A2(n_378),
.B(n_409),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_844),
.A2(n_867),
.B1(n_832),
.B2(n_851),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_889),
.A2(n_386),
.B(n_402),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_769),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_885),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_885),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_890),
.A2(n_386),
.B(n_402),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_908),
.B(n_395),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_828),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_908),
.B(n_389),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_798),
.B(n_389),
.C(n_731),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_760),
.B(n_387),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_857),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_893),
.B(n_97),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_796),
.A2(n_731),
.B1(n_96),
.B2(n_100),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_859),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_845),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_850),
.A2(n_95),
.B(n_198),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_871),
.A2(n_896),
.B(n_843),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_801),
.A2(n_851),
.B(n_867),
.C(n_832),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_871),
.A2(n_202),
.B(n_196),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_763),
.B(n_19),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_890),
.A2(n_193),
.B(n_192),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_909),
.A2(n_183),
.B(n_181),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_789),
.B(n_20),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_784),
.B(n_20),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_859),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_892),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_800),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_892),
.A2(n_176),
.B(n_167),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_801),
.A2(n_159),
.B1(n_154),
.B2(n_144),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_786),
.B(n_22),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_821),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_859),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_800),
.A2(n_814),
.B(n_811),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_839),
.B(n_848),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_883),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_852),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_895),
.B(n_141),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_913),
.A2(n_130),
.B(n_124),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_907),
.B(n_116),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_805),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_793),
.B(n_24),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_805),
.A2(n_105),
.B(n_104),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_916),
.A2(n_30),
.B(n_31),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_897),
.B(n_31),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_818),
.B(n_38),
.Y(n_1048)
);

AO21x1_ASAP7_75t_L g1049 ( 
.A1(n_852),
.A2(n_39),
.B(n_42),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_910),
.B(n_42),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_780),
.B(n_43),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_820),
.B(n_43),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_814),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_904),
.A2(n_918),
.B(n_915),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_826),
.B(n_45),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_779),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_875),
.A2(n_46),
.B(n_47),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_886),
.A2(n_51),
.B(n_54),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_804),
.B(n_54),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_872),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_780),
.A2(n_56),
.B1(n_59),
.B2(n_62),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_884),
.B(n_56),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_SL g1063 ( 
.A(n_770),
.B(n_907),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_861),
.B(n_815),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_785),
.B(n_831),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_901),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_906),
.B(n_888),
.Y(n_1067)
);

AO32x2_ASAP7_75t_L g1068 ( 
.A1(n_855),
.A2(n_768),
.A3(n_779),
.B1(n_869),
.B2(n_902),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_911),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_856),
.A2(n_866),
.B(n_879),
.C(n_840),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_829),
.B(n_865),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_L g1072 ( 
.A1(n_923),
.A2(n_926),
.B(n_924),
.C(n_863),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_917),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_901),
.A2(n_918),
.B(n_915),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_833),
.A2(n_838),
.B(n_858),
.C(n_874),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_920),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_875),
.A2(n_841),
.B(n_827),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_873),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_812),
.B(n_880),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_768),
.B(n_809),
.Y(n_1080)
);

BUFx2_ASAP7_75t_SL g1081 ( 
.A(n_898),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_776),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_813),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_875),
.A2(n_825),
.B(n_907),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_767),
.B(n_766),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_907),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_876),
.B(n_899),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_782),
.A2(n_882),
.B1(n_770),
.B2(n_860),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_903),
.A2(n_761),
.B(n_822),
.C(n_778),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_903),
.B(n_765),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_828),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_761),
.B(n_778),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_761),
.A2(n_620),
.B(n_777),
.C(n_625),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_877),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_823),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_816),
.A2(n_853),
.B(n_862),
.Y(n_1096)
);

NAND2xp33_ASAP7_75t_L g1097 ( 
.A(n_862),
.B(n_672),
.Y(n_1097)
);

INVxp67_ASAP7_75t_SL g1098 ( 
.A(n_830),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_761),
.A2(n_783),
.B1(n_862),
.B2(n_620),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_816),
.A2(n_862),
.B(n_868),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_823),
.Y(n_1101)
);

AO32x2_ASAP7_75t_L g1102 ( 
.A1(n_925),
.A2(n_717),
.A3(n_715),
.B1(n_897),
.B2(n_848),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_843),
.A2(n_853),
.B(n_806),
.Y(n_1103)
);

INVx11_ASAP7_75t_L g1104 ( 
.A(n_895),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_761),
.B(n_778),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_823),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_816),
.A2(n_862),
.B(n_868),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_761),
.B(n_778),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_823),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_1099),
.A2(n_1003),
.A3(n_1089),
.B(n_1107),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_957),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_946),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1020),
.A2(n_970),
.B(n_1074),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_SL g1114 ( 
.A(n_927),
.B(n_1028),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1093),
.A2(n_930),
.B(n_935),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_931),
.B(n_1092),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1066),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_933),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1105),
.B(n_1108),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_952),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1096),
.A2(n_1097),
.B(n_958),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1100),
.A2(n_1107),
.A3(n_934),
.B(n_1051),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1020),
.A2(n_970),
.B(n_1074),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_942),
.B(n_944),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1036),
.A2(n_956),
.B(n_962),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_946),
.B(n_1067),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_945),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_934),
.A2(n_1100),
.B(n_939),
.Y(n_1128)
);

INVx6_ASAP7_75t_L g1129 ( 
.A(n_927),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1094),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_993),
.A2(n_1049),
.A3(n_935),
.B(n_941),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_928),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1021),
.B(n_1083),
.Y(n_1133)
);

OAI33xp33_ASAP7_75t_L g1134 ( 
.A1(n_1009),
.A2(n_1011),
.A3(n_1062),
.B1(n_987),
.B2(n_953),
.B3(n_1071),
.Y(n_1134)
);

BUFx12f_ASAP7_75t_L g1135 ( 
.A(n_1018),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1038),
.B(n_1090),
.Y(n_1136)
);

BUFx4f_ASAP7_75t_L g1137 ( 
.A(n_988),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1090),
.B(n_964),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_927),
.Y(n_1139)
);

BUFx2_ASAP7_75t_R g1140 ( 
.A(n_950),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1014),
.B(n_1078),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_988),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_959),
.A2(n_937),
.B(n_954),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1084),
.A2(n_976),
.B(n_947),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1104),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_986),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1072),
.A2(n_940),
.B(n_943),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_995),
.B(n_1005),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1064),
.B(n_936),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1082),
.B(n_1060),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1087),
.A2(n_1079),
.B(n_932),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1028),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_947),
.A2(n_948),
.B(n_1080),
.Y(n_1153)
);

AO21x1_ASAP7_75t_L g1154 ( 
.A1(n_1070),
.A2(n_1045),
.B(n_1016),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1006),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_991),
.B(n_1012),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_929),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_951),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_992),
.A2(n_1026),
.B(n_1065),
.C(n_1075),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_961),
.A2(n_955),
.B(n_982),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_978),
.A2(n_969),
.B(n_1077),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_939),
.A2(n_1077),
.B(n_1086),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_SL g1163 ( 
.A1(n_1061),
.A2(n_1056),
.B(n_983),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_938),
.B(n_949),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1098),
.A2(n_979),
.B(n_973),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_972),
.A2(n_973),
.B(n_974),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1050),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_997),
.B(n_998),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1037),
.B(n_949),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_988),
.B(n_1081),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1050),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1085),
.B(n_994),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_1013),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1028),
.B(n_971),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_999),
.B(n_1059),
.C(n_975),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1023),
.Y(n_1176)
);

NAND2x1_ASAP7_75t_SL g1177 ( 
.A(n_1088),
.B(n_1035),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1007),
.B(n_1109),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_985),
.A2(n_1106),
.B(n_1101),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_989),
.B(n_996),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_984),
.A2(n_1024),
.A3(n_1031),
.B(n_1046),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1027),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1039),
.A2(n_1022),
.B(n_1019),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1029),
.A2(n_1043),
.B(n_1053),
.Y(n_1184)
);

AND3x4_ASAP7_75t_L g1185 ( 
.A(n_1034),
.B(n_1015),
.C(n_1040),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_960),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_968),
.A2(n_1095),
.B(n_966),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_965),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1001),
.B(n_1030),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1069),
.B(n_1076),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1002),
.A2(n_1044),
.B(n_1048),
.C(n_1033),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1073),
.B(n_967),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_989),
.B(n_996),
.Y(n_1193)
);

AO21x1_ASAP7_75t_L g1194 ( 
.A1(n_1041),
.A2(n_1032),
.B(n_1046),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1025),
.A2(n_984),
.B(n_1091),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1000),
.B(n_1052),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1055),
.B(n_1047),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1004),
.B(n_967),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1010),
.A2(n_1017),
.B1(n_1091),
.B2(n_1042),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1010),
.A2(n_1017),
.B1(n_1042),
.B2(n_1057),
.Y(n_1200)
);

AO21x1_ASAP7_75t_L g1201 ( 
.A1(n_1041),
.A2(n_977),
.B(n_980),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_977),
.B(n_980),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1068),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1019),
.A2(n_1022),
.B1(n_1031),
.B2(n_1024),
.Y(n_1204)
);

AOI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1058),
.A2(n_981),
.B(n_1102),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_990),
.B(n_1102),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1102),
.B(n_1068),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1068),
.A2(n_1096),
.B(n_934),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_927),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_934),
.A2(n_1096),
.B(n_935),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_942),
.B(n_944),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1066),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1021),
.A2(n_1089),
.B(n_1093),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1096),
.A2(n_934),
.B(n_1100),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_931),
.B(n_1092),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_931),
.B(n_1092),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1099),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_942),
.B(n_944),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_931),
.B(n_1092),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1066),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_L g1221 ( 
.A1(n_1087),
.A2(n_761),
.B(n_816),
.C(n_1079),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_931),
.B(n_1092),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_927),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_931),
.B(n_1092),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_957),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_957),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1099),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1096),
.A2(n_816),
.B(n_862),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_933),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_927),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1021),
.A2(n_1049),
.B(n_1045),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_L g1232 ( 
.A(n_1021),
.B(n_761),
.C(n_1051),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1021),
.A2(n_761),
.B1(n_1108),
.B2(n_1105),
.C(n_931),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_931),
.B(n_1092),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_949),
.B(n_1035),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_933),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_933),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_945),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_934),
.A2(n_1096),
.B(n_935),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_934),
.A2(n_816),
.B(n_1100),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_945),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1099),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1099),
.A2(n_1003),
.A3(n_1089),
.B(n_1100),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_931),
.B(n_1092),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1021),
.A2(n_761),
.B(n_1089),
.C(n_931),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1096),
.A2(n_934),
.B(n_1100),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_945),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_931),
.B(n_1092),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_944),
.A2(n_761),
.B1(n_1051),
.B2(n_931),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_931),
.B(n_1092),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1021),
.B(n_761),
.C(n_1051),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1096),
.A2(n_934),
.B(n_1100),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1021),
.A2(n_1099),
.B(n_1003),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_931),
.B(n_1092),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1054),
.A2(n_963),
.B(n_1103),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1021),
.A2(n_761),
.B(n_1089),
.C(n_931),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1021),
.A2(n_761),
.B(n_1089),
.C(n_931),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1021),
.A2(n_761),
.B(n_1089),
.C(n_931),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1021),
.A2(n_761),
.B(n_1089),
.C(n_931),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1066),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1066),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1221),
.A2(n_1151),
.B(n_1256),
.C(n_1232),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1124),
.B(n_1211),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1150),
.B(n_1218),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_SL g1270 ( 
.A1(n_1248),
.A2(n_1264),
.B(n_1263),
.C(n_1262),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1135),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1226),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1252),
.A2(n_1215),
.B(n_1119),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1116),
.B(n_1242),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1228),
.A2(n_1143),
.B(n_1151),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1126),
.B(n_1171),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1141),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1258),
.A2(n_1175),
.B1(n_1233),
.B2(n_1134),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1117),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1145),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1127),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1148),
.Y(n_1282)
);

NOR2xp67_ASAP7_75t_L g1283 ( 
.A(n_1146),
.B(n_1130),
.Y(n_1283)
);

O2A1O1Ixp5_ASAP7_75t_L g1284 ( 
.A1(n_1154),
.A2(n_1194),
.B(n_1243),
.C(n_1227),
.Y(n_1284)
);

INVx3_ASAP7_75t_SL g1285 ( 
.A(n_1141),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1139),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1182),
.B(n_1167),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1148),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1119),
.B(n_1215),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1132),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1233),
.A2(n_1149),
.B1(n_1173),
.B2(n_1156),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1118),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1238),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1143),
.A2(n_1214),
.B(n_1249),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1142),
.B(n_1112),
.Y(n_1295)
);

OR2x4_ASAP7_75t_L g1296 ( 
.A(n_1163),
.B(n_1216),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1217),
.A2(n_1243),
.B(n_1227),
.C(n_1201),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1197),
.B(n_1176),
.Y(n_1298)
);

INVx3_ASAP7_75t_SL g1299 ( 
.A(n_1111),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1140),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1216),
.B(n_1219),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1214),
.A2(n_1249),
.B(n_1257),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1157),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1170),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1170),
.B(n_1225),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1222),
.B(n_1224),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1257),
.A2(n_1121),
.B(n_1162),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1224),
.B(n_1234),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1136),
.B(n_1234),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1136),
.B(n_1246),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_1250),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1261),
.A2(n_1217),
.B(n_1259),
.C(n_1254),
.Y(n_1313)
);

INVx3_ASAP7_75t_SL g1314 ( 
.A(n_1170),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1230),
.B(n_1223),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1120),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1180),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1139),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1246),
.B(n_1251),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1320)
);

INVx3_ASAP7_75t_SL g1321 ( 
.A(n_1129),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1251),
.B(n_1254),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1137),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1147),
.A2(n_1161),
.B(n_1153),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1259),
.B(n_1133),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1139),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1140),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1133),
.B(n_1138),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1128),
.A2(n_1115),
.B(n_1213),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1115),
.A2(n_1159),
.B(n_1153),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1169),
.B(n_1164),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1209),
.B(n_1129),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1165),
.A2(n_1241),
.B(n_1147),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1137),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1168),
.B(n_1138),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1155),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1203),
.A2(n_1185),
.B1(n_1237),
.B2(n_1236),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1209),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1241),
.A2(n_1208),
.B(n_1204),
.Y(n_1339)
);

BUFx4_ASAP7_75t_SL g1340 ( 
.A(n_1198),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1209),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1230),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1193),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1152),
.B(n_1230),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1229),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1208),
.A2(n_1204),
.B(n_1166),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1196),
.B(n_1110),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1191),
.B(n_1174),
.C(n_1161),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1230),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1192),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1206),
.A2(n_1187),
.B(n_1144),
.Y(n_1351)
);

BUFx2_ASAP7_75t_R g1352 ( 
.A(n_1192),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_L g1353 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1188),
.A2(n_1266),
.B1(n_1265),
.B2(n_1186),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1158),
.B(n_1212),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1184),
.B(n_1200),
.C(n_1179),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1231),
.A2(n_1183),
.B1(n_1220),
.B2(n_1178),
.Y(n_1357)
);

OAI21xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1177),
.A2(n_1184),
.B(n_1206),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_1125),
.Y(n_1359)
);

BUFx5_ASAP7_75t_L g1360 ( 
.A(n_1160),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1152),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1202),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1195),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1178),
.B(n_1189),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1110),
.B(n_1245),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1189),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1110),
.B(n_1245),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1114),
.B(n_1205),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1210),
.B(n_1240),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_SL g1370 ( 
.A1(n_1207),
.A2(n_1131),
.B(n_1181),
.C(n_1122),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1131),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1207),
.A2(n_1244),
.B1(n_1255),
.B2(n_1253),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1239),
.B(n_1247),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1260),
.A2(n_1122),
.B(n_1181),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1122),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1226),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1135),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1119),
.B(n_931),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1149),
.B(n_761),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1124),
.B(n_1211),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1119),
.B(n_931),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1140),
.Y(n_1382)
);

AO21x1_ASAP7_75t_L g1383 ( 
.A1(n_1151),
.A2(n_1021),
.B(n_1003),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1235),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1126),
.B(n_1171),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1148),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1139),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1228),
.A2(n_1096),
.B(n_1100),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1139),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1149),
.B(n_761),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1124),
.B(n_1211),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1126),
.B(n_1171),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1139),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1226),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1228),
.A2(n_1096),
.B(n_1100),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1148),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_1012),
.B1(n_1051),
.B2(n_761),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1135),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1124),
.B(n_1211),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1148),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1190),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1117),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1226),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1228),
.A2(n_1096),
.B(n_1100),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1119),
.B(n_931),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1117),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1248),
.A2(n_761),
.B(n_1021),
.C(n_1051),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1190),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1119),
.B(n_931),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1119),
.B(n_931),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1135),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1242),
.Y(n_1412)
);

INVx3_ASAP7_75t_SL g1413 ( 
.A(n_1145),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1228),
.A2(n_1096),
.B(n_1100),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1242),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1119),
.B(n_931),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1235),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1235),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1139),
.Y(n_1419)
);

BUFx4_ASAP7_75t_SL g1420 ( 
.A(n_1111),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1217),
.A2(n_1051),
.B(n_761),
.C(n_1021),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1148),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1232),
.A2(n_1012),
.B1(n_1051),
.B2(n_761),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1119),
.B(n_931),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1235),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1149),
.B(n_761),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1127),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1269),
.B(n_1274),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1342),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1272),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1366),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1376),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1379),
.A2(n_1390),
.B1(n_1426),
.B2(n_1343),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1348),
.A2(n_1375),
.B1(n_1353),
.B2(n_1330),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1316),
.Y(n_1435)
);

BUFx10_ASAP7_75t_L g1436 ( 
.A(n_1300),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1268),
.B(n_1380),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1336),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1397),
.A2(n_1423),
.B1(n_1273),
.B2(n_1296),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1391),
.B(n_1399),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1345),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1412),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1344),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1294),
.A2(n_1308),
.B(n_1302),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1327),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1344),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1279),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1412),
.Y(n_1448)
);

OAI22x1_ASAP7_75t_L g1449 ( 
.A1(n_1320),
.A2(n_1307),
.B1(n_1309),
.B2(n_1305),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1342),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1298),
.B(n_1310),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_SL g1452 ( 
.A(n_1407),
.B(n_1421),
.C(n_1291),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1293),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1342),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1288),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1290),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1359),
.A2(n_1374),
.B(n_1346),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1415),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1312),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1303),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1319),
.B(n_1322),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1312),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1313),
.A2(n_1267),
.B(n_1297),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1402),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1406),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1401),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1408),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1355),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1354),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1354),
.Y(n_1470)
);

BUFx4f_ASAP7_75t_L g1471 ( 
.A(n_1280),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1350),
.Y(n_1472)
);

BUFx2_ASAP7_75t_R g1473 ( 
.A(n_1382),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1409),
.A2(n_1296),
.B1(n_1289),
.B2(n_1301),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1350),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1335),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1333),
.A2(n_1275),
.B(n_1404),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1394),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1311),
.B(n_1287),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1276),
.B(n_1385),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1413),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_SL g1482 ( 
.A1(n_1325),
.A2(n_1383),
.B(n_1328),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1320),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1364),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1351),
.A2(n_1363),
.B(n_1388),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1289),
.B(n_1301),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1317),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1273),
.A2(n_1278),
.B1(n_1424),
.B2(n_1416),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1276),
.B(n_1385),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1332),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1325),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1331),
.B(n_1323),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1328),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1347),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1347),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1395),
.A2(n_1414),
.B(n_1363),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1284),
.A2(n_1339),
.B(n_1351),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1378),
.A2(n_1410),
.B1(n_1424),
.B2(n_1381),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1337),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1317),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1277),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1337),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1286),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1392),
.B(n_1282),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1392),
.B(n_1386),
.Y(n_1505)
);

BUFx8_ASAP7_75t_L g1506 ( 
.A(n_1396),
.Y(n_1506)
);

CKINVDCx11_ASAP7_75t_R g1507 ( 
.A(n_1299),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1331),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1348),
.A2(n_1329),
.B(n_1357),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1285),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1286),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1400),
.B(n_1422),
.Y(n_1512)
);

INVx11_ASAP7_75t_L g1513 ( 
.A(n_1420),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1367),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1371),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1360),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1306),
.B(n_1418),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_R g1518 ( 
.A(n_1403),
.B(n_1334),
.Y(n_1518)
);

BUFx2_ASAP7_75t_R g1519 ( 
.A(n_1271),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1362),
.A2(n_1370),
.B(n_1372),
.Y(n_1520)
);

BUFx8_ASAP7_75t_L g1521 ( 
.A(n_1295),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1324),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1270),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1378),
.A2(n_1416),
.B1(n_1381),
.B2(n_1405),
.Y(n_1524)
);

BUFx2_ASAP7_75t_R g1525 ( 
.A(n_1377),
.Y(n_1525)
);

BUFx10_ASAP7_75t_L g1526 ( 
.A(n_1403),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1405),
.A2(n_1410),
.B1(n_1324),
.B2(n_1356),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1415),
.B(n_1283),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1286),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1365),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1295),
.B(n_1306),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1321),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1373),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1281),
.B(n_1427),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1361),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1356),
.A2(n_1358),
.B1(n_1306),
.B2(n_1352),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1373),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1373),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1358),
.A2(n_1340),
.B1(n_1368),
.B2(n_1411),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1314),
.B(n_1304),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1318),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1369),
.A2(n_1425),
.B(n_1384),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1318),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1318),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1326),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1425),
.A2(n_1418),
.B(n_1417),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1417),
.B(n_1332),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1315),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1398),
.A2(n_1315),
.B1(n_1349),
.B2(n_1341),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1326),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1326),
.A2(n_1338),
.B1(n_1341),
.B2(n_1387),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1338),
.A2(n_1341),
.B1(n_1387),
.B2(n_1389),
.Y(n_1552)
);

BUFx10_ASAP7_75t_L g1553 ( 
.A(n_1387),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1393),
.B(n_1419),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1393),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1274),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1379),
.A2(n_761),
.B1(n_1099),
.B2(n_1051),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1292),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1292),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1312),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1293),
.Y(n_1561)
);

INVx5_ASAP7_75t_L g1562 ( 
.A(n_1342),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1289),
.B(n_1301),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1366),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1342),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1268),
.B(n_1380),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1288),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1272),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1292),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1409),
.A2(n_1252),
.B1(n_761),
.B2(n_1092),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1331),
.B(n_1320),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1292),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1342),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1292),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1292),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1530),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1522),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1514),
.B(n_1494),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1517),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1507),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1490),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1495),
.B(n_1434),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1486),
.B(n_1498),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1498),
.B(n_1451),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1472),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1515),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1475),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1477),
.A2(n_1452),
.B(n_1509),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1557),
.A2(n_1570),
.B(n_1439),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1487),
.B(n_1500),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1533),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1457),
.A2(n_1485),
.B(n_1496),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1434),
.B(n_1487),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1490),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1500),
.B(n_1499),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1537),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1542),
.B(n_1490),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1557),
.A2(n_1433),
.B(n_1463),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1537),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1444),
.A2(n_1520),
.B(n_1527),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1538),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1538),
.Y(n_1604)
);

BUFx2_ASAP7_75t_R g1605 ( 
.A(n_1445),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1437),
.Y(n_1606)
);

BUFx4f_ASAP7_75t_SL g1607 ( 
.A(n_1568),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1556),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1542),
.B(n_1517),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1444),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1431),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1517),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1562),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1474),
.B(n_1563),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1431),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1521),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1462),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1520),
.A2(n_1482),
.B(n_1516),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1497),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1488),
.A2(n_1469),
.B(n_1470),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1440),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1566),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1442),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1493),
.B(n_1491),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1497),
.A2(n_1546),
.B(n_1523),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1435),
.A2(n_1575),
.B(n_1574),
.Y(n_1629)
);

NAND2x1p5_ASAP7_75t_L g1630 ( 
.A(n_1497),
.B(n_1546),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1564),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1632)
);

AO22x1_ASAP7_75t_L g1633 ( 
.A1(n_1521),
.A2(n_1466),
.B1(n_1467),
.B2(n_1468),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1449),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1438),
.B(n_1441),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1448),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1462),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1563),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1458),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1483),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1569),
.B(n_1572),
.Y(n_1642)
);

OAI33xp33_ASAP7_75t_L g1643 ( 
.A1(n_1447),
.A2(n_1460),
.A3(n_1456),
.B1(n_1465),
.B2(n_1464),
.B3(n_1528),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1508),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1488),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1433),
.B(n_1504),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1430),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1571),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1547),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1548),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1571),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1571),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1539),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1539),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1552),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1462),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1531),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1552),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1536),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1455),
.A2(n_1567),
.B1(n_1512),
.B2(n_1492),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1492),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1549),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1541),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1429),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1549),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1562),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1544),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1545),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1513),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1550),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1521),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_SL g1675 ( 
.A(n_1617),
.B(n_1562),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1587),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1577),
.B(n_1505),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1599),
.B(n_1609),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1584),
.B(n_1480),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1587),
.Y(n_1680)
);

BUFx2_ASAP7_75t_SL g1681 ( 
.A(n_1619),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1577),
.B(n_1540),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1632),
.B(n_1551),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1609),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1609),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1622),
.A2(n_1554),
.B(n_1534),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1609),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1614),
.B(n_1429),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1614),
.B(n_1446),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1638),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1629),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1623),
.B(n_1429),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1629),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1591),
.B(n_1454),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1623),
.B(n_1450),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1629),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1634),
.Y(n_1697)
);

INVxp67_ASAP7_75t_SL g1698 ( 
.A(n_1628),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1591),
.B(n_1535),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1622),
.B(n_1511),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1600),
.A2(n_1519),
.B1(n_1525),
.B2(n_1471),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1579),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1576),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1621),
.B(n_1511),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1621),
.B(n_1511),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1621),
.B(n_1511),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1589),
.B(n_1543),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1590),
.A2(n_1660),
.B1(n_1645),
.B2(n_1612),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1589),
.B(n_1543),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1589),
.B(n_1543),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1623),
.B(n_1573),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1671),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1598),
.B(n_1529),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1634),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1580),
.B(n_1471),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1601),
.B(n_1510),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1601),
.B(n_1603),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1630),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1604),
.B(n_1501),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1578),
.B(n_1573),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1617),
.B(n_1561),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1578),
.B(n_1450),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1645),
.B(n_1503),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1682),
.B(n_1608),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1682),
.B(n_1610),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1708),
.B(n_1667),
.C(n_1664),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1708),
.B(n_1667),
.C(n_1664),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1586),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1677),
.B(n_1588),
.Y(n_1731)
);

NOR3xp33_ASAP7_75t_L g1732 ( 
.A(n_1701),
.B(n_1633),
.C(n_1643),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1677),
.B(n_1583),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1701),
.A2(n_1660),
.B1(n_1654),
.B2(n_1653),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1716),
.B(n_1624),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1688),
.B(n_1583),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1697),
.A2(n_1654),
.B1(n_1653),
.B2(n_1615),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1683),
.B(n_1661),
.C(n_1633),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1683),
.B(n_1646),
.C(n_1585),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1684),
.B(n_1595),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1697),
.A2(n_1615),
.B1(n_1652),
.B2(n_1659),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1687),
.B(n_1630),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1688),
.B(n_1640),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1707),
.A2(n_1710),
.B(n_1709),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1687),
.B(n_1630),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1679),
.B(n_1592),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1700),
.B(n_1602),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1679),
.B(n_1689),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1700),
.B(n_1685),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_1655),
.C(n_1658),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1689),
.B(n_1592),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1689),
.B(n_1699),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1715),
.A2(n_1659),
.B(n_1673),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1626),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1700),
.B(n_1602),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1685),
.B(n_1602),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1715),
.A2(n_1625),
.B1(n_1606),
.B2(n_1636),
.C(n_1655),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1723),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1722),
.A2(n_1673),
.B(n_1658),
.Y(n_1760)
);

OAI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1724),
.A2(n_1615),
.B(n_1597),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1721),
.B(n_1635),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1723),
.B(n_1690),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1685),
.B(n_1707),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1722),
.B(n_1649),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1635),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1718),
.B(n_1639),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1717),
.A2(n_1619),
.B1(n_1662),
.B2(n_1597),
.C(n_1674),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1718),
.B(n_1639),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1717),
.A2(n_1619),
.B1(n_1662),
.B2(n_1605),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1709),
.B(n_1642),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1698),
.A2(n_1594),
.B(n_1611),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1709),
.B(n_1642),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1774)
);

NAND2x1_ASAP7_75t_L g1775 ( 
.A(n_1678),
.B(n_1710),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1724),
.B(n_1644),
.C(n_1641),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1676),
.B(n_1650),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1675),
.A2(n_1582),
.B(n_1596),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1676),
.B(n_1650),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1691),
.B(n_1696),
.C(n_1693),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1680),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1692),
.A2(n_1672),
.B1(n_1669),
.B2(n_1670),
.C(n_1627),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1692),
.A2(n_1672),
.B1(n_1669),
.B2(n_1670),
.C(n_1627),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1680),
.B(n_1713),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1704),
.B(n_1648),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1713),
.B(n_1613),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1713),
.B(n_1618),
.Y(n_1789)
);

OAI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1695),
.A2(n_1644),
.B(n_1631),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1783),
.B(n_1686),
.Y(n_1791)
);

AND2x4_ASAP7_75t_SL g1792 ( 
.A(n_1732),
.B(n_1678),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1764),
.B(n_1750),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1778),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1748),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1781),
.B(n_1719),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1749),
.B(n_1686),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1786),
.B(n_1686),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1729),
.B(n_1686),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1771),
.B(n_1691),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1771),
.B(n_1693),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1780),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1773),
.B(n_1678),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1756),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1773),
.B(n_1696),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1725),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1726),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1727),
.B(n_1720),
.C(n_1665),
.Y(n_1808)
);

NAND4xp25_ASAP7_75t_L g1809 ( 
.A(n_1728),
.B(n_1453),
.C(n_1561),
.D(n_1532),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1745),
.B(n_1678),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1775),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1775),
.B(n_1678),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1741),
.B(n_1678),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1737),
.B(n_1733),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1743),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1757),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1735),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1784),
.B(n_1703),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1757),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1743),
.B(n_1719),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1753),
.B(n_1695),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1746),
.B(n_1705),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1746),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1774),
.B(n_1719),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1735),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1774),
.B(n_1719),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1782),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1766),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1772),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1767),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1787),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1785),
.B(n_1703),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1759),
.B(n_1706),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1769),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1752),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1776),
.B(n_1706),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1763),
.B(n_1711),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1788),
.Y(n_1839)
);

AOI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1809),
.A2(n_1740),
.B(n_1739),
.C(n_1770),
.Y(n_1840)
);

BUFx2_ASAP7_75t_SL g1841 ( 
.A(n_1796),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1794),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1822),
.Y(n_1843)
);

NOR2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1809),
.B(n_1581),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1796),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1794),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1799),
.B(n_1797),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1821),
.B(n_1789),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1799),
.B(n_1744),
.Y(n_1849)
);

AOI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1817),
.A2(n_1754),
.B(n_1712),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1810),
.B(n_1776),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1797),
.B(n_1730),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1826),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1762),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1798),
.B(n_1731),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1802),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1810),
.B(n_1765),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1802),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1806),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1807),
.B(n_1751),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1821),
.B(n_1747),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1807),
.B(n_1755),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1839),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1838),
.B(n_1765),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1839),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1838),
.B(n_1768),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1808),
.B(n_1758),
.C(n_1734),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1792),
.A2(n_1736),
.B1(n_1761),
.B2(n_1760),
.C(n_1738),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1798),
.B(n_1711),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1808),
.B(n_1777),
.C(n_1790),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1822),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1822),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1834),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1834),
.Y(n_1874)
);

NOR2xp67_ASAP7_75t_L g1875 ( 
.A(n_1826),
.B(n_1581),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1837),
.B(n_1702),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1800),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1830),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1837),
.B(n_1813),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1836),
.B(n_1714),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1836),
.B(n_1714),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1812),
.B(n_1675),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1812),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1800),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1853),
.B(n_1792),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1843),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1859),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1867),
.A2(n_1792),
.B1(n_1818),
.B2(n_1833),
.C(n_1831),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1870),
.A2(n_1812),
.B1(n_1651),
.B2(n_1742),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1852),
.B(n_1791),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1863),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1840),
.A2(n_1779),
.B(n_1607),
.C(n_1812),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1844),
.A2(n_1835),
.B1(n_1829),
.B2(n_1831),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1882),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1853),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1865),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1852),
.B(n_1791),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1882),
.B(n_1811),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1860),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1842),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1862),
.B(n_1829),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1846),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1864),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1856),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1866),
.B(n_1835),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1882),
.B(n_1811),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1858),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1850),
.A2(n_1868),
.B(n_1845),
.C(n_1875),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1880),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1843),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1854),
.B(n_1814),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1871),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1881),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1873),
.Y(n_1915)
);

NAND2x1_ASAP7_75t_L g1916 ( 
.A(n_1883),
.B(n_1779),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1849),
.A2(n_1833),
.B(n_1818),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1879),
.B(n_1813),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1857),
.A2(n_1651),
.B1(n_1814),
.B2(n_1820),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1879),
.B(n_1803),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1871),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1851),
.B(n_1803),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1849),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1861),
.B(n_1815),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_SL g1925 ( 
.A1(n_1874),
.A2(n_1430),
.B(n_1647),
.C(n_1481),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1872),
.Y(n_1926)
);

NAND2x1_ASAP7_75t_L g1927 ( 
.A(n_1883),
.B(n_1828),
.Y(n_1927)
);

AOI32xp33_ASAP7_75t_L g1928 ( 
.A1(n_1857),
.A2(n_1828),
.A3(n_1825),
.B1(n_1827),
.B2(n_1819),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1872),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1851),
.B(n_1823),
.Y(n_1930)
);

INVx5_ASAP7_75t_L g1931 ( 
.A(n_1900),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1927),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1922),
.B(n_1883),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1887),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1927),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1891),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1906),
.B(n_1847),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1896),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1901),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1904),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1899),
.B(n_1877),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1903),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1922),
.B(n_1876),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1895),
.B(n_1884),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1886),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1905),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1923),
.B(n_1847),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1910),
.B(n_1869),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1930),
.B(n_1876),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1888),
.B(n_1848),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1915),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1930),
.B(n_1855),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1918),
.B(n_1855),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1900),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1909),
.A2(n_1681),
.B1(n_1649),
.B2(n_1663),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1917),
.B(n_1815),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1918),
.B(n_1823),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1912),
.B(n_1902),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1920),
.B(n_1869),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1920),
.B(n_1820),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1909),
.B(n_1824),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1914),
.B(n_1890),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1886),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1893),
.B(n_1825),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1916),
.B(n_1481),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1908),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1889),
.A2(n_1651),
.B1(n_1681),
.B2(n_1649),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1916),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1926),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1931),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1934),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1955),
.A2(n_1885),
.B(n_1928),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1951),
.B(n_1925),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1969),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1954),
.Y(n_1975)
);

OAI222xp33_ASAP7_75t_L g1976 ( 
.A1(n_1955),
.A2(n_1919),
.B1(n_1894),
.B2(n_1907),
.C1(n_1898),
.C2(n_1892),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1940),
.B(n_1925),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1950),
.B(n_1924),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1961),
.B(n_1929),
.C(n_1913),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1934),
.Y(n_1980)
);

AND4x1_ASAP7_75t_L g1981 ( 
.A(n_1965),
.B(n_1907),
.C(n_1568),
.D(n_1478),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1943),
.B(n_1894),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1965),
.B(n_1894),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1964),
.A2(n_1898),
.B1(n_1827),
.B2(n_1825),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1931),
.B(n_1943),
.Y(n_1985)
);

OAI21xp33_ASAP7_75t_SL g1986 ( 
.A1(n_1932),
.A2(n_1897),
.B(n_1890),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1936),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_SL g1988 ( 
.A1(n_1967),
.A2(n_1898),
.B(n_1897),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1931),
.B(n_1911),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1931),
.A2(n_1819),
.B1(n_1816),
.B2(n_1832),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1941),
.A2(n_1518),
.B(n_1911),
.Y(n_1991)
);

OAI31xp33_ASAP7_75t_L g1992 ( 
.A1(n_1968),
.A2(n_1825),
.A3(n_1827),
.B(n_1921),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1958),
.A2(n_1944),
.B1(n_1942),
.B2(n_1938),
.C(n_1939),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_SL g1994 ( 
.A(n_1931),
.B(n_1473),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1933),
.A2(n_1827),
.B1(n_1913),
.B2(n_1921),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1936),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1937),
.B(n_1878),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1931),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1994),
.B(n_1968),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1974),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1973),
.B(n_1977),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1985),
.B(n_1949),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1975),
.B(n_1949),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1985),
.B(n_1933),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1993),
.B(n_1957),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1974),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1978),
.B(n_1957),
.Y(n_2008)
);

OAI21xp33_ASAP7_75t_SL g2009 ( 
.A1(n_1983),
.A2(n_1935),
.B(n_1932),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1971),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1983),
.B(n_1960),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1980),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1972),
.A2(n_1937),
.B1(n_1968),
.B2(n_1947),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1987),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1981),
.B(n_1960),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1996),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1991),
.B(n_1432),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1970),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1998),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1998),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1982),
.B(n_1938),
.Y(n_2021)
);

NAND4xp25_ASAP7_75t_L g2022 ( 
.A(n_2013),
.B(n_1984),
.C(n_1992),
.D(n_1979),
.Y(n_2022)
);

NAND4xp25_ASAP7_75t_L g2023 ( 
.A(n_2001),
.B(n_2003),
.C(n_2005),
.D(n_2015),
.Y(n_2023)
);

OAI21xp33_ASAP7_75t_L g2024 ( 
.A1(n_2002),
.A2(n_1986),
.B(n_1988),
.Y(n_2024)
);

AOI322xp5_ASAP7_75t_L g2025 ( 
.A1(n_2008),
.A2(n_1999),
.A3(n_2010),
.B1(n_2014),
.B2(n_2012),
.C1(n_2016),
.C2(n_2015),
.Y(n_2025)
);

OAI21xp5_ASAP7_75t_SL g2026 ( 
.A1(n_2017),
.A2(n_1976),
.B(n_1995),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_2018),
.B(n_1989),
.Y(n_2027)
);

AOI221x1_ASAP7_75t_L g2028 ( 
.A1(n_2018),
.A2(n_2020),
.B1(n_2019),
.B2(n_2016),
.C(n_2000),
.Y(n_2028)
);

AOI221x1_ASAP7_75t_L g2029 ( 
.A1(n_2019),
.A2(n_1989),
.B1(n_1939),
.B2(n_1946),
.C(n_1966),
.Y(n_2029)
);

OAI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_2009),
.A2(n_1947),
.B1(n_1935),
.B2(n_1990),
.C(n_1942),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2011),
.A2(n_1956),
.B1(n_1966),
.B2(n_1946),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2002),
.A2(n_1997),
.B(n_1969),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_2011),
.A2(n_1952),
.B1(n_1953),
.B2(n_1959),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_2004),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_2021),
.B(n_1432),
.Y(n_2035)
);

NAND2x1p5_ASAP7_75t_L g2036 ( 
.A(n_2027),
.B(n_1532),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_2033),
.B(n_2004),
.Y(n_2037)
);

NAND3xp33_ASAP7_75t_SL g2038 ( 
.A(n_2026),
.B(n_2020),
.C(n_2006),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2034),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2025),
.A2(n_2007),
.B(n_1962),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2028),
.Y(n_2041)
);

OAI322xp33_ASAP7_75t_L g2042 ( 
.A1(n_2031),
.A2(n_1997),
.A3(n_1962),
.B1(n_1963),
.B2(n_1945),
.C1(n_1948),
.C2(n_1952),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2022),
.A2(n_1963),
.B1(n_1945),
.B2(n_1953),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2029),
.Y(n_2044)
);

NOR3xp33_ASAP7_75t_L g2045 ( 
.A(n_2023),
.B(n_1507),
.C(n_1445),
.Y(n_2045)
);

NOR2x1_ASAP7_75t_L g2046 ( 
.A(n_2035),
.B(n_1453),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2024),
.B(n_1959),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2030),
.A2(n_2032),
.B1(n_1948),
.B2(n_1878),
.Y(n_2048)
);

NOR4xp25_ASAP7_75t_L g2049 ( 
.A(n_2041),
.B(n_1459),
.C(n_1560),
.D(n_1637),
.Y(n_2049)
);

NAND3xp33_ASAP7_75t_L g2050 ( 
.A(n_2040),
.B(n_1478),
.C(n_1555),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2038),
.A2(n_2045),
.B1(n_2037),
.B2(n_2044),
.Y(n_2051)
);

NOR2xp67_ASAP7_75t_L g2052 ( 
.A(n_2048),
.B(n_1620),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_2039),
.B(n_2047),
.C(n_2046),
.Y(n_2053)
);

OAI211xp5_ASAP7_75t_SL g2054 ( 
.A1(n_2043),
.A2(n_1555),
.B(n_1478),
.C(n_1620),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_2036),
.A2(n_2042),
.B1(n_1637),
.B2(n_1656),
.C(n_1819),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2051),
.B(n_2036),
.Y(n_2056)
);

NOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2050),
.B(n_1526),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2054),
.A2(n_1436),
.B1(n_1656),
.B2(n_1526),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2053),
.A2(n_1436),
.B1(n_1820),
.B2(n_1830),
.Y(n_2059)
);

INVxp67_ASAP7_75t_SL g2060 ( 
.A(n_2052),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_2055),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2049),
.B(n_1816),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2062),
.B(n_1824),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2057),
.B(n_1565),
.C(n_1506),
.D(n_1616),
.Y(n_2064)
);

OAI321xp33_ASAP7_75t_L g2065 ( 
.A1(n_2056),
.A2(n_2059),
.A3(n_2060),
.B1(n_2058),
.B2(n_2061),
.C(n_1720),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2058),
.A2(n_1820),
.B1(n_1506),
.B2(n_1816),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2062),
.B(n_1801),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2060),
.B(n_1793),
.Y(n_2068)
);

XNOR2xp5_ASAP7_75t_L g2069 ( 
.A(n_2068),
.B(n_1506),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2063),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2067),
.Y(n_2071)
);

XNOR2xp5_ASAP7_75t_L g2072 ( 
.A(n_2064),
.B(n_1665),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2070),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2073),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2074),
.A2(n_2065),
.B(n_2069),
.Y(n_2075)
);

OAI21xp33_ASAP7_75t_L g2076 ( 
.A1(n_2074),
.A2(n_2066),
.B(n_2071),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2075),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2076),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2078),
.A2(n_2072),
.B1(n_1565),
.B2(n_1503),
.C(n_1830),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_2077),
.A2(n_1805),
.B(n_1801),
.Y(n_2080)
);

OA21x2_ASAP7_75t_L g2081 ( 
.A1(n_2079),
.A2(n_2080),
.B(n_1805),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2081),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_R g2083 ( 
.A1(n_2082),
.A2(n_1553),
.B1(n_1503),
.B2(n_1804),
.C(n_1795),
.Y(n_2083)
);

AOI211xp5_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_1503),
.B(n_1666),
.C(n_1668),
.Y(n_2084)
);


endmodule