module fake_jpeg_9595_n_81 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx11_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_1),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_3),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_43),
.C(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_36),
.B1(n_19),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_2),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_65),
.B(n_66),
.C(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_64),
.B1(n_15),
.B2(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_10),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_58),
.C(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_62),
.Y(n_74)
);

OAI322xp33_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_68),
.A3(n_62),
.B1(n_69),
.B2(n_71),
.C1(n_55),
.C2(n_57),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_24),
.C(n_25),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_27),
.B(n_29),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_30),
.B(n_31),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_32),
.B(n_33),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_80),
.Y(n_81)
);


endmodule