module fake_jpeg_21757_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx4_ASAP7_75t_SL g9 ( 
.A(n_3),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_17),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_4),
.B1(n_5),
.B2(n_14),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_6),
.C(n_2),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_2),
.B(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_7),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_22),
.B(n_9),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_8),
.B1(n_7),
.B2(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_26),
.B1(n_30),
.B2(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_22),
.B1(n_15),
.B2(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_37),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_27),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B(n_36),
.Y(n_45)
);

A2O1A1O1Ixp25_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_39),
.B(n_34),
.C(n_33),
.D(n_25),
.Y(n_47)
);

OAI221xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_46),
.B1(n_38),
.B2(n_18),
.C(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_31),
.Y(n_49)
);


endmodule