module fake_netlist_5_1384_n_400 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_58, n_36, n_25, n_53, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_56, n_51, n_11, n_17, n_19, n_57, n_7, n_37, n_59, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_3, n_49, n_52, n_60, n_6, n_39, n_400);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_58;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_56;
input n_51;
input n_11;
input n_17;
input n_19;
input n_57;
input n_7;
input n_37;
input n_59;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_3;
input n_49;
input n_52;
input n_60;
input n_6;
input n_39;

output n_400;

wire n_137;
wire n_294;
wire n_318;
wire n_380;
wire n_82;
wire n_194;
wire n_316;
wire n_389;
wire n_248;
wire n_124;
wire n_86;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_61;
wire n_376;
wire n_127;
wire n_75;
wire n_235;
wire n_226;
wire n_74;
wire n_353;
wire n_351;
wire n_367;
wire n_397;
wire n_111;
wire n_155;
wire n_116;
wire n_284;
wire n_245;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_368;
wire n_321;
wire n_292;
wire n_100;
wire n_212;
wire n_385;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_373;
wire n_67;
wire n_307;
wire n_87;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_375;
wire n_301;
wire n_68;
wire n_93;
wire n_186;
wire n_134;
wire n_191;
wire n_63;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_325;
wire n_132;
wire n_90;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_94;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_95;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_72;
wire n_104;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_313;
wire n_88;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_65;
wire n_78;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_98;
wire n_361;
wire n_363;
wire n_197;
wire n_107;
wire n_69;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_80;
wire n_73;
wire n_277;
wire n_92;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_84;
wire n_130;
wire n_322;
wire n_258;
wire n_79;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_112;
wire n_85;
wire n_239;
wire n_310;
wire n_76;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_102;
wire n_77;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_81;
wire n_118;
wire n_279;
wire n_70;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_345;
wire n_210;
wire n_365;
wire n_91;
wire n_176;
wire n_182;
wire n_143;
wire n_83;
wire n_354;
wire n_237;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_66;
wire n_177;
wire n_359;
wire n_117;
wire n_326;
wire n_233;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_154;
wire n_62;
wire n_148;
wire n_71;
wire n_300;
wire n_159;
wire n_334;
wire n_391;
wire n_175;
wire n_262;
wire n_238;
wire n_99;
wire n_319;
wire n_364;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_64;
wire n_222;
wire n_89;
wire n_115;
wire n_324;
wire n_199;
wire n_187;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_6),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_44),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_38),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_8),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_4),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_60),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_30),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_46),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_31),
.B(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_61),
.B(n_97),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_2),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

AND3x2_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_12),
.C(n_17),
.Y(n_124)
);

OR2x6_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_113),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_18),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_23),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_32),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

CKINVDCx11_ASAP7_75t_R g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_64),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_34),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_103),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_37),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_96),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_43),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_59),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_66),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_132),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

OR2x6_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_78),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_92),
.Y(n_174)
);

NOR2x1p5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_92),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_95),
.B1(n_76),
.B2(n_80),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_95),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_158),
.Y(n_181)
);

AO22x2_ASAP7_75t_L g182 ( 
.A1(n_120),
.A2(n_121),
.B1(n_159),
.B2(n_132),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_121),
.B1(n_144),
.B2(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_162),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_154),
.Y(n_189)
);

OR2x6_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_157),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_166),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_155),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

OR2x6_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_164),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_122),
.B1(n_123),
.B2(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_119),
.B(n_155),
.Y(n_204)
);

NAND2x1p5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_164),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_167),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_161),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_165),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_191),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_144),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

AND2x4_ASAP7_75t_SL g226 ( 
.A(n_173),
.B(n_139),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

AND3x1_ASAP7_75t_SL g231 ( 
.A(n_175),
.B(n_148),
.C(n_140),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_177),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_177),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_124),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_136),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_133),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_137),
.B(n_116),
.C(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_168),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_171),
.B(n_145),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_190),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_232),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_171),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

HAxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_175),
.CON(n_265),
.SN(n_265)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_147),
.B1(n_160),
.B2(n_137),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_216),
.A2(n_147),
.B1(n_160),
.B2(n_171),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_255),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_222),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_201),
.B(n_203),
.C(n_204),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_182),
.B1(n_183),
.B2(n_168),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_234),
.A2(n_147),
.B1(n_160),
.B2(n_183),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

AND3x2_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_203),
.C(n_131),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_182),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_170),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_195),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_227),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_254),
.A2(n_205),
.B1(n_195),
.B2(n_190),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

OAI222xp33_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_199),
.B1(n_173),
.B2(n_131),
.C1(n_134),
.C2(n_151),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_237),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

OR2x6_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_135),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_217),
.B1(n_250),
.B2(n_247),
.Y(n_305)
);

CKINVDCx11_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_147),
.B1(n_160),
.B2(n_124),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_266),
.A2(n_147),
.B1(n_160),
.B2(n_230),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_261),
.A2(n_264),
.B1(n_268),
.B2(n_300),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

OR2x6_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_302),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_221),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_226),
.B(n_220),
.C(n_214),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_282),
.A2(n_229),
.B1(n_230),
.B2(n_134),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_211),
.B1(n_217),
.B2(n_244),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_300),
.A2(n_217),
.B1(n_141),
.B2(n_231),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_278),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_274),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_260),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_286),
.A2(n_248),
.B(n_249),
.C(n_238),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_246),
.B(n_238),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_301),
.A2(n_176),
.B1(n_187),
.B2(n_238),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_258),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_217),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_187),
.B1(n_192),
.B2(n_281),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_192),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_290),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_271),
.B1(n_302),
.B2(n_280),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

OAI221xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_297),
.B1(n_303),
.B2(n_291),
.C(n_279),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_315),
.A2(n_263),
.B(n_275),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_L g346 ( 
.A1(n_315),
.A2(n_271),
.B(n_294),
.C(n_277),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_302),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_267),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_331),
.A2(n_303),
.B1(n_269),
.B2(n_285),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_334),
.A2(n_303),
.B1(n_295),
.B2(n_287),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_326),
.A2(n_265),
.B1(n_262),
.B2(n_292),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_324),
.A2(n_262),
.B1(n_292),
.B2(n_265),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_295),
.B1(n_304),
.B2(n_288),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

OAI221xp5_ASAP7_75t_L g356 ( 
.A1(n_352),
.A2(n_309),
.B1(n_343),
.B2(n_337),
.C(n_350),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_333),
.C(n_284),
.Y(n_357)
);

AOI222xp33_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_299),
.B1(n_329),
.B2(n_325),
.C1(n_310),
.C2(n_307),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_346),
.A2(n_328),
.B(n_305),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_338),
.A2(n_311),
.B1(n_336),
.B2(n_299),
.Y(n_360)
);

OAI33xp33_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_335),
.A3(n_313),
.B1(n_330),
.B2(n_317),
.B3(n_327),
.Y(n_361)
);

AOI31xp67_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_332),
.A3(n_308),
.B(n_307),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_352),
.A2(n_311),
.B1(n_314),
.B2(n_312),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_349),
.A2(n_311),
.B1(n_314),
.B2(n_312),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_284),
.C(n_319),
.Y(n_366)
);

AOI221xp5_ASAP7_75t_SL g367 ( 
.A1(n_347),
.A2(n_316),
.B1(n_308),
.B2(n_304),
.C(n_288),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_316),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_340),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_355),
.Y(n_371)
);

OAI31xp33_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_366),
.A3(n_363),
.B(n_364),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_360),
.Y(n_373)
);

OAI322xp33_ASAP7_75t_SL g374 ( 
.A1(n_358),
.A2(n_341),
.A3(n_342),
.B1(n_344),
.B2(n_348),
.C1(n_351),
.C2(n_347),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_367),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_365),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_370),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_365),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_370),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_359),
.B(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_377),
.A2(n_374),
.B(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_380),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

XNOR2x2_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_378),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_382),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_387),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_390),
.A2(n_389),
.B(n_388),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_392),
.Y(n_393)
);

AND4x1_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_361),
.C(n_391),
.D(n_379),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_395),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_396),
.A2(n_379),
.B1(n_375),
.B2(n_348),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_397),
.B(n_375),
.Y(n_398)
);

AO21x2_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_304),
.B(n_362),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_399),
.A2(n_375),
.B(n_304),
.Y(n_400)
);


endmodule