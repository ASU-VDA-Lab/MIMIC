module real_aes_4831_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_L g28 ( .A(n_0), .B(n_6), .Y(n_28) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
AND2x4_ASAP7_75t_L g34 ( .A(n_1), .B(n_35), .Y(n_34) );
AND2x4_ASAP7_75t_L g43 ( .A(n_1), .B(n_4), .Y(n_43) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_2), .B(n_22), .Y(n_21) );
INVxp67_ASAP7_75t_L g38 ( .A(n_3), .Y(n_38) );
INVx1_ASAP7_75t_L g35 ( .A(n_4), .Y(n_35) );
BUFx6f_ASAP7_75t_L g25 ( .A(n_5), .Y(n_25) );
INVx2_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
INVx1_ASAP7_75t_SL g32 ( .A(n_8), .Y(n_32) );
AND2x4_ASAP7_75t_L g44 ( .A(n_8), .B(n_19), .Y(n_44) );
BUFx3_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_14), .B1(n_26), .B2(n_36), .C(n_39), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_13), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g15 ( .A(n_16), .B(n_18), .C(n_20), .Y(n_15) );
OAI21xp33_ASAP7_75t_L g26 ( .A1(n_16), .A2(n_27), .B(n_29), .Y(n_26) );
AOI211xp5_ASAP7_75t_L g29 ( .A1(n_16), .A2(n_21), .B(n_30), .C(n_34), .Y(n_29) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_17), .A2(n_32), .B(n_33), .Y(n_31) );
INVx1_ASAP7_75t_L g33 ( .A(n_18), .Y(n_33) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVxp67_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
INVx2_ASAP7_75t_SL g22 ( .A(n_23), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g40 ( .A(n_27), .B(n_37), .C(n_41), .Y(n_40) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
INVxp67_ASAP7_75t_SL g30 ( .A(n_31), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
BUFx2_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
AND2x4_ASAP7_75t_L g42 ( .A(n_43), .B(n_44), .Y(n_42) );
endmodule