module fake_jpeg_902_n_481 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_481);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_481;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_49),
.Y(n_130)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_55),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_62),
.B(n_32),
.Y(n_150)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_25),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_43),
.B(n_36),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_80),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_97),
.Y(n_116)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_10),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_23),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_94),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_0),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_27),
.B1(n_20),
.B2(n_35),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_103),
.A2(n_106),
.B1(n_156),
.B2(n_34),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_104),
.A2(n_153),
.B1(n_46),
.B2(n_38),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_27),
.B1(n_26),
.B2(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_28),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_127),
.B(n_154),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_46),
.B(n_1),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_78),
.A2(n_42),
.B1(n_35),
.B2(n_26),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_22),
.B1(n_45),
.B2(n_39),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_54),
.B(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_152),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_81),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_79),
.A2(n_43),
.B1(n_36),
.B2(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_32),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_90),
.A2(n_42),
.B1(n_35),
.B2(n_46),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_160),
.A2(n_205),
.B1(n_167),
.B2(n_143),
.Y(n_222)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_50),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_111),
.A2(n_103),
.B1(n_119),
.B2(n_105),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_169),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_56),
.B1(n_60),
.B2(n_53),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_165),
.A2(n_167),
.B1(n_176),
.B2(n_198),
.Y(n_227)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_106),
.A2(n_45),
.B1(n_22),
.B2(n_39),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_114),
.B(n_100),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_116),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_38),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_187),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_182),
.B(n_149),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_95),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_130),
.A2(n_42),
.B1(n_35),
.B2(n_98),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_196),
.B1(n_202),
.B2(n_203),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_115),
.A2(n_74),
.B(n_72),
.C(n_34),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_190),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_72),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_42),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_35),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_195),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_75),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_133),
.A2(n_73),
.B1(n_65),
.B2(n_61),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_132),
.A2(n_74),
.B1(n_58),
.B2(n_52),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_124),
.A2(n_48),
.B1(n_34),
.B2(n_40),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_129),
.B1(n_122),
.B2(n_158),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_34),
.B1(n_40),
.B2(n_2),
.Y(n_205)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_149),
.A3(n_139),
.B1(n_138),
.B2(n_109),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_203),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_146),
.B1(n_140),
.B2(n_143),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_229),
.B1(n_164),
.B2(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_134),
.C(n_125),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_186),
.C(n_163),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_200),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_203),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_158),
.B1(n_102),
.B2(n_123),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_228),
.A2(n_235),
.B1(n_192),
.B2(n_177),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_148),
.B1(n_141),
.B2(n_145),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_238),
.B1(n_186),
.B2(n_192),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_165),
.B1(n_145),
.B2(n_123),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_163),
.A2(n_129),
.B1(n_108),
.B2(n_121),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_226),
.B(n_211),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_260),
.B(n_224),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_262),
.B1(n_266),
.B2(n_222),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_237),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_255),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_206),
.B(n_214),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_188),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_239),
.C(n_237),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_250),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_188),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_164),
.B1(n_182),
.B2(n_168),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_254),
.B1(n_211),
.B2(n_213),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_203),
.B1(n_193),
.B2(n_169),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_174),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_261),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_206),
.A2(n_220),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_221),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_169),
.B(n_185),
.C(n_195),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_212),
.B(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_209),
.B(n_172),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_267),
.Y(n_294)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_227),
.A2(n_169),
.B1(n_141),
.B2(n_148),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_201),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_269),
.A2(n_272),
.B1(n_274),
.B2(n_290),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_235),
.B1(n_234),
.B2(n_213),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_254),
.A2(n_228),
.B1(n_210),
.B2(n_223),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_210),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_279),
.A2(n_281),
.B1(n_292),
.B2(n_250),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_239),
.B1(n_217),
.B2(n_208),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.C(n_242),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_237),
.C(n_236),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_236),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_249),
.A2(n_238),
.B1(n_231),
.B2(n_218),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_259),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_229),
.B1(n_217),
.B2(n_232),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_252),
.A2(n_169),
.B1(n_233),
.B2(n_232),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_256),
.B1(n_263),
.B2(n_262),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_257),
.B(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_251),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_317),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_260),
.B1(n_241),
.B2(n_240),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_297),
.A2(n_306),
.B1(n_313),
.B2(n_320),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_303),
.C(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_279),
.B1(n_260),
.B2(n_243),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_300),
.A2(n_319),
.B1(n_273),
.B2(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_243),
.C(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_241),
.B1(n_240),
.B2(n_246),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_243),
.C(n_248),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

OAI21x1_ASAP7_75t_R g328 ( 
.A1(n_311),
.A2(n_322),
.B(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_264),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_321),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_316),
.Y(n_333)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_323),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_290),
.A2(n_259),
.B1(n_265),
.B2(n_258),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_255),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_224),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_278),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_339),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_326),
.A2(n_331),
.B1(n_302),
.B2(n_299),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_305),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_269),
.B1(n_272),
.B2(n_287),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_332),
.B(n_343),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_SL g334 ( 
.A(n_297),
.B(n_287),
.C(n_284),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_334),
.B(n_337),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_314),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_294),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_285),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_348),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_301),
.B(n_268),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_346),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_268),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_270),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_300),
.B(n_244),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_349),
.B(n_301),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_304),
.A2(n_291),
.B1(n_277),
.B2(n_280),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_350),
.A2(n_318),
.B1(n_313),
.B2(n_317),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_245),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_324),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_352),
.B(n_358),
.Y(n_382)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_356),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_357),
.A2(n_364),
.B1(n_375),
.B2(n_280),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_324),
.B(n_316),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_328),
.B(n_312),
.CI(n_310),
.CON(n_360),
.SN(n_360)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_361),
.Y(n_397)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_365),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_225),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_376),
.B(n_377),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_277),
.C(n_207),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_338),
.C(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_289),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_351),
.B1(n_326),
.B2(n_350),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_161),
.B(n_199),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_190),
.B(n_194),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_387),
.C(n_388),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_325),
.C(n_339),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_375),
.A2(n_331),
.B1(n_342),
.B2(n_330),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_368),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_393),
.Y(n_404)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_349),
.C(n_348),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_346),
.C(n_225),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_353),
.B(n_215),
.Y(n_389)
);

OAI221xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_374),
.B1(n_362),
.B2(n_365),
.C(n_361),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_346),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_377),
.C(n_359),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_372),
.C(n_376),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_399),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_216),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g400 ( 
.A(n_382),
.B(n_367),
.CI(n_360),
.CON(n_400),
.SN(n_400)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_216),
.Y(n_428)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_SL g431 ( 
.A(n_403),
.B(n_409),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_382),
.B(n_370),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_196),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_392),
.A2(n_357),
.B1(n_356),
.B2(n_360),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_411),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_280),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_384),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_379),
.Y(n_413)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_413),
.Y(n_435)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_415),
.Y(n_434)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_253),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_418),
.Y(n_429)
);

OAI221xp5_ASAP7_75t_L g417 ( 
.A1(n_395),
.A2(n_391),
.B1(n_390),
.B2(n_380),
.C(n_398),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_417),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_388),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_408),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_419),
.B(n_170),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_383),
.B1(n_399),
.B2(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_401),
.C(n_409),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_425),
.Y(n_437)
);

BUFx6f_ASAP7_75t_SL g425 ( 
.A(n_410),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_403),
.A2(n_383),
.B1(n_253),
.B2(n_162),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_432),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_427),
.B(n_184),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_400),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_406),
.A2(n_204),
.B1(n_215),
.B2(n_177),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_166),
.C(n_173),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_404),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_439),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_420),
.B(n_418),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_440),
.B(n_433),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_SL g441 ( 
.A1(n_422),
.A2(n_400),
.B(n_405),
.C(n_404),
.Y(n_441)
);

AOI21xp33_ASAP7_75t_L g458 ( 
.A1(n_441),
.A2(n_427),
.B(n_425),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_443),
.B(n_445),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_449),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_121),
.C(n_112),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_191),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_446),
.B(n_448),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_431),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_429),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_424),
.B(n_112),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_108),
.B1(n_34),
.B2(n_40),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_451),
.A2(n_453),
.B(n_0),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_456),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_447),
.A2(n_428),
.B1(n_435),
.B2(n_421),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_455),
.B(n_450),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_0),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_460),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_441),
.B(n_438),
.Y(n_460)
);

A2O1A1O1Ixp25_ASAP7_75t_L g461 ( 
.A1(n_454),
.A2(n_436),
.B(n_444),
.C(n_2),
.D(n_4),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_461),
.A2(n_467),
.B(n_462),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_0),
.C(n_1),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_1),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_8),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_1),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_470),
.B(n_471),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_468),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_4),
.B(n_6),
.Y(n_476)
);

AOI322xp5_ASAP7_75t_L g473 ( 
.A1(n_462),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_469),
.C(n_5),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_7),
.C(n_8),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_6),
.B(n_7),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g479 ( 
.A(n_477),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_475),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_478),
.B(n_8),
.Y(n_481)
);


endmodule