module fake_jpeg_31767_n_494 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_49),
.Y(n_148)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_50),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_23),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_48),
.B1(n_47),
.B2(n_30),
.Y(n_117)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_25),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_92),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_40),
.B1(n_48),
.B2(n_47),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_1),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_91),
.Y(n_106)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_96),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_23),
.B1(n_39),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_99),
.A2(n_107),
.B1(n_108),
.B2(n_124),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_102),
.B(n_118),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_40),
.B1(n_32),
.B2(n_23),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_117),
.A2(n_8),
.B(n_10),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_38),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_23),
.B1(n_39),
.B2(n_42),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_132),
.B1(n_139),
.B2(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_140),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_75),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_34),
.B1(n_43),
.B2(n_36),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_150),
.B1(n_96),
.B2(n_94),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_52),
.A2(n_35),
.B1(n_30),
.B2(n_18),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_95),
.B(n_33),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_54),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_153),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_69),
.A2(n_46),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_4),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_76),
.B1(n_72),
.B2(n_56),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_157),
.A2(n_167),
.B1(n_208),
.B2(n_111),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_108),
.A2(n_61),
.B1(n_63),
.B2(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_158),
.A2(n_177),
.B1(n_193),
.B2(n_203),
.Y(n_216)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_163),
.B(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_84),
.B1(n_71),
.B2(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_101),
.B(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_169),
.B(n_174),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_97),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_175),
.B(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_65),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_106),
.B(n_5),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_212),
.Y(n_221)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_49),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_51),
.C(n_88),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_199),
.C(n_210),
.Y(n_220)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_192),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_100),
.A2(n_46),
.B1(n_7),
.B2(n_8),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_46),
.C(n_7),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_131),
.B(n_46),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_98),
.B(n_6),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_209),
.B(n_211),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_100),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_205),
.Y(n_235)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_145),
.A2(n_141),
.B1(n_133),
.B2(n_152),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_116),
.B1(n_141),
.B2(n_152),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_110),
.B(n_10),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_117),
.B(n_10),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_116),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_219),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_128),
.C(n_154),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_161),
.C(n_200),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_170),
.B1(n_166),
.B2(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_257),
.B1(n_258),
.B2(n_167),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_248),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_145),
.B1(n_121),
.B2(n_156),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_212),
.B1(n_187),
.B2(n_183),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_210),
.A2(n_104),
.B1(n_154),
.B2(n_156),
.Y(n_248)
);

MAJx3_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_104),
.C(n_11),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_252),
.A2(n_220),
.B(n_219),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_122),
.B1(n_119),
.B2(n_104),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_177),
.A2(n_109),
.B1(n_105),
.B2(n_12),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_10),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_13),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_267),
.B1(n_282),
.B2(n_254),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_173),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_265),
.B(n_271),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_161),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_304),
.C(n_260),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_296),
.B1(n_254),
.B2(n_244),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_273),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_206),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

AOI32xp33_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_161),
.A3(n_192),
.B1(n_204),
.B2(n_194),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_191),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_280),
.Y(n_334)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_215),
.A2(n_161),
.B1(n_196),
.B2(n_180),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_242),
.B1(n_232),
.B2(n_244),
.Y(n_312)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_234),
.A2(n_213),
.B1(n_205),
.B2(n_181),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_179),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_216),
.A2(n_201),
.B1(n_198),
.B2(n_196),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_109),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_283),
.B(n_295),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_222),
.B(n_186),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_289),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_252),
.A2(n_159),
.B(n_105),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_285),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_286)
);

NAND2x1p5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_248),
.A2(n_13),
.B(n_15),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_288),
.A2(n_246),
.B(n_230),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_222),
.B(n_13),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_221),
.B(n_219),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_290),
.B(n_292),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_261),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_217),
.B(n_15),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_221),
.B(n_16),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_243),
.A2(n_16),
.B1(n_17),
.B2(n_233),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_229),
.Y(n_299)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_220),
.B(n_16),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_301),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_237),
.B(n_17),
.Y(n_301)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_226),
.B(n_236),
.C(n_261),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_235),
.B(n_226),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_256),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_253),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_235),
.B1(n_242),
.B2(n_225),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_309),
.A2(n_315),
.B(n_323),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_317),
.B1(n_269),
.B2(n_305),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_312),
.A2(n_314),
.B1(n_332),
.B2(n_340),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_263),
.A2(n_254),
.B1(n_228),
.B2(n_249),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_283),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_331),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_280),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_328),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_266),
.A2(n_246),
.B(n_253),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_275),
.A2(n_250),
.B1(n_260),
.B2(n_247),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_250),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_338),
.C(n_343),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_275),
.A2(n_218),
.B1(n_224),
.B2(n_247),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_266),
.A2(n_218),
.B(n_224),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_342),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_268),
.B(n_290),
.C(n_281),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_302),
.A2(n_296),
.B1(n_266),
.B2(n_264),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_344),
.A2(n_281),
.B1(n_278),
.B2(n_285),
.Y(n_355)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_302),
.B1(n_264),
.B2(n_273),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_355),
.B1(n_364),
.B2(n_365),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_351),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_349),
.A2(n_350),
.B1(n_363),
.B2(n_366),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_305),
.B1(n_288),
.B2(n_281),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_320),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_352),
.B(n_360),
.Y(n_386)
);

OAI32xp33_ASAP7_75t_L g353 ( 
.A1(n_308),
.A2(n_285),
.A3(n_270),
.B1(n_265),
.B2(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_339),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_300),
.C(n_283),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_362),
.C(n_369),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_271),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_358),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_274),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_283),
.C(n_304),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_308),
.A2(n_305),
.B1(n_301),
.B2(n_293),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_307),
.A2(n_272),
.B1(n_277),
.B2(n_298),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_307),
.A2(n_287),
.B1(n_292),
.B2(n_306),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_311),
.A2(n_284),
.B1(n_294),
.B2(n_289),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_367),
.Y(n_399)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_286),
.C(n_299),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_324),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_286),
.C(n_299),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_376),
.C(n_323),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_319),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_334),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_303),
.C(n_325),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_380),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_384),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_348),
.B(n_337),
.Y(n_382)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_359),
.B(n_331),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_387),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_339),
.C(n_325),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_392),
.C(n_395),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_309),
.B(n_321),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_371),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_341),
.C(n_342),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_327),
.B1(n_314),
.B2(n_310),
.Y(n_393)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_393),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_341),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_357),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_374),
.A2(n_315),
.B(n_376),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_401),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_326),
.B(n_337),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_402),
.A2(n_366),
.B1(n_326),
.B2(n_327),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_315),
.B1(n_324),
.B2(n_330),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_375),
.B1(n_345),
.B2(n_364),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_409),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_369),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_416),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_355),
.C(n_363),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.C(n_421),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_392),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_417),
.A2(n_418),
.B1(n_381),
.B2(n_382),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_385),
.A2(n_345),
.B1(n_365),
.B2(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_419),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_384),
.C(n_379),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_350),
.C(n_349),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_387),
.B(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_426),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_370),
.C(n_368),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_380),
.C(n_378),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_396),
.B1(n_385),
.B2(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_435),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_443),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_436),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_407),
.B1(n_418),
.B2(n_423),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_404),
.B1(n_390),
.B2(n_381),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_403),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_403),
.C(n_400),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_445),
.C(n_427),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_422),
.B(n_400),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_442),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_389),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_421),
.B(n_389),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_412),
.A2(n_361),
.B1(n_346),
.B2(n_399),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_417),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_399),
.C(n_330),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_438),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_440),
.B(n_424),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_448),
.B(n_456),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_413),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_445),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_451),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_454),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_428),
.A2(n_413),
.B(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_455),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_438),
.C(n_437),
.Y(n_456)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_460),
.A2(n_435),
.B1(n_429),
.B2(n_443),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_467),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_450),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_464),
.A2(n_465),
.B1(n_449),
.B2(n_333),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_457),
.A2(n_329),
.B1(n_333),
.B2(n_336),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_450),
.B(n_439),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_469),
.B(n_471),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_428),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_466),
.A2(n_447),
.B(n_452),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_472),
.B(n_477),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_478),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_410),
.C(n_436),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_458),
.B(n_429),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_467),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_468),
.C(n_410),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_483),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_461),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_474),
.Y(n_487)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g488 ( 
.A1(n_486),
.A2(n_484),
.B(n_477),
.C(n_415),
.D(n_481),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_478),
.C(n_453),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_489),
.B(n_453),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_465),
.B(n_336),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_492),
.A2(n_303),
.B(n_409),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_493),
.Y(n_494)
);


endmodule