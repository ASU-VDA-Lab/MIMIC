module fake_jpeg_2358_n_557 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_557);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_54),
.B(n_83),
.Y(n_161)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_99),
.Y(n_130)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_33),
.B1(n_49),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_23),
.B1(n_46),
.B2(n_39),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_33),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_11),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_53),
.CON(n_134),
.SN(n_134)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_102),
.B(n_23),
.Y(n_163)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_104),
.Y(n_148)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_53),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_107),
.B1(n_31),
.B2(n_41),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_48),
.B1(n_43),
.B2(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_108),
.A2(n_114),
.B1(n_121),
.B2(n_122),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_26),
.B1(n_50),
.B2(n_42),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_112),
.A2(n_115),
.B1(n_159),
.B2(n_165),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_48),
.B1(n_43),
.B2(n_24),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_86),
.B1(n_90),
.B2(n_68),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_54),
.A2(n_26),
.B1(n_50),
.B2(n_42),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_118),
.A2(n_114),
.B(n_122),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_48),
.B1(n_43),
.B2(n_24),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_134),
.A2(n_17),
.B(n_16),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_147),
.B1(n_154),
.B2(n_164),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_27),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_143),
.B(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_56),
.A2(n_38),
.B1(n_30),
.B2(n_20),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_94),
.A2(n_38),
.B1(n_46),
.B2(n_39),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_59),
.B(n_46),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_39),
.B1(n_23),
.B2(n_41),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_58),
.A2(n_41),
.B1(n_31),
.B2(n_36),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_93),
.A2(n_41),
.B1(n_31),
.B2(n_2),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_41),
.B1(n_31),
.B2(n_36),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_166),
.A2(n_172),
.B1(n_44),
.B2(n_18),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_79),
.B(n_14),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_0),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_91),
.A2(n_41),
.B1(n_31),
.B2(n_2),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_176),
.Y(n_250)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_177),
.Y(n_275)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_132),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_179),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_180),
.Y(n_285)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_130),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_185),
.B(n_194),
.Y(n_274)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_191),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_119),
.B(n_107),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_196),
.B(n_197),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_137),
.Y(n_199)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_115),
.A2(n_106),
.B1(n_103),
.B2(n_97),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_154),
.B1(n_165),
.B2(n_172),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_218),
.Y(n_253)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_207),
.Y(n_292)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_212),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_13),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_213),
.Y(n_265)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_219),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_13),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_217),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_111),
.B(n_150),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_133),
.A2(n_95),
.B1(n_31),
.B2(n_36),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_220),
.A2(n_15),
.B1(n_17),
.B2(n_179),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_110),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_223),
.Y(n_283)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_141),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_222),
.Y(n_293)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_225),
.Y(n_296)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_109),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_226),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_12),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_231),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_228),
.Y(n_284)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_126),
.B(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_12),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_110),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_237),
.B1(n_44),
.B2(n_18),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_290),
.B1(n_215),
.B2(n_182),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_166),
.C(n_108),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_243),
.B(n_257),
.C(n_269),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_113),
.B1(n_159),
.B2(n_152),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_251),
.B1(n_272),
.B2(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_113),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_260),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_249),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_155),
.B1(n_152),
.B2(n_139),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_44),
.B1(n_37),
.B2(n_13),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_256),
.A2(n_289),
.B1(n_294),
.B2(n_248),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_155),
.C(n_139),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_0),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_222),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_5),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_190),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_276),
.A2(n_297),
.B1(n_290),
.B2(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_190),
.B(n_4),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_186),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_208),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_241),
.B(n_282),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_208),
.A2(n_6),
.B1(n_15),
.B2(n_17),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_207),
.A2(n_15),
.B1(n_17),
.B2(n_209),
.Y(n_289)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_220),
.A2(n_193),
.B1(n_181),
.B2(n_223),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_299),
.A2(n_312),
.B1(n_314),
.B2(n_318),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_245),
.B(n_219),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_300),
.B(n_311),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_334),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_303),
.A2(n_327),
.B1(n_338),
.B2(n_339),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_210),
.B(n_192),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_304),
.A2(n_333),
.B(n_347),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_243),
.A2(n_184),
.B(n_189),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_307),
.A2(n_325),
.B(n_285),
.Y(n_363)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_175),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_277),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_245),
.B(n_230),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_269),
.B1(n_242),
.B2(n_279),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_313),
.B(n_320),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_235),
.B1(n_226),
.B2(n_183),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_275),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_315),
.B(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_180),
.B1(n_188),
.B2(n_246),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_341),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_321),
.B(n_331),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_263),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_322),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_323),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_247),
.A2(n_251),
.B1(n_254),
.B2(n_280),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_324),
.A2(n_329),
.B1(n_335),
.B2(n_287),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_262),
.A2(n_283),
.B(n_294),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_257),
.B(n_265),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_262),
.A2(n_258),
.B1(n_293),
.B2(n_275),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_262),
.A2(n_250),
.B1(n_271),
.B2(n_292),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_284),
.A2(n_240),
.B(n_270),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_255),
.B(n_268),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_292),
.A2(n_281),
.B1(n_259),
.B2(n_291),
.Y(n_335)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_252),
.B(n_281),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_344),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_255),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_322),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g345 ( 
.A(n_248),
.B(n_244),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_345),
.A2(n_295),
.B(n_267),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_346),
.Y(n_385)
);

AOI22x1_ASAP7_75t_SL g347 ( 
.A1(n_252),
.A2(n_295),
.B1(n_273),
.B2(n_266),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_300),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_351),
.Y(n_393)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_355),
.B(n_381),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_358),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_363),
.A2(n_364),
.B(n_381),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_304),
.A2(n_325),
.B(n_310),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_286),
.B1(n_266),
.B2(n_285),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_365),
.A2(n_380),
.B1(n_336),
.B2(n_317),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_377),
.B1(n_382),
.B2(n_343),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_287),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_386),
.C(n_341),
.Y(n_410)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_303),
.A2(n_333),
.B(n_329),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_384),
.B(n_341),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_312),
.A2(n_299),
.B1(n_319),
.B2(n_307),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_301),
.B(n_311),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_356),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_305),
.A2(n_302),
.B1(n_316),
.B2(n_340),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_303),
.A2(n_301),
.B(n_306),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_324),
.A2(n_318),
.B1(n_330),
.B2(n_314),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_327),
.A2(n_345),
.B(n_330),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_374),
.B(n_345),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_392),
.B(n_408),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_394),
.A2(n_400),
.B1(n_409),
.B2(n_415),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_388),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_396),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_388),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_399),
.A2(n_359),
.B(n_378),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_308),
.B1(n_309),
.B2(n_347),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_401),
.B(n_411),
.Y(n_433)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_342),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_375),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_377),
.A2(n_298),
.B1(n_337),
.B2(n_336),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_423),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_386),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_371),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_412),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_335),
.C(n_328),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_421),
.C(n_360),
.Y(n_448)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_417),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_419),
.B(n_366),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_358),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_420),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_384),
.C(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_367),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_422),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_367),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_389),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_424),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_352),
.B(n_378),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_352),
.Y(n_429)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_351),
.B1(n_383),
.B2(n_372),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_435),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_412),
.A2(n_383),
.B1(n_353),
.B2(n_363),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_397),
.A2(n_361),
.B1(n_383),
.B2(n_368),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_402),
.B1(n_422),
.B2(n_391),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_438),
.A2(n_392),
.B(n_408),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_359),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_440),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_361),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_397),
.A2(n_387),
.B1(n_373),
.B2(n_390),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_447),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_400),
.A2(n_373),
.B1(n_360),
.B2(n_376),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_441),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_354),
.C(n_357),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_452),
.C(n_398),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_354),
.C(n_357),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_399),
.A2(n_376),
.B(n_366),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_453),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_455),
.B(n_423),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_409),
.A2(n_420),
.B1(n_402),
.B2(n_416),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_456),
.A2(n_395),
.B(n_407),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_458),
.B(n_479),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_393),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_464),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_445),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_467),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_465),
.C(n_466),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_393),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_398),
.C(n_396),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_426),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_407),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_470),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_481),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_472),
.A2(n_475),
.B1(n_480),
.B2(n_437),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_425),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_449),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_436),
.A2(n_424),
.B1(n_391),
.B2(n_405),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_403),
.C(n_406),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_478),
.C(n_428),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_414),
.C(n_418),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_415),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_427),
.A2(n_431),
.B1(n_430),
.B2(n_446),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_438),
.A2(n_430),
.B(n_456),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_471),
.A2(n_446),
.B(n_433),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_483),
.B(n_487),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_474),
.A2(n_431),
.B1(n_427),
.B2(n_432),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_484),
.A2(n_472),
.B1(n_481),
.B2(n_479),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_453),
.C(n_435),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_497),
.C(n_499),
.Y(n_505)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

OAI221xp5_ASAP7_75t_L g506 ( 
.A1(n_496),
.A2(n_473),
.B1(n_464),
.B2(n_482),
.C(n_461),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_466),
.C(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_469),
.Y(n_498)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_434),
.C(n_428),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_442),
.C(n_447),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_501),
.C(n_490),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_443),
.C(n_437),
.Y(n_501)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_469),
.Y(n_504)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_506),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_495),
.B(n_468),
.Y(n_507)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_513),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_508),
.A2(n_511),
.B1(n_486),
.B2(n_520),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_485),
.A2(n_459),
.B1(n_444),
.B2(n_451),
.Y(n_509)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_484),
.A2(n_475),
.B1(n_443),
.B2(n_451),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_493),
.A2(n_444),
.B(n_458),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_492),
.B(n_501),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_502),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_503),
.A2(n_488),
.B1(n_492),
.B2(n_500),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_508),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_519),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_490),
.B(n_489),
.Y(n_519)
);

O2A1O1Ixp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_499),
.B(n_517),
.C(n_497),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_524),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_527),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_486),
.C(n_505),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_533),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_511),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_529),
.A2(n_507),
.B1(n_530),
.B2(n_531),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_512),
.A2(n_515),
.B(n_514),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_514),
.B(n_510),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_519),
.C(n_513),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_536),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_527),
.B(n_510),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_537),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_529),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_540),
.B(n_542),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_524),
.A2(n_528),
.B(n_532),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_525),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_533),
.B(n_523),
.Y(n_542)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_543),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_535),
.C(n_523),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_544),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_SL g549 ( 
.A(n_546),
.B(n_534),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_549),
.A2(n_538),
.B(n_545),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_552),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_550),
.C(n_538),
.Y(n_554)
);

BUFx24_ASAP7_75t_SL g555 ( 
.A(n_554),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_541),
.C(n_526),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_526),
.Y(n_557)
);


endmodule