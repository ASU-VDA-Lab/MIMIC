module fake_jpeg_16206_n_78 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_14),
.B1(n_26),
.B2(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_1),
.B(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_59),
.B(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_3),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_41),
.B(n_43),
.C(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_31),
.B1(n_15),
.B2(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_8),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_31),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_57),
.C(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_5),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B(n_62),
.Y(n_72)
);

OAI221xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_66),
.B1(n_69),
.B2(n_63),
.C(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_9),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.C(n_27),
.Y(n_78)
);


endmodule