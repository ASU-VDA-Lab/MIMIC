module real_jpeg_31337_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_0),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_0),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_2),
.Y(n_108)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_67),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_3),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_3),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_13),
.B1(n_64),
.B2(n_68),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_48),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_8),
.B(n_68),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_8),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_10),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2x1_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_84),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_10),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_84),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_10),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_12),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_13),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_13),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_13),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_13),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_13),
.B(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_14),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_14),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_15),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_15),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_15),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_15),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_15),
.B(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_214),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_R g17 ( 
.A(n_18),
.B(n_211),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_159),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_19),
.B(n_159),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.C(n_140),
.Y(n_19)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_20),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_21),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_52),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_23),
.B(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_25),
.B(n_33),
.C(n_34),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_31),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_31),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_37),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_38),
.B(n_52),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.C(n_47),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_39),
.A2(n_47),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_42),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_43),
.B(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_45),
.Y(n_329)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_51),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_53),
.B(n_58),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_57),
.B(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_57),
.B(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_58),
.B(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_59),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_82),
.Y(n_60)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_71),
.B2(n_81),
.Y(n_61)
);

OA21x2_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_130),
.B(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_63),
.B(n_180),
.C(n_181),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_67),
.Y(n_342)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_77),
.Y(n_327)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_78),
.Y(n_180)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_162),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_97),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_86),
.Y(n_291)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_95),
.C(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_95),
.A2(n_96),
.B1(n_102),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_98),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_115),
.C(n_129),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_99),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_109),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_100),
.A2(n_101),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_102),
.Y(n_277)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_103),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_262)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_107),
.B(n_285),
.Y(n_349)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_114),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_115),
.B(n_129),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_121),
.C(n_127),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_121),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_140),
.B(n_247),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_143),
.C(n_158),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_153),
.C(n_157),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_157),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_183),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_182),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_179),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_194),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_193),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_189),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_189),
.B(n_266),
.Y(n_303)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_191),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_194)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_204),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_202),
.Y(n_357)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_208),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_249),
.B(n_370),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_245),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_218),
.B(n_245),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_243),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_241),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_241),
.B1(n_242),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.C(n_236),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_227),
.A2(n_228),
.B1(n_236),
.B2(n_237),
.Y(n_311)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_278),
.B(n_369),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_253),
.B(n_255),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.C(n_263),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_257),
.B(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_260),
.B(n_263),
.Y(n_367)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.C(n_275),
.Y(n_263)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_268),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_270),
.A2(n_275),
.B1(n_276),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_363),
.B(n_368),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_318),
.B(n_362),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_304),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_281),
.B(n_304),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_295),
.C(n_303),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_282),
.B(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_292),
.C(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_297),
.A2(n_300),
.B1(n_301),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_312),
.B1(n_316),
.B2(n_317),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_317),
.C(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_333),
.B(n_361),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_330),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_330),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.C(n_328),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_321),
.A2(n_322),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_347),
.B(n_360),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_338),
.Y(n_360)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_339),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_354),
.B(n_359),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_358),
.Y(n_359)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_366),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);


endmodule