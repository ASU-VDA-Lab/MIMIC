module real_jpeg_24186_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_0),
.B(n_2),
.Y(n_160)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_2),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_2),
.B(n_25),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_5),
.B(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_75),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_56),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_33),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_29),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_5),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_5),
.B(n_256),
.Y(n_345)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_8),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_8),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_8),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_29),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_8),
.B(n_25),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_8),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_9),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_9),
.B(n_56),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_9),
.B(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_29),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_9),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_9),
.B(n_38),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_10),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_171),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_10),
.B(n_75),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_10),
.B(n_56),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_10),
.B(n_33),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_12),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_12),
.B(n_33),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_115),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_12),
.B(n_75),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_12),
.B(n_56),
.Y(n_337)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_36),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_14),
.B(n_115),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_14),
.B(n_75),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_14),
.B(n_33),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_14),
.B(n_29),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_56),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_25),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_17),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_17),
.B(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_17),
.B(n_75),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_17),
.B(n_29),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_17),
.B(n_25),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_58),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.C(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_52),
.C(n_54),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_49),
.B1(n_54),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_39),
.B(n_156),
.Y(n_215)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_43),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_43),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_44),
.B(n_150),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_44),
.B(n_251),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_53),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_72),
.C(n_74),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_54),
.A2(n_74),
.B1(n_79),
.B2(n_332),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_55),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_55),
.B(n_73),
.Y(n_264)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_81),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_59),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.C(n_77),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_60),
.B(n_376),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_61),
.B(n_81),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.CI(n_64),
.CON(n_61),
.SN(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.C(n_69),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_65),
.B(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_71),
.B(n_77),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_72),
.B(n_357),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_74),
.A2(n_303),
.B1(n_304),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_74),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_74),
.B(n_303),
.C(n_330),
.Y(n_361)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_380),
.C(n_381),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_371),
.C(n_372),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_349),
.C(n_350),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_325),
.C(n_326),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_293),
.C(n_294),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_258),
.C(n_259),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_221),
.C(n_222),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_191),
.C(n_192),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_165),
.C(n_166),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_126),
.C(n_137),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_107),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_102),
.C(n_107),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_97),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_105),
.C(n_106),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_108),
.B(n_118),
.C(n_119),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_111),
.Y(n_254)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_115),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_125),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_136),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_161),
.C(n_162),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_146),
.C(n_153),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_144),
.C(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.C(n_158),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_180),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_181),
.C(n_190),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_175),
.C(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_174),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_176),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.CI(n_179),
.CON(n_176),
.SN(n_176)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_207),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_196),
.C(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_203),
.C(n_206),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_198),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.CI(n_201),
.CON(n_198),
.SN(n_198)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_200),
.C(n_201),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_214),
.C(n_219),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_246),
.C(n_247),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_242),
.B2(n_257),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_243),
.C(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_227),
.C(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_235),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_231),
.C(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_239),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_252),
.C(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_291),
.B2(n_292),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_282),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_282),
.C(n_291),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_271),
.C(n_272),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_275),
.B1(n_276),
.B2(n_281),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_278),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_300),
.C(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_297),
.C(n_324),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_311),
.B2(n_324),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_306),
.C(n_307),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_307),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.CI(n_310),
.CON(n_307),
.SN(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_323),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_319),
.C(n_321),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_320),
.A2(n_321),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_346),
.C(n_347),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_348),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_339),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_339),
.C(n_348),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_334),
.C(n_335),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_335),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.CI(n_338),
.CON(n_335),
.SN(n_335)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_337),
.C(n_338),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.C(n_343),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_353),
.C(n_363),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_362),
.B2(n_363),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_360),
.C(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_366),
.C(n_369),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_372)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_375),
.C(n_379),
.Y(n_380)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);


endmodule