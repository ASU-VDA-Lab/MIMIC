module fake_jpeg_4743_n_157 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_157);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_22),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_20),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_47),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_51),
.Y(n_68)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_22),
.B1(n_31),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_61),
.B1(n_34),
.B2(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_35),
.B1(n_16),
.B2(n_17),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_53),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_25),
.B1(n_19),
.B2(n_42),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_42),
.B1(n_43),
.B2(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_97),
.B1(n_32),
.B2(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_60),
.C(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_43),
.C(n_57),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_74),
.B(n_72),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_80),
.B(n_86),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_110),
.B1(n_84),
.B2(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_93),
.B1(n_94),
.B2(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_117),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_25),
.B(n_19),
.C(n_57),
.D(n_38),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_27),
.B(n_23),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_101),
.B(n_99),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_102),
.C(n_55),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_106),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_131),
.C(n_113),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_115),
.C(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.C(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_122),
.B1(n_114),
.B2(n_119),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_102),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_32),
.A3(n_23),
.B1(n_28),
.B2(n_27),
.C(n_24),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_130),
.B(n_71),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_133),
.C(n_69),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_28),
.C(n_49),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_148),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_142),
.B1(n_49),
.B2(n_14),
.Y(n_149)
);

OAI321xp33_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_3),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_11),
.B(n_4),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_9),
.Y(n_157)
);


endmodule