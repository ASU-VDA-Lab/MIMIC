module fake_jpeg_17542_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_25),
.B1(n_18),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_45),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_25),
.B(n_13),
.C(n_22),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_48),
.B(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_25),
.B1(n_18),
.B2(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_18),
.B1(n_13),
.B2(n_23),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_17),
.B1(n_15),
.B2(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_62),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_34),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_15),
.B1(n_28),
.B2(n_24),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_40),
.C(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_78),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_70),
.B(n_65),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_28),
.B(n_33),
.C(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_58),
.C(n_57),
.Y(n_86)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_88),
.B(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_77),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_66),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_95),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_93),
.B(n_70),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_81),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_24),
.B1(n_20),
.B2(n_10),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_4),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_83),
.B1(n_91),
.B2(n_79),
.Y(n_111)
);

OAI322xp33_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_103),
.A3(n_108),
.B1(n_96),
.B2(n_93),
.C1(n_90),
.C2(n_83),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_86),
.C(n_43),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_71),
.A3(n_68),
.B1(n_80),
.B2(n_76),
.C1(n_34),
.C2(n_43),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_78),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_68),
.B(n_24),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_55),
.B(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_67),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_9),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_100),
.C(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_118),
.B1(n_99),
.B2(n_24),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.C(n_118),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_124),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_116),
.C(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_130),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_112),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_131),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_117),
.B(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_42),
.C(n_46),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_42),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_137),
.C(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_42),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_132),
.C(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_6),
.C(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_8),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_139),
.Y(n_143)
);


endmodule