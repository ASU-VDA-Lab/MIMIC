module real_aes_18314_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_456;
wire n_156;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_0), .A2(n_452), .B(n_456), .C(n_461), .Y(n_451) );
INVx1_ASAP7_75t_L g509 ( .A(n_0), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_1), .A2(n_30), .B1(n_105), .B2(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g481 ( .A(n_2), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_2), .B(n_447), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_3), .A2(n_9), .B1(n_145), .B2(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g540 ( .A(n_4), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_5), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_6), .A2(n_10), .B1(n_89), .B2(n_147), .Y(n_200) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_7), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_8), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_11), .A2(n_38), .B1(n_436), .B2(n_444), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_11), .A2(n_14), .B1(n_516), .B2(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g492 ( .A(n_12), .Y(n_492) );
INVx1_ASAP7_75t_L g502 ( .A(n_12), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_13), .A2(n_76), .B1(n_145), .B2(n_164), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_14), .A2(n_59), .B1(n_472), .B2(n_475), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_15), .A2(n_27), .B1(n_178), .B2(n_179), .Y(n_177) );
INVx2_ASAP7_75t_L g494 ( .A(n_16), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_17), .B(n_146), .Y(n_216) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_18), .A2(n_41), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g466 ( .A(n_19), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_20), .Y(n_171) );
INVx1_ASAP7_75t_L g548 ( .A(n_21), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_22), .A2(n_34), .B1(n_111), .B2(n_113), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_23), .A2(n_40), .B1(n_113), .B2(n_145), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_24), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_25), .B(n_178), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_26), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_28), .A2(n_67), .B1(n_105), .B2(n_127), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_29), .A2(n_33), .B1(n_105), .B2(n_149), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_31), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_32), .A2(n_42), .B1(n_145), .B2(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_34), .Y(n_635) );
INVx2_ASAP7_75t_L g528 ( .A(n_35), .Y(n_528) );
INVx1_ASAP7_75t_L g587 ( .A(n_35), .Y(n_587) );
INVx1_ASAP7_75t_L g557 ( .A(n_36), .Y(n_557) );
INVx2_ASAP7_75t_L g626 ( .A(n_37), .Y(n_626) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_38), .A2(n_59), .B1(n_488), .B2(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g564 ( .A(n_39), .Y(n_564) );
INVx1_ASAP7_75t_L g559 ( .A(n_43), .Y(n_559) );
BUFx3_ASAP7_75t_L g490 ( .A(n_44), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_45), .A2(n_56), .B1(n_111), .B2(n_167), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_46), .A2(n_58), .B1(n_105), .B2(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g546 ( .A(n_47), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_48), .A2(n_75), .B1(n_145), .B2(n_147), .Y(n_144) );
AND2x4_ASAP7_75t_L g82 ( .A(n_49), .B(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_49), .Y(n_595) );
INVx1_ASAP7_75t_L g119 ( .A(n_50), .Y(n_119) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_51), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_52), .Y(n_614) );
INVx1_ASAP7_75t_L g83 ( .A(n_53), .Y(n_83) );
INVx1_ASAP7_75t_L g566 ( .A(n_54), .Y(n_566) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_55), .Y(n_440) );
INVx1_ASAP7_75t_L g462 ( .A(n_57), .Y(n_462) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_60), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g87 ( .A(n_61), .Y(n_87) );
BUFx3_ASAP7_75t_L g610 ( .A(n_62), .Y(n_610) );
INVx1_ASAP7_75t_L g555 ( .A(n_63), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_64), .A2(n_74), .B1(n_113), .B2(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_65), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
INVx1_ASAP7_75t_L g443 ( .A(n_68), .Y(n_443) );
BUFx3_ASAP7_75t_L g447 ( .A(n_68), .Y(n_447) );
INVx1_ASAP7_75t_L g604 ( .A(n_69), .Y(n_604) );
INVx1_ASAP7_75t_L g485 ( .A(n_70), .Y(n_485) );
INVx2_ASAP7_75t_L g537 ( .A(n_70), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_71), .B(n_116), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_72), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_73), .B(n_146), .Y(n_219) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_75), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_430), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_84), .Y(n_80) );
AO31x2_ASAP7_75t_L g102 ( .A1(n_81), .A2(n_103), .A3(n_115), .B(n_120), .Y(n_102) );
INVx2_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_81), .A2(n_124), .A3(n_176), .B(n_184), .Y(n_175) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_81), .A2(n_141), .A3(n_199), .B(n_202), .Y(n_198) );
BUFx10_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_83), .Y(n_597) );
INVxp67_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AO21x1_ASAP7_75t_L g644 ( .A1(n_85), .A2(n_596), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_88), .Y(n_85) );
INVx6_ASAP7_75t_L g114 ( .A(n_86), .Y(n_114) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_86), .A2(n_149), .B(n_215), .C(n_216), .Y(n_214) );
BUFx8_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx3_ASAP7_75t_L g105 ( .A(n_92), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_92), .Y(n_106) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_92), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
INVx2_ASAP7_75t_L g128 ( .A(n_92), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_92), .Y(n_146) );
INVx1_ASAP7_75t_L g165 ( .A(n_92), .Y(n_165) );
INVx1_ASAP7_75t_L g180 ( .A(n_92), .Y(n_180) );
INVx1_ASAP7_75t_L g183 ( .A(n_92), .Y(n_183) );
BUFx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NOR2x1p5_ASAP7_75t_L g95 ( .A(n_96), .B(n_340), .Y(n_95) );
NAND4xp75_ASAP7_75t_L g96 ( .A(n_97), .B(n_285), .C(n_305), .D(n_321), .Y(n_96) );
NOR2x1p5_ASAP7_75t_SL g97 ( .A(n_98), .B(n_255), .Y(n_97) );
NAND4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_194), .C(n_232), .D(n_241), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_100), .B(n_155), .Y(n_99) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_122), .Y(n_100) );
AND2x4_ASAP7_75t_L g365 ( .A(n_101), .B(n_292), .Y(n_365) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_102), .Y(n_208) );
INVx2_ASAP7_75t_L g226 ( .A(n_102), .Y(n_226) );
AND2x2_ASAP7_75t_L g249 ( .A(n_102), .B(n_211), .Y(n_249) );
OR2x2_ASAP7_75t_L g304 ( .A(n_102), .B(n_123), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B1(n_110), .B2(n_114), .Y(n_103) );
INVx1_ASAP7_75t_L g147 ( .A(n_105), .Y(n_147) );
INVx4_ASAP7_75t_L g149 ( .A(n_105), .Y(n_149) );
INVx1_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_107), .A2(n_114), .B1(n_163), .B2(n_166), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_107), .A2(n_114), .B1(n_177), .B2(n_181), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_107), .A2(n_114), .B1(n_190), .B2(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g178 ( .A(n_112), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_114), .A2(n_126), .B1(n_129), .B2(n_131), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_114), .A2(n_144), .B1(n_148), .B2(n_150), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_114), .A2(n_150), .B1(n_200), .B2(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_114), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_117), .B(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_117), .B(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_117), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g212 ( .A(n_117), .Y(n_212) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
AND2x2_ASAP7_75t_L g222 ( .A(n_122), .B(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g372 ( .A(n_122), .B(n_249), .Y(n_372) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_139), .Y(n_122) );
OR2x2_ASAP7_75t_L g209 ( .A(n_123), .B(n_210), .Y(n_209) );
BUFx2_ASAP7_75t_L g240 ( .A(n_123), .Y(n_240) );
AND2x2_ASAP7_75t_L g246 ( .A(n_123), .B(n_140), .Y(n_246) );
INVx1_ASAP7_75t_L g264 ( .A(n_123), .Y(n_264) );
INVx2_ASAP7_75t_L g293 ( .A(n_123), .Y(n_293) );
AO31x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .A3(n_133), .B(n_135), .Y(n_123) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_SL g150 ( .A(n_132), .Y(n_150) );
AO31x2_ASAP7_75t_L g188 ( .A1(n_133), .A2(n_168), .A3(n_189), .B(n_192), .Y(n_188) );
INVx2_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_SL g220 ( .A(n_134), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx2_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_136), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
INVx2_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx3_ASAP7_75t_L g269 ( .A(n_139), .Y(n_269) );
INVx2_ASAP7_75t_L g274 ( .A(n_139), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_139), .B(n_225), .Y(n_279) );
AND2x2_ASAP7_75t_L g302 ( .A(n_139), .B(n_281), .Y(n_302) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_139), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_139), .B(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx2_ASAP7_75t_L g291 ( .A(n_140), .Y(n_291) );
AND2x2_ASAP7_75t_L g339 ( .A(n_140), .B(n_293), .Y(n_339) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_143), .A3(n_151), .B(n_153), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AO31x2_ASAP7_75t_L g161 ( .A1(n_151), .A2(n_162), .A3(n_168), .B(n_170), .Y(n_161) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_173), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_157), .B(n_283), .Y(n_330) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_158), .B(n_283), .Y(n_327) );
INVx1_ASAP7_75t_L g428 ( .A(n_158), .Y(n_428) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g378 ( .A(n_159), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g231 ( .A(n_160), .Y(n_231) );
OR2x2_ASAP7_75t_L g312 ( .A(n_160), .B(n_187), .Y(n_312) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g254 ( .A(n_161), .Y(n_254) );
AND2x4_ASAP7_75t_L g260 ( .A(n_161), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_172), .B(n_193), .Y(n_192) );
AOI32xp33_ASAP7_75t_L g398 ( .A1(n_173), .A2(n_301), .A3(n_399), .B1(n_401), .B2(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g347 ( .A(n_174), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_186), .Y(n_174) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
OR2x2_ASAP7_75t_L g229 ( .A(n_175), .B(n_188), .Y(n_229) );
INVx1_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
AND2x2_ASAP7_75t_L g253 ( .A(n_175), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g259 ( .A(n_175), .Y(n_259) );
INVx2_ASAP7_75t_L g284 ( .A(n_175), .Y(n_284) );
AND2x2_ASAP7_75t_L g403 ( .A(n_175), .B(n_198), .Y(n_403) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_186), .B(n_236), .Y(n_323) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g197 ( .A(n_188), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g252 ( .A(n_188), .Y(n_252) );
INVx2_ASAP7_75t_L g261 ( .A(n_188), .Y(n_261) );
AND2x4_ASAP7_75t_L g283 ( .A(n_188), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_188), .Y(n_375) );
AOI22x1_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_204), .B1(n_222), .B2(n_227), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_197), .B(n_353), .C(n_354), .D(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_197), .B(n_253), .Y(n_383) );
INVx4_ASAP7_75t_SL g236 ( .A(n_198), .Y(n_236) );
BUFx2_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_198), .B(n_244), .Y(n_362) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g324 ( .A(n_206), .B(n_273), .Y(n_324) );
NOR2x1_ASAP7_75t_L g206 ( .A(n_207), .B(n_209), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x4_ASAP7_75t_L g247 ( .A(n_210), .B(n_225), .Y(n_247) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_211), .B(n_226), .Y(n_271) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_221), .Y(n_211) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_212), .A2(n_213), .B(n_221), .Y(n_266) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .B(n_220), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_223), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g289 ( .A(n_223), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g328 ( .A(n_224), .B(n_246), .Y(n_328) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g371 ( .A(n_226), .B(n_281), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_227), .A2(n_344), .B1(n_346), .B2(n_349), .C(n_351), .Y(n_343) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g237 ( .A(n_229), .Y(n_237) );
OR2x2_ASAP7_75t_L g337 ( .A(n_229), .B(n_276), .Y(n_337) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_238), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_233), .A2(n_359), .B1(n_363), .B2(n_366), .Y(n_358) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
AND2x4_ASAP7_75t_L g282 ( .A(n_234), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g394 ( .A(n_234), .B(n_312), .Y(n_394) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g242 ( .A(n_236), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_236), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g317 ( .A(n_236), .B(n_254), .Y(n_317) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_236), .Y(n_334) );
INVx1_ASAP7_75t_L g348 ( .A(n_236), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_236), .B(n_261), .Y(n_391) );
AND2x4_ASAP7_75t_L g298 ( .A(n_237), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g296 ( .A(n_239), .Y(n_296) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_240), .B(n_281), .Y(n_280) );
NAND2x1_ASAP7_75t_L g400 ( .A(n_240), .B(n_302), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B1(n_248), .B2(n_250), .Y(n_241) );
AND2x2_ASAP7_75t_L g267 ( .A(n_242), .B(n_260), .Y(n_267) );
INVx1_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
AND2x2_ASAP7_75t_L g415 ( .A(n_242), .B(n_276), .Y(n_415) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x4_ASAP7_75t_SL g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g248 ( .A(n_246), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g388 ( .A(n_246), .Y(n_388) );
AND2x2_ASAP7_75t_L g405 ( .A(n_246), .B(n_265), .Y(n_405) );
AND2x2_ASAP7_75t_L g421 ( .A(n_246), .B(n_371), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_247), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g344 ( .A(n_247), .B(n_345), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_247), .A2(n_337), .B1(n_352), .B2(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g307 ( .A(n_249), .Y(n_307) );
AND2x2_ASAP7_75t_L g338 ( .A(n_249), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_249), .B(n_345), .Y(n_367) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g373 ( .A(n_253), .B(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_253), .A2(n_277), .B1(n_382), .B2(n_384), .Y(n_381) );
INVx3_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
AND2x2_ASAP7_75t_L g408 ( .A(n_254), .B(n_261), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_272), .Y(n_255) );
AOI32xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .A3(n_265), .B1(n_267), .B2(n_268), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_259), .Y(n_354) );
INVx1_ASAP7_75t_L g379 ( .A(n_259), .Y(n_379) );
INVx3_ASAP7_75t_L g335 ( .A(n_260), .Y(n_335) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_263), .A2(n_411), .B1(n_412), .B2(n_413), .C(n_414), .Y(n_410) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g387 ( .A(n_265), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g423 ( .A(n_265), .B(n_384), .Y(n_423) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g281 ( .A(n_266), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g295 ( .A(n_268), .B(n_296), .Y(n_295) );
AO22x1_ASAP7_75t_L g325 ( .A1(n_268), .A2(n_326), .B1(n_328), .B2(n_329), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_268), .B(n_296), .Y(n_429) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g345 ( .A(n_269), .Y(n_345) );
INVx1_ASAP7_75t_L g355 ( .A(n_269), .Y(n_355) );
AND2x2_ASAP7_75t_L g275 ( .A(n_270), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_271), .Y(n_357) );
INVx1_ASAP7_75t_L g397 ( .A(n_271), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_277), .C(n_282), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2x1p5_ASAP7_75t_L g384 ( .A(n_274), .B(n_304), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_275), .B(n_334), .Y(n_411) );
AOI31xp33_ASAP7_75t_L g294 ( .A1(n_276), .A2(n_295), .A3(n_297), .B(n_300), .Y(n_294) );
INVx4_ASAP7_75t_L g353 ( .A(n_276), .Y(n_353) );
OR2x2_ASAP7_75t_L g390 ( .A(n_276), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x4_ASAP7_75t_L g292 ( .A(n_281), .B(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_317), .Y(n_319) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_286), .B(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g412 ( .A(n_289), .Y(n_412) );
INVx1_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
AND2x2_ASAP7_75t_L g349 ( .A(n_292), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .A3(n_309), .B1(n_313), .B2(n_316), .C1(n_318), .C2(n_320), .Y(n_306) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI211x1_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_325), .C(n_331), .Y(n_321) );
INVx1_ASAP7_75t_L g426 ( .A(n_322), .Y(n_426) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OA21x2_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_336), .B(n_338), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g401 ( .A(n_335), .Y(n_401) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp33_ASAP7_75t_L g396 ( .A(n_339), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_409), .Y(n_340) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_376), .C(n_392), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_358), .C(n_368), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_345), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_349), .A2(n_405), .B(n_406), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_353), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_353), .B(n_403), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_354), .B(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_355), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g414 ( .A1(n_365), .A2(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B(n_381), .C(n_385), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_387), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_398), .C(n_404), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_403), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g420 ( .A(n_408), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_418), .C(n_425), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_422), .B(n_424), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_R g425 ( .A1(n_426), .A2(n_427), .B(n_429), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_593), .B1(n_598), .B2(n_640), .C(n_641), .Y(n_430) );
INVx1_ASAP7_75t_L g640 ( .A(n_432), .Y(n_640) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_SL g433 ( .A(n_434), .B(n_486), .C(n_532), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_451), .A3(n_471), .B(n_479), .Y(n_434) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_442), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
BUFx4f_ASAP7_75t_L g542 ( .A(n_438), .Y(n_542) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_L g450 ( .A(n_440), .Y(n_450) );
NAND2x1_ASAP7_75t_L g455 ( .A(n_440), .B(n_441), .Y(n_455) );
AND2x2_ASAP7_75t_L g460 ( .A(n_440), .B(n_441), .Y(n_460) );
INVx1_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
AND2x2_ASAP7_75t_L g477 ( .A(n_440), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g552 ( .A(n_440), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_441), .B(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
INVx2_ASAP7_75t_L g478 ( .A(n_441), .Y(n_478) );
OR2x2_ASAP7_75t_L g551 ( .A(n_441), .B(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g476 ( .A(n_442), .B(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
AND2x2_ASAP7_75t_L g457 ( .A(n_445), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g473 ( .A(n_446), .Y(n_473) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
AND2x4_ASAP7_75t_L g468 ( .A(n_447), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g562 ( .A(n_447), .B(n_481), .Y(n_562) );
INVx8_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx5_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_455), .Y(n_554) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_466), .B2(n_467), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_462), .A2(n_504), .B1(n_509), .B2(n_510), .Y(n_503) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g531 ( .A(n_484), .Y(n_531) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI31xp33_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_497), .A3(n_515), .B(n_525), .Y(n_486) );
OR2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_493), .Y(n_488) );
OR2x4_ASAP7_75t_L g495 ( .A(n_489), .B(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
BUFx4f_ASAP7_75t_L g589 ( .A(n_489), .Y(n_589) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_L g500 ( .A(n_490), .B(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_490), .Y(n_508) );
INVx2_ASAP7_75t_L g521 ( .A(n_490), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_490), .B(n_502), .Y(n_524) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g520 ( .A(n_492), .Y(n_520) );
INVx1_ASAP7_75t_L g496 ( .A(n_493), .Y(n_496) );
AND2x4_ASAP7_75t_L g514 ( .A(n_493), .B(n_500), .Y(n_514) );
OR2x6_ASAP7_75t_L g522 ( .A(n_493), .B(n_523), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_493), .B(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g624 ( .A(n_493), .B(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g506 ( .A(n_494), .Y(n_506) );
NAND2xp33_ASAP7_75t_SL g570 ( .A(n_494), .B(n_528), .Y(n_570) );
AND2x2_ASAP7_75t_L g517 ( .A(n_496), .B(n_518), .Y(n_517) );
NAND3xp33_ASAP7_75t_SL g497 ( .A(n_498), .B(n_503), .C(n_513), .Y(n_497) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g512 ( .A(n_502), .Y(n_512) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g510 ( .A(n_505), .B(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_508), .B(n_512), .Y(n_575) );
INVx2_ASAP7_75t_L g623 ( .A(n_508), .Y(n_623) );
BUFx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
CKINVDCx8_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g581 ( .A(n_524), .Y(n_581) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g625 ( .A(n_528), .Y(n_625) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_531), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g569 ( .A(n_531), .B(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_567), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_539), .A3(n_547), .B1(n_556), .B2(n_560), .B3(n_563), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
OR2x2_ASAP7_75t_L g585 ( .A(n_536), .B(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_543), .B2(n_546), .Y(n_539) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_540), .A2(n_557), .B1(n_572), .B2(n_574), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_541), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g565 ( .A(n_545), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_546), .A2(n_559), .B1(n_589), .B2(n_590), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_553), .B2(n_555), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_548), .A2(n_564), .B1(n_577), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_549), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_556) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_554), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_555), .A2(n_566), .B1(n_583), .B2(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI33xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .A3(n_576), .B1(n_582), .B2(n_585), .B3(n_588), .Y(n_567) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g631 ( .A(n_570), .Y(n_631) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_575), .Y(n_592) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g584 ( .A(n_580), .Y(n_584) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g633 ( .A(n_595), .Y(n_633) );
BUFx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_597), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g645 ( .A(n_597), .B(n_633), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_616), .B1(n_634), .B2(n_636), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_599), .A2(n_617), .B1(n_634), .B2(n_643), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_611), .B1(n_612), .B2(n_615), .Y(n_605) );
INVx1_ASAP7_75t_L g615 ( .A(n_606), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
CKINVDCx14_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx12f_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx8_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_626), .B(n_627), .C(n_632), .Y(n_619) );
AND2x2_ASAP7_75t_L g639 ( .A(n_620), .B(n_627), .Y(n_639) );
INVx4_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x6_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_622), .B(n_628), .C(n_631), .Y(n_627) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx3_ASAP7_75t_L g630 ( .A(n_626), .Y(n_630) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g638 ( .A(n_632), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_634), .A2(n_640), .B1(n_642), .B2(n_644), .Y(n_641) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g643 ( .A(n_636), .Y(n_643) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
endmodule