module real_aes_2148_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g225 ( .A(n_0), .B(n_132), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_1), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_2), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_3), .B(n_121), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_4), .B(n_130), .Y(n_466) );
INVx1_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_6), .B(n_121), .Y(n_178) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_7), .B(n_127), .Y(n_171) );
INVx1_ASAP7_75t_L g151 ( .A(n_8), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_9), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_10), .Y(n_728) );
AND2x2_ASAP7_75t_L g176 ( .A(n_11), .B(n_111), .Y(n_176) );
AND2x2_ASAP7_75t_L g459 ( .A(n_12), .B(n_168), .Y(n_459) );
AND2x2_ASAP7_75t_L g468 ( .A(n_13), .B(n_143), .Y(n_468) );
INVx2_ASAP7_75t_L g112 ( .A(n_14), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_15), .B(n_130), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_16), .Y(n_425) );
AOI221x1_ASAP7_75t_L g165 ( .A1(n_17), .A2(n_115), .B1(n_166), .B2(n_168), .C(n_170), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_18), .B(n_121), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_19), .B(n_121), .Y(n_506) );
INVx1_ASAP7_75t_L g428 ( .A(n_20), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_21), .A2(n_89), .B1(n_121), .B2(n_153), .Y(n_447) );
AOI221xp5_ASAP7_75t_SL g114 ( .A1(n_22), .A2(n_36), .B1(n_115), .B2(n_121), .C(n_128), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_23), .A2(n_115), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_24), .B(n_132), .Y(n_181) );
OR2x2_ASAP7_75t_L g113 ( .A(n_25), .B(n_88), .Y(n_113) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_25), .A2(n_88), .B(n_112), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_26), .B(n_130), .Y(n_142) );
INVxp67_ASAP7_75t_L g164 ( .A(n_27), .Y(n_164) );
AND2x2_ASAP7_75t_L g214 ( .A(n_28), .B(n_110), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_29), .A2(n_115), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_30), .A2(n_168), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_31), .B(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_32), .A2(n_115), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_33), .B(n_130), .Y(n_501) );
AND2x2_ASAP7_75t_L g116 ( .A(n_34), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g127 ( .A(n_34), .B(n_120), .Y(n_127) );
INVx1_ASAP7_75t_L g160 ( .A(n_34), .Y(n_160) );
OR2x6_ASAP7_75t_L g426 ( .A(n_35), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_37), .B(n_121), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_38), .A2(n_81), .B1(n_115), .B2(n_158), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_39), .B(n_130), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_40), .B(n_121), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_41), .B(n_132), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_42), .A2(n_115), .B(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_43), .A2(n_71), .B1(n_720), .B2(n_721), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_43), .Y(n_720) );
AND2x2_ASAP7_75t_L g228 ( .A(n_44), .B(n_110), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_45), .B(n_132), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_46), .B(n_110), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_47), .B(n_121), .Y(n_518) );
INVx1_ASAP7_75t_L g119 ( .A(n_48), .Y(n_119) );
INVx1_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_49), .B(n_130), .Y(n_457) );
AND2x2_ASAP7_75t_L g487 ( .A(n_50), .B(n_110), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_51), .B(n_121), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_52), .B(n_132), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_53), .B(n_132), .Y(n_500) );
AND2x2_ASAP7_75t_L g192 ( .A(n_54), .B(n_110), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_55), .B(n_121), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_56), .B(n_130), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_57), .B(n_121), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_58), .A2(n_115), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_59), .B(n_111), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_60), .B(n_132), .Y(n_189) );
AND2x2_ASAP7_75t_L g512 ( .A(n_61), .B(n_111), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_62), .A2(n_115), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_63), .B(n_130), .Y(n_182) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_64), .B(n_143), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_65), .B(n_132), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_66), .A2(n_101), .B1(n_729), .B2(n_740), .C1(n_755), .C2(n_757), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_66), .A2(n_69), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_66), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_67), .B(n_132), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_68), .A2(n_91), .B1(n_115), .B2(n_158), .Y(n_448) );
INVx1_ASAP7_75t_L g744 ( .A(n_69), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_70), .B(n_130), .Y(n_509) );
INVx1_ASAP7_75t_L g721 ( .A(n_71), .Y(n_721) );
INVx1_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_73), .B(n_132), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_74), .A2(n_115), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_75), .A2(n_115), .B(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_76), .A2(n_115), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g503 ( .A(n_77), .B(n_111), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_78), .B(n_110), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_79), .B(n_121), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_80), .A2(n_83), .B1(n_121), .B2(n_153), .Y(n_197) );
INVx1_ASAP7_75t_L g429 ( .A(n_82), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_84), .B(n_132), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_85), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g480 ( .A(n_86), .B(n_143), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_87), .A2(n_115), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_90), .B(n_130), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_92), .A2(n_115), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_93), .B(n_130), .Y(n_478) );
INVxp67_ASAP7_75t_L g167 ( .A(n_94), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_95), .B(n_121), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_96), .B(n_130), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_97), .A2(n_115), .B(n_140), .Y(n_139) );
BUFx2_ASAP7_75t_L g511 ( .A(n_98), .Y(n_511) );
BUFx2_ASAP7_75t_L g737 ( .A(n_99), .Y(n_737) );
BUFx2_ASAP7_75t_SL g761 ( .A(n_99), .Y(n_761) );
OAI222xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_718), .B1(n_719), .B2(n_722), .C1(n_725), .C2(n_728), .Y(n_101) );
OA22x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_421), .B1(n_430), .B2(n_434), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_104), .A2(n_430), .B1(n_435), .B2(n_724), .Y(n_723) );
INVx4_ASAP7_75t_L g747 ( .A(n_104), .Y(n_747) );
OR2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_334), .Y(n_104) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_244), .C(n_284), .Y(n_105) );
O2A1O1Ixp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_146), .B(n_173), .C(n_200), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_107), .B(n_249), .Y(n_283) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_135), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g219 ( .A(n_109), .Y(n_219) );
INVx2_ASAP7_75t_L g235 ( .A(n_109), .Y(n_235) );
OR2x2_ASAP7_75t_L g247 ( .A(n_109), .B(n_136), .Y(n_247) );
AND2x2_ASAP7_75t_L g261 ( .A(n_109), .B(n_220), .Y(n_261) );
INVx1_ASAP7_75t_L g289 ( .A(n_109), .Y(n_289) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_109), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_109), .B(n_136), .Y(n_395) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_134), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_110), .Y(n_191) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_110), .A2(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_110), .A2(n_475), .B(n_476), .Y(n_474) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x4_ASAP7_75t_L g152 ( .A(n_112), .B(n_113), .Y(n_152) );
AND2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
BUFx3_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
AND2x6_ASAP7_75t_L g132 ( .A(n_117), .B(n_123), .Y(n_132) );
INVx2_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
AND2x4_ASAP7_75t_L g158 ( .A(n_118), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g130 ( .A(n_119), .B(n_125), .Y(n_130) );
INVx2_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g172 ( .A(n_122), .Y(n_172) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_131), .B(n_133), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_132), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_133), .A2(n_141), .B(n_142), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_133), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_133), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_133), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_133), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_133), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_133), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_133), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_133), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_133), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_133), .A2(n_521), .B(n_522), .Y(n_520) );
OR2x2_ASAP7_75t_L g216 ( .A(n_135), .B(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_135), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_135), .B(n_218), .Y(n_356) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g146 ( .A(n_136), .B(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g215 ( .A(n_136), .B(n_148), .Y(n_215) );
OR2x2_ASAP7_75t_L g234 ( .A(n_136), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g263 ( .A(n_136), .Y(n_263) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_136), .B(n_148), .Y(n_302) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_136), .Y(n_306) );
OR2x2_ASAP7_75t_L g323 ( .A(n_136), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g333 ( .A(n_136), .B(n_240), .Y(n_333) );
INVx1_ASAP7_75t_L g362 ( .A(n_136), .Y(n_362) );
OR2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_145), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_143), .Y(n_137) );
INVx2_ASAP7_75t_SL g195 ( .A(n_143), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_143), .A2(n_506), .B(n_507), .Y(n_505) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_146), .B(n_291), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_147), .B(n_220), .Y(n_237) );
AND2x2_ASAP7_75t_L g249 ( .A(n_147), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g267 ( .A(n_147), .B(n_234), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_147), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g240 ( .A(n_148), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g262 ( .A(n_148), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g297 ( .A(n_148), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_148), .B(n_220), .Y(n_321) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_165), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B1(n_158), .B2(n_163), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_152), .B(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_152), .B(n_167), .Y(n_166) );
NOR3xp33_ASAP7_75t_L g170 ( .A(n_152), .B(n_171), .C(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_152), .A2(n_518), .B(n_519), .Y(n_517) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_157), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g496 ( .A(n_168), .Y(n_496) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21x1_ASAP7_75t_L g221 ( .A1(n_169), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_169), .A2(n_453), .B(n_459), .Y(n_452) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_183), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_174), .B(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g270 ( .A(n_174), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_174), .B(n_184), .Y(n_275) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_174), .B(n_291), .C(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g338 ( .A(n_174), .B(n_243), .Y(n_338) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g205 ( .A(n_175), .B(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_SL g242 ( .A(n_175), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
OR2x2_ASAP7_75t_L g281 ( .A(n_175), .B(n_271), .Y(n_281) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_175), .Y(n_298) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_175), .B(n_204), .Y(n_316) );
AND2x4_ASAP7_75t_L g331 ( .A(n_175), .B(n_207), .Y(n_331) );
AND2x2_ASAP7_75t_L g345 ( .A(n_175), .B(n_184), .Y(n_345) );
OR2x2_ASAP7_75t_L g366 ( .A(n_175), .B(n_193), .Y(n_366) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
AND2x2_ASAP7_75t_L g420 ( .A(n_183), .B(n_298), .Y(n_420) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
AND2x4_ASAP7_75t_L g243 ( .A(n_184), .B(n_206), .Y(n_243) );
INVx2_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
AND2x2_ASAP7_75t_L g259 ( .A(n_184), .B(n_204), .Y(n_259) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_184), .Y(n_292) );
OR2x2_ASAP7_75t_L g315 ( .A(n_184), .B(n_207), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_184), .B(n_207), .Y(n_318) );
INVx1_ASAP7_75t_L g327 ( .A(n_184), .Y(n_327) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_191), .A2(n_208), .B(n_214), .Y(n_207) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_191), .A2(n_208), .B(n_214), .Y(n_271) );
AOI21x1_ASAP7_75t_L g461 ( .A1(n_191), .A2(n_462), .B(n_468), .Y(n_461) );
AND2x2_ASAP7_75t_L g230 ( .A(n_193), .B(n_207), .Y(n_230) );
BUFx2_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
AND2x2_ASAP7_75t_L g374 ( .A(n_193), .B(n_254), .Y(n_374) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_194), .Y(n_204) );
AOI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_215), .B1(n_216), .B2(n_229), .C(n_231), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_205), .Y(n_202) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_203), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_203), .B(n_270), .Y(n_310) );
OR2x2_ASAP7_75t_L g322 ( .A(n_203), .B(n_318), .Y(n_322) );
OR2x2_ASAP7_75t_L g325 ( .A(n_203), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g414 ( .A(n_203), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g253 ( .A(n_204), .B(n_254), .Y(n_253) );
OA33x2_ASAP7_75t_L g286 ( .A1(n_204), .A2(n_247), .A3(n_287), .B1(n_290), .B2(n_293), .B3(n_296), .Y(n_286) );
OR2x2_ASAP7_75t_L g317 ( .A(n_204), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g341 ( .A(n_204), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g349 ( .A(n_204), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g369 ( .A(n_204), .B(n_243), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_204), .B(n_258), .Y(n_407) );
INVx2_ASAP7_75t_L g277 ( .A(n_205), .Y(n_277) );
AOI322xp5_ASAP7_75t_L g347 ( .A1(n_205), .A2(n_260), .A3(n_348), .B1(n_351), .B2(n_352), .C1(n_354), .C2(n_356), .Y(n_347) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_207), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_213), .Y(n_208) );
OR2x2_ASAP7_75t_L g329 ( .A(n_215), .B(n_308), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_215), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g402 ( .A(n_215), .Y(n_402) );
INVx1_ASAP7_75t_SL g268 ( .A(n_216), .Y(n_268) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g301 ( .A(n_218), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g241 ( .A(n_220), .Y(n_241) );
INVx1_ASAP7_75t_L g250 ( .A(n_220), .Y(n_250) );
INVx1_ASAP7_75t_L g291 ( .A(n_220), .Y(n_291) );
OR2x2_ASAP7_75t_L g308 ( .A(n_220), .B(n_235), .Y(n_308) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_220), .Y(n_383) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_SL g352 ( .A(n_230), .B(n_353), .Y(n_352) );
OAI21xp5_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_238), .B(n_242), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_232), .A2(n_306), .B(n_307), .C(n_309), .Y(n_305) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_236), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g370 ( .A(n_234), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_235), .Y(n_239) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g394 ( .A(n_237), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_240), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g371 ( .A(n_240), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_240), .B(n_362), .Y(n_379) );
INVx3_ASAP7_75t_SL g304 ( .A(n_243), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B1(n_255), .B2(n_260), .C(n_264), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_250), .Y(n_295) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_253), .A2(n_280), .B(n_352), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_253), .B(n_331), .Y(n_384) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_254), .Y(n_272) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_258), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g393 ( .A(n_258), .B(n_315), .Y(n_393) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g342 ( .A(n_261), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .B(n_273), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx2_ASAP7_75t_L g415 ( .A(n_270), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_271), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g344 ( .A(n_271), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_272), .B(n_294), .Y(n_293) );
OAI31xp33_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_276), .A3(n_278), .B(n_282), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_277), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g355 ( .A(n_279), .B(n_281), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_279), .B(n_331), .Y(n_410) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR5xp2_ASAP7_75t_L g284 ( .A(n_285), .B(n_299), .C(n_311), .D(n_320), .E(n_328), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_289), .B(n_291), .Y(n_324) );
INVx1_ASAP7_75t_L g364 ( .A(n_289), .Y(n_364) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_289), .Y(n_401) );
INVx1_ASAP7_75t_L g353 ( .A(n_292), .Y(n_353) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI321xp33_ASAP7_75t_L g336 ( .A1(n_297), .A2(n_337), .A3(n_339), .B1(n_343), .B2(n_346), .C(n_347), .Y(n_336) );
INVx1_ASAP7_75t_L g390 ( .A(n_298), .Y(n_390) );
OAI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B(n_305), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_301), .A2(n_374), .B1(n_381), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g409 ( .A(n_302), .B(n_383), .Y(n_409) );
INVx1_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_317), .B(n_319), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_318), .A2(n_329), .B1(n_330), .B2(n_332), .Y(n_328) );
INVx1_ASAP7_75t_L g391 ( .A(n_318), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_323), .B2(n_325), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_327), .B(n_331), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_329), .A2(n_406), .B1(n_408), .B2(n_410), .C(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_329), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_330), .A2(n_387), .B1(n_394), .B2(n_396), .C(n_397), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_332), .A2(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_385), .Y(n_334) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_357), .C(n_375), .Y(n_335) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_338), .Y(n_404) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g403 ( .A(n_346), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_348), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_365), .B(n_367), .Y(n_359) );
INVxp67_ASAP7_75t_L g417 ( .A(n_360), .Y(n_417) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g372 ( .A(n_363), .Y(n_372) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_372), .B2(n_373), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_380), .Y(n_375) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g418 ( .A(n_381), .Y(n_418) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_405), .C(n_416), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_392), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_403), .B(n_404), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_409), .A2(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
INVx4_ASAP7_75t_SL g724 ( .A(n_422), .Y(n_724) );
INVx3_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
AND2x6_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OR2x6_ASAP7_75t_SL g432 ( .A(n_425), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g727 ( .A(n_425), .B(n_426), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_425), .B(n_433), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_426), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
CKINVDCx11_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
INVx4_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OR2x6_ASAP7_75t_L g435 ( .A(n_436), .B(n_655), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_571), .C(n_608), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_539), .C(n_554), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_484), .B1(n_513), .B2(n_525), .C(n_526), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_469), .Y(n_440) );
OAI22xp33_ASAP7_75t_SL g599 ( .A1(n_441), .A2(n_563), .B1(n_600), .B2(n_603), .Y(n_599) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .Y(n_441) );
OAI21xp33_ASAP7_75t_SL g609 ( .A1(n_442), .A2(n_610), .B(n_616), .Y(n_609) );
OR2x2_ASAP7_75t_L g638 ( .A(n_442), .B(n_471), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_442), .B(n_558), .Y(n_639) );
INVx2_ASAP7_75t_L g670 ( .A(n_442), .Y(n_670) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_443), .B(n_530), .Y(n_651) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g525 ( .A(n_444), .B(n_452), .Y(n_525) );
BUFx3_ASAP7_75t_L g551 ( .A(n_444), .Y(n_551) );
AND2x2_ASAP7_75t_L g687 ( .A(n_444), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g710 ( .A(n_444), .B(n_472), .Y(n_710) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
AND2x4_ASAP7_75t_L g483 ( .A(n_445), .B(n_446), .Y(n_483) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_450), .B(n_472), .Y(n_630) );
INVx1_ASAP7_75t_L g667 ( .A(n_450), .Y(n_667) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
AND2x2_ASAP7_75t_L g482 ( .A(n_451), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g688 ( .A(n_451), .Y(n_688) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g531 ( .A(n_452), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_452), .B(n_460), .Y(n_532) );
AND2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_473), .Y(n_553) );
AND2x2_ASAP7_75t_L g635 ( .A(n_452), .B(n_461), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_458), .Y(n_453) );
AND2x4_ASAP7_75t_SL g528 ( .A(n_460), .B(n_473), .Y(n_528) );
INVx1_ASAP7_75t_L g559 ( .A(n_460), .Y(n_559) );
INVx2_ASAP7_75t_L g567 ( .A(n_460), .Y(n_567) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_460), .Y(n_591) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_461), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_482), .Y(n_469) );
AND2x2_ASAP7_75t_L g706 ( .A(n_470), .B(n_569), .Y(n_706) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_472), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g617 ( .A(n_472), .B(n_532), .Y(n_617) );
AND2x2_ASAP7_75t_L g634 ( .A(n_472), .B(n_635), .Y(n_634) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g558 ( .A(n_473), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
AND2x2_ASAP7_75t_L g618 ( .A(n_473), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g625 ( .A(n_473), .B(n_626), .Y(n_625) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_473), .B(n_531), .Y(n_640) );
BUFx2_ASAP7_75t_L g650 ( .A(n_473), .Y(n_650) );
AND2x2_ASAP7_75t_L g675 ( .A(n_473), .B(n_635), .Y(n_675) );
AND2x2_ASAP7_75t_L g696 ( .A(n_473), .B(n_697), .Y(n_696) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_480), .Y(n_473) );
INVx1_ASAP7_75t_L g627 ( .A(n_481), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_482), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g657 ( .A(n_482), .B(n_528), .Y(n_657) );
INVx3_ASAP7_75t_L g564 ( .A(n_483), .Y(n_564) );
AND2x2_ASAP7_75t_L g697 ( .A(n_483), .B(n_619), .Y(n_697) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_485), .A2(n_527), .B1(n_532), .B2(n_533), .Y(n_526) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
INVx4_ASAP7_75t_L g524 ( .A(n_486), .Y(n_524) );
INVx2_ASAP7_75t_L g561 ( .A(n_486), .Y(n_561) );
NAND2x1_ASAP7_75t_L g587 ( .A(n_486), .B(n_504), .Y(n_587) );
OR2x2_ASAP7_75t_L g602 ( .A(n_486), .B(n_537), .Y(n_602) );
OR2x2_ASAP7_75t_SL g629 ( .A(n_486), .B(n_601), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_486), .B(n_516), .Y(n_642) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_486), .Y(n_663) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g542 ( .A(n_494), .Y(n_542) );
AND2x2_ASAP7_75t_L g674 ( .A(n_494), .B(n_648), .Y(n_674) );
NOR2x1_ASAP7_75t_SL g494 ( .A(n_495), .B(n_504), .Y(n_494) );
AND2x2_ASAP7_75t_L g515 ( .A(n_495), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g691 ( .A(n_495), .B(n_614), .Y(n_691) );
AO21x1_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B(n_503), .Y(n_495) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_496), .A2(n_497), .B(n_503), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
OR2x2_ASAP7_75t_L g523 ( .A(n_504), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g534 ( .A(n_504), .B(n_524), .Y(n_534) );
AND2x2_ASAP7_75t_L g580 ( .A(n_504), .B(n_537), .Y(n_580) );
OR2x2_ASAP7_75t_L g601 ( .A(n_504), .B(n_516), .Y(n_601) );
INVx2_ASAP7_75t_SL g607 ( .A(n_504), .Y(n_607) );
AND2x2_ASAP7_75t_L g613 ( .A(n_504), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g623 ( .A(n_504), .B(n_606), .Y(n_623) );
BUFx2_ASAP7_75t_L g645 ( .A(n_504), .Y(n_645) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .Y(n_504) );
INVx2_ASAP7_75t_L g692 ( .A(n_513), .Y(n_692) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
OR2x2_ASAP7_75t_L g717 ( .A(n_514), .B(n_561), .Y(n_717) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_515), .B(n_524), .Y(n_583) );
AND2x2_ASAP7_75t_L g654 ( .A(n_515), .B(n_534), .Y(n_654) );
INVx1_ASAP7_75t_L g536 ( .A(n_516), .Y(n_536) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
INVx1_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
INVx2_ASAP7_75t_L g614 ( .A(n_516), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_524), .B(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g604 ( .A(n_524), .Y(n_604) );
INVx2_ASAP7_75t_SL g680 ( .A(n_525), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_527), .A2(n_582), .B1(n_584), .B2(n_588), .Y(n_581) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g708 ( .A(n_528), .B(n_564), .Y(n_708) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_530), .B(n_574), .Y(n_653) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g619 ( .A(n_531), .B(n_567), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_532), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g562 ( .A(n_533), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_533), .A2(n_677), .B1(n_681), .B2(n_683), .C(n_685), .Y(n_676) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g546 ( .A(n_534), .B(n_547), .Y(n_546) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_534), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_534), .B(n_577), .Y(n_632) );
INVx1_ASAP7_75t_SL g628 ( .A(n_535), .Y(n_628) );
AOI221xp5_ASAP7_75t_SL g656 ( .A1(n_535), .A2(n_546), .B1(n_657), .B2(n_658), .C(n_661), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_535), .A2(n_607), .A3(n_634), .B1(n_690), .B2(n_692), .C1(n_693), .C2(n_696), .Y(n_689) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
BUFx2_ASAP7_75t_L g556 ( .A(n_536), .Y(n_556) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
INVx2_ASAP7_75t_L g606 ( .A(n_537), .Y(n_606) );
AND2x2_ASAP7_75t_L g647 ( .A(n_537), .B(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OA21x2_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_546), .B(n_549), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_540), .A2(n_710), .B(n_711), .C(n_715), .Y(n_709) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OR2x2_ASAP7_75t_L g598 ( .A(n_542), .B(n_560), .Y(n_598) );
OR2x2_ASAP7_75t_L g682 ( .A(n_542), .B(n_577), .Y(n_682) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g622 ( .A(n_544), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g700 ( .A(n_547), .Y(n_700) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OR2x2_ASAP7_75t_L g555 ( .A(n_551), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_591), .Y(n_590) );
OAI322xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .A3(n_560), .B1(n_562), .B2(n_563), .C1(n_568), .C2(n_570), .Y(n_554) );
INVx1_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
OR2x2_ASAP7_75t_L g568 ( .A(n_557), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_557), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g579 ( .A(n_561), .B(n_580), .Y(n_579) );
OAI32xp33_ASAP7_75t_L g624 ( .A1(n_561), .A2(n_625), .A3(n_628), .B1(n_629), .B2(n_630), .Y(n_624) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g569 ( .A(n_564), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_564), .B(n_627), .Y(n_626) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_564), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g690 ( .A(n_564), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_569), .B(n_635), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_592), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_581), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g641 ( .A(n_580), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_583), .A2(n_603), .B1(n_705), .B2(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_585), .A2(n_632), .B(n_633), .C(n_636), .Y(n_631) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx3_ASAP7_75t_L g713 ( .A(n_587), .Y(n_713) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g594 ( .A(n_591), .Y(n_594) );
AO21x1_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_599), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g659 ( .A(n_594), .Y(n_659) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_600), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g615 ( .A(n_602), .Y(n_615) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g672 ( .A(n_605), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_631), .C(n_643), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_612), .A2(n_674), .B(n_675), .Y(n_673) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g648 ( .A(n_614), .Y(n_648) );
O2A1O1Ixp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_618), .B(n_620), .C(n_624), .Y(n_616) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_626), .Y(n_716) );
INVx2_ASAP7_75t_L g701 ( .A(n_629), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_630), .A2(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g695 ( .A(n_635), .Y(n_695) );
OAI31xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .A3(n_640), .B(n_641), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g714 ( .A(n_642), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_649), .B(n_652), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g664 ( .A(n_647), .Y(n_664) );
AOI21xp33_ASAP7_75t_SL g711 ( .A1(n_649), .A2(n_712), .B(n_714), .Y(n_711) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx2_ASAP7_75t_L g679 ( .A(n_650), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_650), .B(n_670), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_650), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g660 ( .A(n_651), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND5xp2_ASAP7_75t_L g655 ( .A(n_656), .B(n_676), .C(n_689), .D(n_698), .E(n_709), .Y(n_655) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B1(n_668), .B2(n_671), .C(n_673), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B(n_704), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_738), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_SL g756 ( .A(n_735), .B(n_737), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_735), .A2(n_759), .B(n_762), .Y(n_758) );
INVx1_ASAP7_75t_SL g754 ( .A(n_738), .Y(n_754) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx3_ASAP7_75t_L g752 ( .A(n_739), .Y(n_752) );
BUFx2_ASAP7_75t_L g763 ( .A(n_739), .Y(n_763) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_748), .C(n_753), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_742), .A2(n_747), .B(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_749), .B(n_754), .Y(n_753) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
CKINVDCx9p33_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
CKINVDCx11_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
CKINVDCx8_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule