module fake_jpeg_1557_n_241 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_16),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_0),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_1),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_64),
.Y(n_86)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_99),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_18),
.B1(n_25),
.B2(n_22),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_87),
.B1(n_34),
.B2(n_23),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_29),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_61),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_29),
.B1(n_36),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_84),
.B1(n_92),
.B2(n_93),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_29),
.B1(n_36),
.B2(n_25),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_17),
.B1(n_20),
.B2(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_27),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_108),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_30),
.B(n_33),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_121),
.B(n_98),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_110),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_65),
.B1(n_52),
.B2(n_44),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_63),
.B1(n_53),
.B2(n_42),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_129),
.B1(n_75),
.B2(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_96),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_35),
.B(n_59),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_23),
.B1(n_34),
.B2(n_19),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_23),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_70),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_19),
.C(n_3),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_1),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_68),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_154),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_102),
.B1(n_110),
.B2(n_103),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_102),
.B1(n_114),
.B2(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_14),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_66),
.A3(n_88),
.B1(n_83),
.B2(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_83),
.C(n_73),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_119),
.C(n_112),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_116),
.B(n_111),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_95),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_95),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_121),
.B(n_117),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_145),
.B(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_159),
.B(n_175),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_104),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_132),
.B1(n_153),
.B2(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_136),
.B1(n_132),
.B2(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_169),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_119),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_174),
.C(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_146),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_179),
.B1(n_185),
.B2(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_190),
.C(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_151),
.B1(n_144),
.B2(n_135),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_130),
.B(n_142),
.C(n_139),
.D(n_146),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_147),
.A3(n_148),
.B1(n_105),
.B2(n_66),
.C1(n_71),
.C2(n_120),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_175),
.B(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_188),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_71),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_158),
.B1(n_173),
.B2(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_198),
.B1(n_203),
.B2(n_205),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_200),
.C(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_199),
.C(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_156),
.B1(n_148),
.B2(n_138),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_138),
.C(n_109),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_127),
.A3(n_133),
.B1(n_120),
.B2(n_90),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_177),
.C(n_180),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_204),
.Y(n_218)
);

AOI31xp67_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_197),
.A3(n_195),
.B(n_181),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_206),
.A2(n_179),
.B1(n_180),
.B2(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_224),
.B(n_14),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_13),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_220),
.Y(n_230)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_191),
.B(n_189),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_214),
.B(n_211),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_203),
.B(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_215),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_228),
.Y(n_234)
);

OAI221xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_6),
.B1(n_10),
.B2(n_230),
.C(n_228),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_221),
.C(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_10),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_10),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_234),
.B(n_235),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_237),
.C(n_239),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);


endmodule