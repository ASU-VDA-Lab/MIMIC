module fake_jpeg_29047_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_7),
.A2(n_3),
.B1(n_1),
.B2(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx6p67_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_20),
.CI(n_13),
.CON(n_25),
.SN(n_25)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_17),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_16),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_23),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_13),
.B(n_17),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_11),
.C(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_29),
.B(n_25),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_27),
.B(n_25),
.C(n_28),
.Y(n_33)
);


endmodule