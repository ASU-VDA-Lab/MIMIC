module fake_netlist_5_925_n_5259 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_678, n_664, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_5259);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_5259;

wire n_924;
wire n_977;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_882;
wire n_2384;
wire n_3156;
wire n_696;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_870;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1994;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_4294;
wire n_1732;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_727;
wire n_5210;
wire n_4967;
wire n_957;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_4452;
wire n_4348;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_802;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_3178;
wire n_873;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_1726;
wire n_3035;
wire n_5194;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_1109;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_1742;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_3691;
wire n_3628;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1012;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_1061;
wire n_2931;
wire n_5185;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_695;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_951;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_4330;
wire n_3695;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_902;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_858;
wire n_2985;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_705;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_906;
wire n_919;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_2878;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_967;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_2637;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_5173;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_984;
wire n_694;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_849;
wire n_1786;
wire n_4997;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_5243;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_1174;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_3135;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_985;
wire n_3404;
wire n_3217;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_5214;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_4881;
wire n_5089;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_927;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_915;
wire n_864;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_4483;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_897;
wire n_1428;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_857;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_1017;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5216;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_765;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_701;
wire n_1023;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_1060;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_842;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_749;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_4679;
wire n_4115;
wire n_726;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_905;
wire n_5077;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_1028;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_1089;
wire n_5217;
wire n_1004;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_1528;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_1545;
wire n_2374;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_4197;
wire n_4829;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_926;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_1072;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_913;
wire n_3833;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5108;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_750;
wire n_742;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_700;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_764;
wire n_1424;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_1432;
wire n_3875;
wire n_4003;
wire n_2402;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_4682;
wire n_3708;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_1188;
wire n_3957;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_1110;
wire n_3123;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_866;
wire n_5198;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_693;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_710;
wire n_3090;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_737;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_1225;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_699;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_2135;
wire n_3493;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_730;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_2839;
wire n_1588;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_251),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_340),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_556),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_292),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_150),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_687),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_204),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_214),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_179),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_476),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_289),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_56),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_599),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_207),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_98),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_385),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_687),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_647),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_672),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_361),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_312),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_533),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_316),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_416),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_680),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_128),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_334),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_288),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_402),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_130),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_648),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_9),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_394),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_262),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_518),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_109),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_530),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_410),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_533),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_146),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_670),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_275),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_480),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_374),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_544),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_632),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_511),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_388),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_498),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_201),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_610),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_587),
.Y(n_745)
);

BUFx5_ASAP7_75t_L g746 ( 
.A(n_345),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_235),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_127),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_563),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_206),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_47),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_460),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_500),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_389),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_601),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_652),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_202),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_657),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_573),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_222),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_592),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_195),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_206),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_665),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_329),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_378),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_491),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_417),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_137),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_78),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_608),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_139),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_103),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_511),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_330),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_312),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_320),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_243),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_108),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_122),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_371),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_347),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_95),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_106),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_33),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_664),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_418),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_391),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_549),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_23),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_18),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_454),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_178),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_204),
.Y(n_795)
);

CKINVDCx14_ASAP7_75t_R g796 ( 
.A(n_210),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_83),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_101),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_393),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_110),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_452),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_227),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_566),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_256),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_40),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_531),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_584),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_316),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_23),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_273),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_690),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_683),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_240),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_427),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_12),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_256),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_91),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_280),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_137),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_372),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_314),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_175),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_469),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_590),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_153),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_671),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_348),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_181),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_515),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_89),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_609),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_57),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_186),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_461),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_100),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_290),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_323),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_616),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_318),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_570),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_311),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_250),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_415),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_303),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_332),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_231),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_269),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_327),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_90),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_383),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_655),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_666),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_184),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_534),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_330),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_303),
.Y(n_856)
);

BUFx10_ASAP7_75t_L g857 ( 
.A(n_606),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_162),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_667),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_343),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_399),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_406),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_548),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_386),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_482),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_321),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_30),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_649),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_238),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_437),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_635),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_180),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_547),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_54),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_279),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_431),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_566),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_337),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_448),
.Y(n_879)
);

CKINVDCx14_ASAP7_75t_R g880 ( 
.A(n_257),
.Y(n_880)
);

BUFx10_ASAP7_75t_L g881 ( 
.A(n_158),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_506),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_258),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_673),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_227),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_634),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_240),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_81),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_335),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_216),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_198),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_58),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_596),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_30),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_524),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_471),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_444),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_609),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_143),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_596),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_166),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_521),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_170),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_480),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_476),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_23),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_170),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_314),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_669),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_628),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_266),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_195),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_620),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_318),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_254),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_284),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_223),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_214),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_487),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_296),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_570),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_281),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_219),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_2),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_194),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_11),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_337),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_372),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_457),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_123),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_95),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_6),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_4),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_229),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_384),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_433),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_598),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_423),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_654),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_283),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_249),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_460),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_615),
.Y(n_943)
);

BUFx5_ASAP7_75t_L g944 ( 
.A(n_557),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_524),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_53),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_417),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_207),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_628),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_66),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_458),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_611),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_450),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_441),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_354),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_310),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_616),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_203),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_152),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_127),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_517),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_458),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_464),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_264),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_494),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_442),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_329),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_678),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_258),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_248),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_383),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_682),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_565),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_275),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_466),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_644),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_493),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_640),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_76),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_167),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_113),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_287),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_188),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_595),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_247),
.Y(n_985)
);

BUFx8_ASAP7_75t_SL g986 ( 
.A(n_35),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_272),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_600),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_390),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_263),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_232),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_369),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_370),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_157),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_629),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_111),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_210),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_621),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_291),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_246),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_668),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_108),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_428),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_78),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_637),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_646),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_584),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_242),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_64),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_228),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_684),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_469),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_276),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_301),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_652),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_441),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_6),
.Y(n_1017)
);

BUFx8_ASAP7_75t_SL g1018 ( 
.A(n_108),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_470),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_13),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_346),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_613),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_253),
.Y(n_1023)
);

INVxp33_ASAP7_75t_L g1024 ( 
.A(n_57),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_289),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_248),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_447),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_503),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_746),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_746),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_986),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_1018),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_849),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_746),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_796),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_746),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_880),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_746),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_733),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_746),
.Y(n_1040)
);

CKINVDCx14_ASAP7_75t_R g1041 ( 
.A(n_835),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_746),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_839),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_849),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_746),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_736),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_944),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_910),
.B(n_0),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_944),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_944),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_719),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_944),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_944),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_944),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_725),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_725),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_725),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_725),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_725),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_729),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_729),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_759),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_729),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_729),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_729),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_839),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_809),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_824),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_693),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_809),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_809),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_809),
.Y(n_1074)
);

INVxp33_ASAP7_75t_SL g1075 ( 
.A(n_761),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_809),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_817),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_817),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_817),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_719),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_988),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_1005),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_817),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_817),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_760),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_708),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_762),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_1002),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_751),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_770),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_779),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_783),
.Y(n_1092)
);

INVxp33_ASAP7_75t_L g1093 ( 
.A(n_698),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_791),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_797),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_798),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_705),
.B(n_1),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_805),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_766),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_867),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_709),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_768),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_697),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_769),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_771),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_989),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_774),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_775),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1004),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_776),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_839),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1002),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_700),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_839),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_700),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_839),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_723),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_742),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_723),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_742),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_709),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_921),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_777),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_921),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_983),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_912),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_983),
.Y(n_1128)
);

INVxp33_ASAP7_75t_SL g1129 ( 
.A(n_748),
.Y(n_1129)
);

INVxp33_ASAP7_75t_SL g1130 ( 
.A(n_748),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_912),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_773),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_912),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_912),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_912),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_784),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_960),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_792),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_927),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_927),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_927),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_927),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_815),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_717),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_781),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_927),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_965),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_965),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_965),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_782),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_965),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_787),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1024),
.B(n_800),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_965),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_785),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_709),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_789),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_794),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_960),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_785),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_926),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_786),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_926),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_830),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_874),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_979),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_888),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_894),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_906),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_699),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_924),
.Y(n_1171)
);

CKINVDCx16_ASAP7_75t_R g1172 ( 
.A(n_786),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_795),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_780),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_701),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_801),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_715),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_979),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_715),
.Y(n_1179)
);

INVxp33_ASAP7_75t_L g1180 ( 
.A(n_706),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_767),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_707),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_802),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_804),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_711),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_714),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_807),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_810),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_724),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_752),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_812),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_813),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_726),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_754),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_767),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_816),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_755),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_818),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_981),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_819),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_820),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_823),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_786),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_756),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_763),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_764),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_765),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_823),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_778),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_790),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_981),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_829),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_793),
.Y(n_1213)
);

BUFx5_ASAP7_75t_L g1214 ( 
.A(n_803),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_832),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_892),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_799),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_806),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_808),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1009),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_753),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_821),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_828),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_758),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_831),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_814),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_833),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_825),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_788),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_829),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_SL g1231 ( 
.A(n_799),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_836),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_826),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_827),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_844),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_811),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_840),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_852),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_837),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_854),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_838),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_856),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_864),
.Y(n_1243)
);

CKINVDCx16_ASAP7_75t_R g1244 ( 
.A(n_799),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_822),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_822),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_868),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1009),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_869),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_872),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_841),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_843),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_875),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_845),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_879),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_883),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_851),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_853),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_834),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_885),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_842),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_886),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_822),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_855),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_840),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_887),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_895),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_847),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_898),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_846),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_905),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_914),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_857),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_847),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_857),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_915),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_919),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_858),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_934),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_859),
.Y(n_1280)
);

CKINVDCx14_ASAP7_75t_R g1281 ( 
.A(n_857),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_936),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_862),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_848),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_939),
.Y(n_1285)
);

CKINVDCx14_ASAP7_75t_R g1286 ( 
.A(n_862),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_863),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_866),
.Y(n_1288)
);

CKINVDCx16_ASAP7_75t_R g1289 ( 
.A(n_862),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_911),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_949),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_881),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_954),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_881),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_860),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_961),
.Y(n_1296)
);

INVxp33_ASAP7_75t_L g1297 ( 
.A(n_962),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_865),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_964),
.Y(n_1299)
);

CKINVDCx16_ASAP7_75t_R g1300 ( 
.A(n_881),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_967),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_873),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_876),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_971),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_878),
.Y(n_1305)
);

INVxp33_ASAP7_75t_L g1306 ( 
.A(n_973),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_882),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_884),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_890),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_999),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_975),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_976),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_891),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_991),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_995),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_997),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1006),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1008),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_893),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1010),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_877),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1022),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_899),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1026),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_903),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_896),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_913),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1027),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_897),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_848),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_900),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_850),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_850),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_889),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_889),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_902),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_901),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_901),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_922),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_904),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_922),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_951),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_951),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_980),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_978),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_978),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_907),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_984),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_908),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_984),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_999),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_909),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_999),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_800),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_712),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_712),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_870),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_916),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_1017),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_870),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1007),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_1014),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1007),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_917),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_772),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_918),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_930),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_920),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_923),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_925),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_928),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_929),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1017),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_931),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_935),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_932),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_938),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_940),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_941),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_943),
.Y(n_1380)
);

CKINVDCx14_ASAP7_75t_R g1381 ( 
.A(n_933),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_945),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_947),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_948),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_952),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_946),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_953),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_955),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1020),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_713),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_956),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_957),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_958),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1057),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1071),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1058),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1035),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1059),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1071),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1035),
.B(n_950),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1037),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1060),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1061),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1063),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1390),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1132),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1136),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1039),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1062),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1065),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1375),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1066),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1364),
.B(n_1028),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1067),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1366),
.B(n_1020),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1103),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1069),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1072),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1037),
.B(n_694),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1103),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1138),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1073),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1074),
.Y(n_1423)
);

CKINVDCx14_ASAP7_75t_R g1424 ( 
.A(n_1281),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_694),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1144),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1144),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1193),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1077),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1143),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1078),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1079),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1083),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1084),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1164),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1131),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1165),
.Y(n_1437)
);

INVxp67_ASAP7_75t_SL g1438 ( 
.A(n_1375),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1193),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1134),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1135),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_L g1442 ( 
.A(n_1364),
.B(n_0),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1139),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1140),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1142),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1031),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1149),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1151),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1063),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_R g1450 ( 
.A(n_1381),
.B(n_695),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1221),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1221),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1224),
.Y(n_1453)
);

INVxp33_ASAP7_75t_SL g1454 ( 
.A(n_1032),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1076),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1167),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1168),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1051),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1076),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1169),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1043),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1224),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1148),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1148),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1117),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1112),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1112),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1115),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_R g1469 ( 
.A(n_1171),
.B(n_695),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1375),
.B(n_1364),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1236),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1115),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1085),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1085),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1127),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1236),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1127),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1259),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1087),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1133),
.Y(n_1480)
);

INVxp33_ASAP7_75t_SL g1481 ( 
.A(n_1032),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1087),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_L g1483 ( 
.A(n_1099),
.B(n_1102),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1375),
.B(n_696),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1133),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1141),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1099),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1141),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1102),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1147),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1039),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1105),
.B(n_696),
.Y(n_1492)
);

CKINVDCx16_ASAP7_75t_R g1493 ( 
.A(n_1362),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1118),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1105),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1385),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1106),
.B(n_0),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1106),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1147),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1154),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1108),
.B(n_702),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1120),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1108),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1259),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1107),
.B(n_716),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1154),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1117),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1043),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1117),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1113),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1354),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1109),
.B(n_702),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1044),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1109),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1111),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_1111),
.B(n_1),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1043),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1124),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1170),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1385),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1175),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1295),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1182),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1185),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1186),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1189),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_R g1527 ( 
.A(n_1124),
.B(n_703),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1190),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1368),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1145),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1145),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1295),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1150),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1194),
.Y(n_1534)
);

CKINVDCx16_ASAP7_75t_R g1535 ( 
.A(n_1286),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1150),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_L g1537 ( 
.A(n_1152),
.B(n_1),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1152),
.B(n_703),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1046),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1197),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1204),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1205),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1157),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1298),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1374),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1298),
.Y(n_1546)
);

INVxp33_ASAP7_75t_SL g1547 ( 
.A(n_1046),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1157),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1206),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1044),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1369),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1302),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1064),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1207),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1209),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1158),
.B(n_704),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1158),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1210),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1173),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1213),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1218),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1302),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1173),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1219),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1064),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1226),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1228),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1070),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1159),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1043),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1176),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1176),
.B(n_704),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1183),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1183),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1184),
.B(n_710),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1184),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1374),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1043),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1321),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1068),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1233),
.Y(n_1581)
);

INVxp33_ASAP7_75t_L g1582 ( 
.A(n_1178),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1321),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1234),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1235),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1229),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1187),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1101),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1238),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1240),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1187),
.B(n_2),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1242),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1323),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1323),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1325),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1243),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1068),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1247),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1249),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1250),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1068),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1188),
.Y(n_1602)
);

CKINVDCx16_ASAP7_75t_R g1603 ( 
.A(n_1172),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1253),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1325),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1070),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1255),
.Y(n_1607)
);

INVxp33_ASAP7_75t_SL g1608 ( 
.A(n_1081),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_1244),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1256),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1260),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1262),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1188),
.B(n_1191),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1191),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1211),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1192),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1266),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1081),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1327),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1327),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1192),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1267),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1269),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1344),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1196),
.B(n_710),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1370),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1271),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1371),
.B(n_718),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1068),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1272),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1276),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1248),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1196),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1277),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1198),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1279),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1282),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1068),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1198),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1344),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1386),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_1386),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1285),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1291),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1200),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1293),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1296),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1299),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1372),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1080),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1301),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1246),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1200),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1304),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1311),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1137),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1166),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1201),
.Y(n_1658)
);

INVxp33_ASAP7_75t_SL g1659 ( 
.A(n_1082),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1312),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1314),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1263),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1201),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1283),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1222),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1289),
.Y(n_1666)
);

CKINVDCx16_ASAP7_75t_R g1667 ( 
.A(n_1294),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1300),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1222),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1315),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1082),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1316),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1378),
.B(n_1379),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1223),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1317),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1223),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1318),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1320),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1322),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1261),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1225),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1324),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1225),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1227),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1227),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1328),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1232),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1270),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_1174),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1232),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1116),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1382),
.B(n_718),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1239),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1215),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_1216),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1239),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1119),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1123),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1241),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1461),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1510),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1404),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1404),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1466),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1470),
.B(n_1367),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1463),
.B(n_1177),
.Y(n_1706)
);

INVx5_ASAP7_75t_L g1707 ( 
.A(n_1461),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1461),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1461),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1689),
.A2(n_1695),
.B1(n_1694),
.B2(n_1680),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1464),
.B(n_1177),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1467),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1691),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1442),
.B(n_1179),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1697),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1638),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1586),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1411),
.B(n_1367),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1638),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1638),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1438),
.B(n_1179),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1698),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1513),
.B(n_1181),
.Y(n_1723)
);

NAND2xp33_ASAP7_75t_L g1724 ( 
.A(n_1673),
.B(n_1214),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1468),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1529),
.B(n_1387),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1505),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1472),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1638),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1519),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1475),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1405),
.B(n_1129),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1551),
.B(n_1388),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1626),
.B(n_1391),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1649),
.B(n_1129),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1469),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1513),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1477),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1521),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1550),
.B(n_1181),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1436),
.A2(n_1030),
.B(n_1029),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1492),
.A2(n_1075),
.B1(n_1251),
.B2(n_1241),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1601),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1689),
.A2(n_1130),
.B1(n_1075),
.B2(n_1041),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1480),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1485),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1601),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1415),
.A2(n_1130),
.B1(n_1376),
.B2(n_1252),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1523),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1486),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1601),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1524),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1425),
.B(n_1484),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1508),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1488),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1424),
.B(n_1376),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1490),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_R g1758 ( 
.A(n_1527),
.B(n_1665),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1413),
.B(n_1251),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1694),
.A2(n_721),
.B1(n_722),
.B2(n_720),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1499),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1695),
.A2(n_1680),
.B1(n_1688),
.B2(n_1671),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1500),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1525),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1550),
.B(n_1195),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1506),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1508),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1449),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1496),
.B(n_1195),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1526),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1520),
.B(n_1392),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1517),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1517),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1582),
.B(n_1156),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1528),
.B(n_1230),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1465),
.Y(n_1776)
);

NOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1465),
.B(n_1393),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1509),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1628),
.A2(n_1049),
.B(n_1036),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1534),
.B(n_1230),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1501),
.B(n_1156),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1455),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1540),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1570),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1459),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1541),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1570),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1542),
.B(n_1549),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1578),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1554),
.B(n_1268),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1509),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1555),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1578),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1580),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1688),
.A2(n_721),
.B1(n_722),
.B2(n_720),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1558),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1560),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1561),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1512),
.B(n_1275),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1580),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1597),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1564),
.B(n_1268),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1566),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1538),
.B(n_1556),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1567),
.B(n_1274),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1507),
.B(n_1034),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1581),
.B(n_1274),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1584),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1419),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1597),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1585),
.B(n_1335),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1629),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1629),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1572),
.B(n_1275),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1440),
.Y(n_1815)
);

OA21x2_ASAP7_75t_L g1816 ( 
.A1(n_1441),
.A2(n_1040),
.B(n_1038),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1394),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1443),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1589),
.B(n_1335),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1396),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1398),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1402),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1403),
.B(n_1042),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1590),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1483),
.B(n_1114),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_1395),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1575),
.B(n_1252),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1592),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1450),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1535),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1625),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1692),
.A2(n_1049),
.B(n_1036),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1409),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1444),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1458),
.B(n_1254),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1410),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1493),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1494),
.B(n_1254),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1596),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1412),
.B(n_1045),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1414),
.B(n_1047),
.Y(n_1841)
);

INVx5_ASAP7_75t_L g1842 ( 
.A(n_1445),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1417),
.B(n_1050),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1418),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1422),
.B(n_1054),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1598),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1447),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1613),
.A2(n_1257),
.B1(n_1264),
.B2(n_1258),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1423),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1429),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1671),
.A2(n_1093),
.B1(n_728),
.B2(n_730),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1652),
.A2(n_728),
.B1(n_730),
.B2(n_727),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1431),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1502),
.B(n_1257),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1448),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1432),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1599),
.B(n_1160),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1397),
.Y(n_1858)
);

CKINVDCx11_ASAP7_75t_R g1859 ( 
.A(n_1395),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1569),
.A2(n_1264),
.B1(n_1278),
.B2(n_1258),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1600),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1433),
.Y(n_1862)
);

OAI21x1_ASAP7_75t_L g1863 ( 
.A1(n_1434),
.A2(n_1053),
.B(n_1052),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1604),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1607),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1400),
.A2(n_1278),
.B1(n_1287),
.B2(n_1280),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1610),
.Y(n_1867)
);

AND2x6_ASAP7_75t_L g1868 ( 
.A(n_1611),
.B(n_1055),
.Y(n_1868)
);

BUFx8_ASAP7_75t_L g1869 ( 
.A(n_1545),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1612),
.B(n_1160),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1617),
.B(n_1088),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1615),
.B(n_1280),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1622),
.B(n_1056),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1623),
.B(n_1088),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1627),
.B(n_1033),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1630),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1631),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1634),
.B(n_1636),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1637),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1643),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1644),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1632),
.B(n_1287),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1646),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1650),
.B(n_1288),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1647),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1648),
.A2(n_1053),
.B(n_1052),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1651),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1654),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1656),
.B(n_1288),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1657),
.B(n_1303),
.Y(n_1890)
);

CKINVDCx6p67_ASAP7_75t_R g1891 ( 
.A(n_1588),
.Y(n_1891)
);

OA21x2_ASAP7_75t_L g1892 ( 
.A1(n_1655),
.A2(n_1365),
.B(n_1126),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1660),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1547),
.A2(n_1305),
.B1(n_1307),
.B2(n_1303),
.Y(n_1894)
);

CKINVDCx14_ASAP7_75t_R g1895 ( 
.A(n_1652),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1661),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1670),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1672),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1497),
.A2(n_1307),
.B1(n_1308),
.B2(n_1305),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1675),
.Y(n_1900)
);

AND2x6_ASAP7_75t_L g1901 ( 
.A(n_1677),
.B(n_1153),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1678),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1679),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1516),
.A2(n_1309),
.B1(n_1313),
.B2(n_1308),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1682),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1547),
.A2(n_1309),
.B1(n_1319),
.B2(n_1313),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1686),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1608),
.A2(n_1319),
.B1(n_1329),
.B2(n_1326),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1511),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1406),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1407),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1537),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1591),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1397),
.A2(n_1329),
.B1(n_1331),
.B2(n_1326),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1421),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1681),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1684),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1687),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1430),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1408),
.B(n_1033),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1491),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1435),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1437),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1608),
.A2(n_1331),
.B1(n_1340),
.B2(n_1336),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1401),
.A2(n_1340),
.B1(n_1347),
.B2(n_1336),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1539),
.A2(n_1342),
.B(n_1212),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1456),
.B(n_1347),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1457),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1553),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1659),
.A2(n_1349),
.B1(n_1358),
.B2(n_1352),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1565),
.B(n_1086),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1568),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1456),
.B(n_1349),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1606),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_SL g1935 ( 
.A1(n_1662),
.A2(n_731),
.B1(n_732),
.B2(n_727),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1460),
.B(n_1352),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1473),
.B(n_1358),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1474),
.B(n_1377),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1618),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1479),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1482),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1487),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1489),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1495),
.B(n_1089),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1498),
.B(n_1146),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1401),
.A2(n_1380),
.B1(n_1383),
.B2(n_1377),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1503),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1514),
.B(n_1380),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1515),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1518),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1530),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1531),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1533),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1536),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1543),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1548),
.B(n_1090),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1557),
.B(n_1091),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1559),
.B(n_1146),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1563),
.B(n_1146),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1571),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1573),
.Y(n_1961)
);

INVx5_ASAP7_75t_L g1962 ( 
.A(n_1603),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1659),
.A2(n_1383),
.B1(n_1384),
.B2(n_1290),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1574),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1576),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1587),
.B(n_1384),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1602),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1454),
.B(n_1231),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1614),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1616),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1621),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1633),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1635),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1639),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1645),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1653),
.Y(n_1976)
);

AND2x6_ASAP7_75t_L g1977 ( 
.A(n_1454),
.B(n_1203),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1658),
.A2(n_1389),
.B1(n_1220),
.B2(n_1199),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1663),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1665),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1669),
.B(n_1092),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1669),
.A2(n_1122),
.B1(n_1310),
.B2(n_1162),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1662),
.A2(n_732),
.B1(n_734),
.B2(n_731),
.Y(n_1983)
);

OA21x2_ASAP7_75t_L g1984 ( 
.A1(n_1699),
.A2(n_1128),
.B(n_1125),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1674),
.B(n_1146),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1674),
.B(n_1203),
.Y(n_1986)
);

AND2x6_ASAP7_75t_L g1987 ( 
.A(n_1481),
.B(n_1217),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1577),
.Y(n_1988)
);

BUFx10_ASAP7_75t_L g1989 ( 
.A(n_1936),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1753),
.A2(n_1683),
.B1(n_1685),
.B2(n_1676),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1717),
.B(n_1676),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1831),
.B(n_1683),
.Y(n_1992)
);

OAI22xp33_ASAP7_75t_R g1993 ( 
.A1(n_1735),
.A2(n_1097),
.B1(n_942),
.B2(n_871),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_SL g1994 ( 
.A1(n_1759),
.A2(n_1690),
.B1(n_1693),
.B2(n_1685),
.Y(n_1994)
);

AO22x1_ASAP7_75t_L g1995 ( 
.A1(n_1804),
.A2(n_1693),
.B1(n_1696),
.B2(n_1690),
.Y(n_1995)
);

AO22x2_ASAP7_75t_L g1996 ( 
.A1(n_1860),
.A2(n_1748),
.B1(n_1809),
.B2(n_1914),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1705),
.A2(n_1736),
.B1(n_1733),
.B2(n_1734),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1702),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1886),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1732),
.B(n_1696),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1726),
.A2(n_1699),
.B1(n_1609),
.B2(n_1667),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1762),
.A2(n_1642),
.B1(n_1641),
.B2(n_1416),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1702),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1718),
.B(n_1214),
.Y(n_2004)
);

NAND3x1_ASAP7_75t_L g2005 ( 
.A(n_1894),
.B(n_1353),
.C(n_1351),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1781),
.B(n_1664),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1759),
.A2(n_735),
.B1(n_737),
.B2(n_734),
.Y(n_2007)
);

AO22x2_ASAP7_75t_L g2008 ( 
.A1(n_1925),
.A2(n_937),
.B1(n_1012),
.B2(n_741),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1901),
.A2(n_1446),
.B1(n_1481),
.B2(n_1214),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1703),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1901),
.A2(n_1446),
.B1(n_1214),
.B2(n_1048),
.Y(n_2011)
);

OAI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1735),
.A2(n_1025),
.B1(n_737),
.B2(n_738),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1703),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1717),
.B(n_1217),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1771),
.A2(n_1297),
.B1(n_1306),
.B2(n_1180),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1901),
.A2(n_1214),
.B1(n_1668),
.B2(n_1666),
.Y(n_2016)
);

OR2x6_ASAP7_75t_L g2017 ( 
.A(n_1911),
.B(n_1121),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1912),
.A2(n_1273),
.B1(n_1292),
.B2(n_1245),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1704),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1737),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1727),
.B(n_1359),
.Y(n_2021)
);

OA22x2_ASAP7_75t_L g2022 ( 
.A1(n_1760),
.A2(n_738),
.B1(n_970),
.B2(n_750),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1886),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1769),
.B(n_1214),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1769),
.B(n_1721),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1901),
.A2(n_1214),
.B1(n_1668),
.B2(n_1666),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1886),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1901),
.A2(n_1208),
.B1(n_1237),
.B2(n_1202),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1863),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1863),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1913),
.A2(n_1273),
.B1(n_1292),
.B2(n_1245),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1704),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1727),
.B(n_1359),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1774),
.B(n_1359),
.Y(n_2034)
);

OA22x2_ASAP7_75t_L g2035 ( 
.A1(n_1795),
.A2(n_739),
.B1(n_972),
.B2(n_757),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1732),
.A2(n_1208),
.B1(n_1237),
.B2(n_1202),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_SL g2037 ( 
.A1(n_1985),
.A2(n_739),
.B1(n_740),
.B2(n_735),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1799),
.A2(n_743),
.B1(n_744),
.B2(n_740),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1814),
.B(n_1373),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1866),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_SL g2041 ( 
.A1(n_1895),
.A2(n_1641),
.B1(n_1642),
.B2(n_1416),
.Y(n_2041)
);

OAI22xp33_ASAP7_75t_SL g2042 ( 
.A1(n_1730),
.A2(n_747),
.B1(n_749),
.B2(n_745),
.Y(n_2042)
);

OA22x2_ASAP7_75t_L g2043 ( 
.A1(n_1742),
.A2(n_749),
.B1(n_990),
.B2(n_969),
.Y(n_2043)
);

AO22x2_ASAP7_75t_L g2044 ( 
.A1(n_1946),
.A2(n_1121),
.B1(n_1356),
.B2(n_1355),
.Y(n_2044)
);

OAI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1806),
.A2(n_750),
.B1(n_757),
.B2(n_747),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1984),
.A2(n_1208),
.B1(n_1237),
.B2(n_1202),
.Y(n_2046)
);

AO22x2_ASAP7_75t_L g2047 ( 
.A1(n_1980),
.A2(n_1357),
.B1(n_1361),
.B2(n_1360),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_1984),
.A2(n_1208),
.B1(n_1237),
.B2(n_1202),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1848),
.A2(n_959),
.B1(n_963),
.B2(n_861),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_R g2050 ( 
.A1(n_1854),
.A2(n_1095),
.B1(n_1096),
.B2(n_1094),
.Y(n_2050)
);

INVx8_ASAP7_75t_L g2051 ( 
.A(n_1962),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1920),
.B(n_1373),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1712),
.Y(n_2053)
);

OAI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1902),
.A2(n_959),
.B1(n_963),
.B2(n_861),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1712),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1725),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1725),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1728),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1827),
.A2(n_968),
.B1(n_969),
.B2(n_966),
.Y(n_2059)
);

AO22x2_ASAP7_75t_L g2060 ( 
.A1(n_1899),
.A2(n_1363),
.B1(n_1114),
.B2(n_1100),
.Y(n_2060)
);

AO22x2_ASAP7_75t_L g2061 ( 
.A1(n_1904),
.A2(n_1104),
.B1(n_1110),
.B2(n_1098),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1984),
.A2(n_1208),
.B1(n_1237),
.B2(n_1202),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1728),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1920),
.B(n_1373),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1920),
.B(n_1155),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1854),
.B(n_1399),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1835),
.B(n_1161),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1981),
.A2(n_968),
.B1(n_970),
.B2(n_966),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1731),
.Y(n_2069)
);

AO22x2_ASAP7_75t_L g2070 ( 
.A1(n_1916),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1769),
.A2(n_1981),
.B1(n_1724),
.B2(n_1872),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1902),
.A2(n_1903),
.B1(n_1978),
.B2(n_1982),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1931),
.B(n_972),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_SL g2074 ( 
.A(n_1939),
.B(n_974),
.Y(n_2074)
);

AOI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1981),
.A2(n_1265),
.B1(n_1284),
.B2(n_1330),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1838),
.B(n_1163),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1721),
.B(n_1265),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1882),
.B(n_1332),
.Y(n_2078)
);

AND2x6_ASAP7_75t_L g2079 ( 
.A(n_1756),
.B(n_1333),
.Y(n_2079)
);

OAI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1903),
.A2(n_977),
.B1(n_982),
.B2(n_974),
.Y(n_2080)
);

OAI22xp33_ASAP7_75t_SL g2081 ( 
.A1(n_1739),
.A2(n_982),
.B1(n_985),
.B2(n_977),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1884),
.B(n_1334),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1737),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_SL g2084 ( 
.A1(n_1749),
.A2(n_987),
.B1(n_990),
.B2(n_985),
.Y(n_2084)
);

AND2x2_ASAP7_75t_SL g2085 ( 
.A(n_1927),
.B(n_1933),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1724),
.A2(n_1284),
.B1(n_1265),
.B2(n_1337),
.Y(n_2086)
);

AO22x2_ASAP7_75t_L g2087 ( 
.A1(n_1916),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1731),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1889),
.B(n_1338),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_SL g2090 ( 
.A1(n_1752),
.A2(n_1770),
.B1(n_1783),
.B2(n_1764),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1738),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1738),
.Y(n_2092)
);

OAI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1786),
.A2(n_1796),
.B1(n_1797),
.B2(n_1792),
.Y(n_2093)
);

AOI22x1_ASAP7_75t_SL g2094 ( 
.A1(n_1826),
.A2(n_1420),
.B1(n_1426),
.B2(n_1399),
.Y(n_2094)
);

OAI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1963),
.A2(n_992),
.B1(n_993),
.B2(n_987),
.Y(n_2095)
);

INVx8_ASAP7_75t_L g2096 ( 
.A(n_1962),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1890),
.B(n_1339),
.Y(n_2097)
);

OAI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1865),
.A2(n_993),
.B1(n_994),
.B2(n_992),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1745),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_1871),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1745),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1909),
.Y(n_2102)
);

AO22x2_ASAP7_75t_L g2103 ( 
.A1(n_1917),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_2103)
);

AO22x2_ASAP7_75t_L g2104 ( 
.A1(n_1918),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_2104)
);

NAND3x1_ASAP7_75t_L g2105 ( 
.A(n_1906),
.B(n_1343),
.C(n_1341),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1746),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_1826),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1865),
.A2(n_998),
.B1(n_1000),
.B2(n_994),
.Y(n_2108)
);

NAND3x1_ASAP7_75t_L g2109 ( 
.A(n_1908),
.B(n_1346),
.C(n_1345),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1721),
.B(n_1265),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1909),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1706),
.Y(n_2112)
);

XNOR2xp5_ASAP7_75t_L g2113 ( 
.A(n_1837),
.B(n_1420),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_1706),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1746),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1750),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1872),
.A2(n_1284),
.B1(n_1265),
.B2(n_1348),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1944),
.B(n_1350),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_SL g2119 ( 
.A1(n_1895),
.A2(n_1427),
.B1(n_1428),
.B2(n_1426),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1944),
.B(n_1212),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1944),
.B(n_1212),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1750),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1956),
.B(n_1342),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1956),
.B(n_1342),
.Y(n_2124)
);

OAI22xp33_ASAP7_75t_SL g2125 ( 
.A1(n_1798),
.A2(n_1000),
.B1(n_1001),
.B2(n_998),
.Y(n_2125)
);

OAI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_1867),
.A2(n_1003),
.B1(n_1011),
.B2(n_1001),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1956),
.B(n_1003),
.Y(n_2127)
);

OAI22xp33_ASAP7_75t_SL g2128 ( 
.A1(n_1803),
.A2(n_1013),
.B1(n_1015),
.B2(n_1011),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1755),
.Y(n_2129)
);

OAI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_1867),
.A2(n_1015),
.B1(n_1016),
.B2(n_1013),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1755),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_1957),
.A2(n_1284),
.B1(n_1019),
.B2(n_1021),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1757),
.Y(n_2133)
);

OA22x2_ASAP7_75t_L g2134 ( 
.A1(n_1852),
.A2(n_1019),
.B1(n_1021),
.B2(n_1016),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1957),
.B(n_1023),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1957),
.A2(n_1284),
.B1(n_1023),
.B2(n_1146),
.Y(n_2136)
);

OAI22xp33_ASAP7_75t_SL g2137 ( 
.A1(n_1808),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1788),
.A2(n_1428),
.B1(n_1439),
.B2(n_1427),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1706),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_1988),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1892),
.A2(n_1451),
.B1(n_1452),
.B2(n_1439),
.Y(n_2141)
);

OAI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_1876),
.A2(n_1452),
.B1(n_1453),
.B2(n_1451),
.Y(n_2142)
);

OR2x6_ASAP7_75t_L g2143 ( 
.A(n_1911),
.B(n_1453),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1788),
.A2(n_1471),
.B1(n_1476),
.B2(n_1462),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1757),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1761),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1761),
.Y(n_2147)
);

AO22x2_ASAP7_75t_L g2148 ( 
.A1(n_1940),
.A2(n_1941),
.B1(n_1951),
.B2(n_1942),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_1711),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1763),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1939),
.B(n_1938),
.Y(n_2151)
);

AO22x2_ASAP7_75t_L g2152 ( 
.A1(n_1952),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2152)
);

AO22x2_ASAP7_75t_L g2153 ( 
.A1(n_1953),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1788),
.A2(n_1471),
.B1(n_1476),
.B2(n_1462),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1763),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_1878),
.A2(n_1504),
.B1(n_1522),
.B2(n_1478),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1766),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_1878),
.A2(n_1504),
.B1(n_1522),
.B2(n_1478),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1766),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1711),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1986),
.B(n_1532),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1768),
.Y(n_2162)
);

OA22x2_ASAP7_75t_L g2163 ( 
.A1(n_1935),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1966),
.B(n_1552),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1931),
.B(n_1552),
.Y(n_2165)
);

AO22x2_ASAP7_75t_L g2166 ( 
.A1(n_1955),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1878),
.A2(n_1544),
.B1(n_1546),
.B2(n_1532),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_1710),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1768),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1931),
.B(n_1583),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_1876),
.A2(n_1546),
.B1(n_1562),
.B2(n_1544),
.Y(n_2171)
);

OR2x6_ASAP7_75t_L g2172 ( 
.A(n_1911),
.B(n_1562),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1711),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1723),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1782),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1782),
.Y(n_2176)
);

OAI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_1824),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2177)
);

BUFx10_ASAP7_75t_L g2178 ( 
.A(n_1936),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1892),
.A2(n_1583),
.B1(n_1593),
.B2(n_1579),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1986),
.B(n_1619),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1785),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1785),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1875),
.B(n_1619),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1787),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_1937),
.B(n_1579),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_1937),
.B(n_1593),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1787),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1820),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1875),
.B(n_1640),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1820),
.Y(n_2190)
);

OAI22xp33_ASAP7_75t_SL g2191 ( 
.A1(n_1828),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1948),
.B(n_1594),
.Y(n_2192)
);

OAI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_1877),
.A2(n_1595),
.B1(n_1605),
.B2(n_1594),
.Y(n_2193)
);

OAI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_1877),
.A2(n_1605),
.B1(n_1620),
.B2(n_1595),
.Y(n_2194)
);

OAI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_1880),
.A2(n_1893),
.B1(n_1896),
.B2(n_1887),
.Y(n_2195)
);

OAI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_1880),
.A2(n_1624),
.B1(n_1640),
.B2(n_1620),
.Y(n_2196)
);

AO22x2_ASAP7_75t_L g2197 ( 
.A1(n_1967),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1875),
.B(n_1624),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_1871),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1839),
.A2(n_138),
.B1(n_139),
.B2(n_136),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1821),
.Y(n_2201)
);

OR2x6_ASAP7_75t_L g2202 ( 
.A(n_1911),
.B(n_16),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1964),
.B(n_685),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1909),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1821),
.Y(n_2205)
);

AO22x2_ASAP7_75t_L g2206 ( 
.A1(n_1969),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1846),
.A2(n_138),
.B1(n_140),
.B2(n_136),
.Y(n_2207)
);

INVx8_ASAP7_75t_L g2208 ( 
.A(n_1962),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1861),
.A2(n_141),
.B1(n_142),
.B2(n_140),
.Y(n_2209)
);

OA22x2_ASAP7_75t_L g2210 ( 
.A1(n_1983),
.A2(n_1924),
.B1(n_1930),
.B2(n_1744),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_1723),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1864),
.A2(n_142),
.B1(n_143),
.B2(n_141),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_1879),
.A2(n_145),
.B1(n_146),
.B2(n_144),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1964),
.B(n_144),
.Y(n_2214)
);

OAI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_1887),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1822),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1892),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1948),
.B(n_680),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1723),
.B(n_681),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1822),
.Y(n_2220)
);

BUFx10_ASAP7_75t_L g2221 ( 
.A(n_1829),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_1881),
.A2(n_147),
.B1(n_148),
.B2(n_145),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1800),
.Y(n_2223)
);

OAI22xp33_ASAP7_75t_SL g2224 ( 
.A1(n_1885),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1833),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_SL g2226 ( 
.A1(n_1858),
.A2(n_29),
.B1(n_37),
.B2(n_20),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1897),
.A2(n_148),
.B1(n_149),
.B2(n_147),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_1900),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_2228)
);

AO22x2_ASAP7_75t_L g2229 ( 
.A1(n_1972),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1740),
.B(n_689),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1740),
.B(n_689),
.Y(n_2231)
);

BUFx10_ASAP7_75t_L g2232 ( 
.A(n_1829),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1800),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_1945),
.B(n_22),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1813),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1909),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_1701),
.A2(n_152),
.B1(n_153),
.B2(n_151),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1740),
.B(n_675),
.Y(n_2238)
);

OAI22xp33_ASAP7_75t_SL g2239 ( 
.A1(n_1958),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1833),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1959),
.B(n_24),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1713),
.A2(n_155),
.B1(n_156),
.B2(n_154),
.Y(n_2242)
);

OAI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1893),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2243)
);

INVxp33_ASAP7_75t_L g2244 ( 
.A(n_1851),
.Y(n_2244)
);

AO22x2_ASAP7_75t_L g2245 ( 
.A1(n_1973),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1921),
.B(n_27),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_1765),
.B(n_679),
.Y(n_2247)
);

OA22x2_ASAP7_75t_L g2248 ( 
.A1(n_1929),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1776),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_2249)
);

AOI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_1715),
.A2(n_155),
.B1(n_156),
.B2(n_154),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1722),
.A2(n_158),
.B1(n_159),
.B2(n_157),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_SL g2252 ( 
.A1(n_1858),
.A2(n_38),
.B1(n_46),
.B2(n_28),
.Y(n_2252)
);

AO22x2_ASAP7_75t_L g2253 ( 
.A1(n_1949),
.A2(n_1954),
.B1(n_1950),
.B2(n_1965),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1844),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1765),
.B(n_690),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_1776),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2256)
);

OAI22xp33_ASAP7_75t_SL g2257 ( 
.A1(n_1932),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1765),
.B(n_159),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_1977),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_2259)
);

OAI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_1896),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1947),
.B(n_676),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_1977),
.A2(n_1987),
.B1(n_1868),
.B2(n_1714),
.Y(n_2262)
);

OAI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_1898),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2263)
);

AO22x2_ASAP7_75t_L g2264 ( 
.A1(n_1949),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_1947),
.B(n_678),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_1977),
.A2(n_161),
.B1(n_163),
.B2(n_160),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1714),
.B(n_36),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_SL g2268 ( 
.A1(n_1934),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2268)
);

AO22x2_ASAP7_75t_L g2269 ( 
.A1(n_1950),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2269)
);

OR2x6_ASAP7_75t_L g2270 ( 
.A(n_1919),
.B(n_39),
.Y(n_2270)
);

OAI22xp33_ASAP7_75t_SL g2271 ( 
.A1(n_1898),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_1977),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_2272)
);

OAI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_1905),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1813),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1922),
.B(n_1923),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_1954),
.B(n_691),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1977),
.A2(n_165),
.B1(n_166),
.B2(n_164),
.Y(n_2277)
);

BUFx10_ASAP7_75t_L g2278 ( 
.A(n_1830),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_1965),
.B(n_674),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1844),
.Y(n_2280)
);

AO22x2_ASAP7_75t_L g2281 ( 
.A1(n_1970),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2281)
);

AOI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_1987),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1970),
.B(n_676),
.Y(n_2283)
);

AO22x2_ASAP7_75t_L g2284 ( 
.A1(n_1975),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1714),
.B(n_44),
.Y(n_2285)
);

OAI22xp33_ASAP7_75t_SL g2286 ( 
.A1(n_1905),
.A2(n_1907),
.B1(n_1976),
.B2(n_1975),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_1987),
.A2(n_169),
.B1(n_171),
.B2(n_168),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1817),
.B(n_44),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_1922),
.B(n_1923),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_1987),
.A2(n_172),
.B1(n_173),
.B2(n_171),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1741),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_1775),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1849),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1976),
.B(n_684),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1849),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1850),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_SL g2297 ( 
.A1(n_1907),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1943),
.B(n_691),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_1775),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_1859),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_1883),
.B(n_48),
.Y(n_2301)
);

AO22x2_ASAP7_75t_L g2302 ( 
.A1(n_1910),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1857),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1741),
.Y(n_2304)
);

AOI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_1987),
.A2(n_173),
.B1(n_174),
.B2(n_172),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_1883),
.A2(n_1888),
.B1(n_1758),
.B2(n_1968),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_1868),
.A2(n_175),
.B1(n_176),
.B2(n_174),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1868),
.A2(n_177),
.B1(n_178),
.B2(n_176),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1741),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2218),
.A2(n_1868),
.B1(n_1888),
.B2(n_1883),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2174),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2100),
.B(n_1778),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2174),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_2014),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_2211),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1997),
.B(n_1817),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2306),
.B(n_1919),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2184),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2184),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2071),
.B(n_2286),
.Y(n_2320)
);

AND2x6_ASAP7_75t_L g2321 ( 
.A(n_2262),
.B(n_1919),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2211),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2187),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2067),
.B(n_1871),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2102),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2112),
.Y(n_2326)
);

NAND2xp33_ASAP7_75t_SL g2327 ( 
.A(n_2298),
.B(n_1943),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2107),
.B(n_1988),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2112),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2076),
.B(n_1874),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2275),
.A2(n_1758),
.B1(n_1868),
.B2(n_1883),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2078),
.B(n_1874),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2114),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2289),
.B(n_1919),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2234),
.A2(n_1888),
.B1(n_1850),
.B2(n_1856),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2114),
.Y(n_2336)
);

INVxp67_ASAP7_75t_SL g2337 ( 
.A(n_2025),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2187),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2000),
.B(n_1928),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2120),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2223),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2223),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2233),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2139),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_L g2345 ( 
.A(n_2102),
.B(n_2111),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2139),
.Y(n_2346)
);

AND3x1_ASAP7_75t_L g2347 ( 
.A(n_2141),
.B(n_1825),
.C(n_1777),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2149),
.Y(n_2348)
);

AOI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2241),
.A2(n_1888),
.B1(n_1853),
.B2(n_1856),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2233),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_2020),
.B(n_1778),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_2102),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2235),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2235),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_2121),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2274),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2082),
.B(n_1836),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2274),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1999),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_2094),
.Y(n_2360)
);

AO21x2_ASAP7_75t_L g2361 ( 
.A1(n_2029),
.A2(n_1832),
.B(n_1779),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2149),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2160),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1999),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2111),
.B(n_1928),
.Y(n_2365)
);

INVxp67_ASAP7_75t_L g2366 ( 
.A(n_1991),
.Y(n_2366)
);

OAI21xp33_ASAP7_75t_SL g2367 ( 
.A1(n_2023),
.A2(n_1926),
.B(n_1832),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2160),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2089),
.B(n_1874),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2023),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_1992),
.B(n_1928),
.Y(n_2371)
);

NOR2x1p5_ASAP7_75t_L g2372 ( 
.A(n_2052),
.B(n_1891),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_2083),
.B(n_1791),
.Y(n_2373)
);

INVx3_ASAP7_75t_L g2374 ( 
.A(n_2303),
.Y(n_2374)
);

INVx2_ASAP7_75t_SL g2375 ( 
.A(n_2123),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2173),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2303),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2173),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2032),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2027),
.Y(n_2380)
);

AND2x2_ASAP7_75t_SL g2381 ( 
.A(n_2259),
.B(n_1928),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2027),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2032),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2053),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_2219),
.A2(n_1853),
.B1(n_1836),
.B2(n_1818),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2124),
.Y(n_2386)
);

INVxp33_ASAP7_75t_L g2387 ( 
.A(n_2140),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2097),
.B(n_1873),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2029),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2053),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2057),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2111),
.B(n_1943),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_2204),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2083),
.B(n_1791),
.Y(n_2394)
);

INVx4_ASAP7_75t_L g2395 ( 
.A(n_2204),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2065),
.B(n_1815),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2057),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2188),
.B(n_1815),
.Y(n_2398)
);

INVxp67_ASAP7_75t_L g2399 ( 
.A(n_2034),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2030),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2030),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2058),
.Y(n_2402)
);

INVx4_ASAP7_75t_L g2403 ( 
.A(n_2204),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2058),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2039),
.A2(n_1818),
.B1(n_1834),
.B2(n_1815),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2083),
.B(n_1962),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2063),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2063),
.Y(n_2408)
);

BUFx2_ASAP7_75t_L g2409 ( 
.A(n_2165),
.Y(n_2409)
);

INVx5_ASAP7_75t_L g2410 ( 
.A(n_2236),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2092),
.Y(n_2411)
);

NAND3xp33_ASAP7_75t_L g2412 ( 
.A(n_2066),
.B(n_1960),
.C(n_1943),
.Y(n_2412)
);

AND2x2_ASAP7_75t_SL g2413 ( 
.A(n_2266),
.B(n_1960),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2118),
.B(n_1960),
.Y(n_2414)
);

NAND2xp33_ASAP7_75t_L g2415 ( 
.A(n_2236),
.B(n_1960),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2051),
.Y(n_2416)
);

INVx4_ASAP7_75t_L g2417 ( 
.A(n_2236),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2190),
.B(n_1815),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_1990),
.B(n_1971),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2092),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2151),
.B(n_1961),
.Y(n_2421)
);

OAI22xp33_ASAP7_75t_L g2422 ( 
.A1(n_2141),
.A2(n_2179),
.B1(n_2210),
.B2(n_2009),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2106),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_2051),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2170),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2230),
.A2(n_1818),
.B1(n_1847),
.B2(n_1834),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_2161),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_1998),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2231),
.A2(n_1818),
.B1(n_1847),
.B2(n_1834),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_2072),
.B(n_1961),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2106),
.Y(n_2431)
);

CKINVDCx14_ASAP7_75t_R g2432 ( 
.A(n_2041),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2115),
.Y(n_2433)
);

AND3x1_ASAP7_75t_L g2434 ( 
.A(n_2179),
.B(n_1859),
.C(n_1869),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_2085),
.B(n_1961),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2201),
.B(n_1834),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2205),
.B(n_1847),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2115),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2003),
.Y(n_2439)
);

NAND2xp33_ASAP7_75t_L g2440 ( 
.A(n_2079),
.B(n_1961),
.Y(n_2440)
);

INVx2_ASAP7_75t_SL g2441 ( 
.A(n_2253),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2122),
.Y(n_2442)
);

BUFx3_ASAP7_75t_L g2443 ( 
.A(n_2096),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2122),
.Y(n_2444)
);

INVx5_ASAP7_75t_L g2445 ( 
.A(n_2079),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2133),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2133),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2064),
.B(n_1971),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2216),
.B(n_1847),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2146),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2146),
.Y(n_2451)
);

AOI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2253),
.A2(n_1862),
.B1(n_1855),
.B2(n_1926),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2150),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2276),
.B(n_1971),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_2096),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2150),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2021),
.B(n_1971),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2010),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2159),
.Y(n_2459)
);

INVxp67_ASAP7_75t_SL g2460 ( 
.A(n_2077),
.Y(n_2460)
);

INVx3_ASAP7_75t_L g2461 ( 
.A(n_2013),
.Y(n_2461)
);

INVx3_ASAP7_75t_L g2462 ( 
.A(n_2291),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2291),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2220),
.B(n_1855),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2225),
.B(n_1855),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2159),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2019),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2238),
.A2(n_1862),
.B1(n_1855),
.B2(n_1823),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2304),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2011),
.B(n_1974),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2055),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2304),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2279),
.B(n_1974),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_SL g2474 ( 
.A1(n_1996),
.A2(n_1979),
.B1(n_1974),
.B2(n_1910),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2309),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2240),
.B(n_1862),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2283),
.B(n_1974),
.Y(n_2477)
);

NAND2xp33_ASAP7_75t_L g2478 ( 
.A(n_2079),
.B(n_1979),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2056),
.Y(n_2479)
);

AOI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2247),
.A2(n_1862),
.B1(n_1840),
.B2(n_1843),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2199),
.B(n_1915),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2069),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2088),
.Y(n_2483)
);

OR2x2_ASAP7_75t_SL g2484 ( 
.A(n_1993),
.B(n_1979),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_2195),
.B(n_1979),
.Y(n_2485)
);

INVxp33_ASAP7_75t_SL g2486 ( 
.A(n_2113),
.Y(n_2486)
);

INVx5_ASAP7_75t_L g2487 ( 
.A(n_2079),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2309),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2208),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2033),
.B(n_1915),
.Y(n_2490)
);

INVx2_ASAP7_75t_SL g2491 ( 
.A(n_2255),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2091),
.Y(n_2492)
);

INVx4_ASAP7_75t_L g2493 ( 
.A(n_2208),
.Y(n_2493)
);

INVxp33_ASAP7_75t_L g2494 ( 
.A(n_2183),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2099),
.Y(n_2495)
);

XNOR2xp5_ASAP7_75t_L g2496 ( 
.A(n_2094),
.B(n_1837),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2101),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2258),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2116),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2254),
.B(n_1841),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2129),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2131),
.Y(n_2502)
);

INVx4_ASAP7_75t_L g2503 ( 
.A(n_2280),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2145),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2147),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2189),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2278),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2155),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2024),
.B(n_1754),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2294),
.B(n_1857),
.Y(n_2510)
);

NAND3xp33_ASAP7_75t_L g2511 ( 
.A(n_2185),
.B(n_1830),
.C(n_1869),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_2198),
.Y(n_2512)
);

BUFx10_ASAP7_75t_L g2513 ( 
.A(n_2186),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2157),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2162),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2203),
.B(n_1754),
.Y(n_2516)
);

INVx1_ASAP7_75t_SL g2517 ( 
.A(n_2164),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2169),
.Y(n_2518)
);

NAND2xp33_ASAP7_75t_L g2519 ( 
.A(n_2214),
.B(n_1754),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2175),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2293),
.B(n_1845),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2050),
.A2(n_1816),
.B1(n_1775),
.B2(n_1790),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2176),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_2090),
.B(n_1754),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2181),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2127),
.B(n_1857),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2182),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2295),
.B(n_1751),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2093),
.B(n_1767),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2296),
.B(n_1870),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_2050),
.A2(n_1816),
.B1(n_1780),
.B2(n_1802),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_1994),
.B(n_1767),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_1995),
.B(n_1891),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2110),
.B(n_1751),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_2016),
.B(n_1767),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2288),
.B(n_1747),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_2105),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2028),
.B(n_1816),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2015),
.B(n_1747),
.Y(n_2539)
);

AND2x6_ASAP7_75t_L g2540 ( 
.A(n_2217),
.B(n_1767),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_2017),
.B(n_1870),
.Y(n_2541)
);

INVx5_ASAP7_75t_L g2542 ( 
.A(n_2017),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2004),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2267),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2285),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2264),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2264),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2117),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_1989),
.B(n_1869),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2026),
.B(n_1789),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_1989),
.B(n_1747),
.Y(n_2551)
);

OR2x6_ASAP7_75t_L g2552 ( 
.A(n_2143),
.B(n_1779),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2178),
.B(n_1870),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2301),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2135),
.B(n_1780),
.Y(n_2555)
);

AOI22xp33_ASAP7_75t_L g2556 ( 
.A1(n_1993),
.A2(n_1790),
.B1(n_1802),
.B2(n_1780),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2061),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2061),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2047),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_SL g2560 ( 
.A(n_2278),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2269),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2073),
.B(n_1790),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_1996),
.A2(n_2148),
.B1(n_2060),
.B2(n_2006),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2046),
.B(n_1802),
.Y(n_2564)
);

BUFx10_ASAP7_75t_L g2565 ( 
.A(n_2192),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2109),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2047),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2075),
.Y(n_2568)
);

OAI21xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2292),
.A2(n_1773),
.B(n_1772),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2269),
.Y(n_2570)
);

CKINVDCx20_ASAP7_75t_R g2571 ( 
.A(n_2119),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2143),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2036),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2202),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2148),
.A2(n_1807),
.B1(n_1811),
.B2(n_1805),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2248),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2281),
.Y(n_2577)
);

OR2x6_ASAP7_75t_L g2578 ( 
.A(n_2172),
.B(n_1805),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2012),
.B(n_1807),
.C(n_1805),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2178),
.B(n_1807),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2043),
.A2(n_1819),
.B1(n_1811),
.B2(n_1743),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_2261),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2281),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2086),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2048),
.Y(n_2585)
);

INVx2_ASAP7_75t_SL g2586 ( 
.A(n_2265),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2172),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2062),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2007),
.B(n_1789),
.Y(n_2589)
);

AND2x6_ASAP7_75t_L g2590 ( 
.A(n_2217),
.B(n_1789),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2136),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2132),
.B(n_1811),
.Y(n_2592)
);

OAI22xp33_ASAP7_75t_SL g2593 ( 
.A1(n_2202),
.A2(n_1819),
.B1(n_51),
.B2(n_49),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2284),
.Y(n_2594)
);

OR2x6_ASAP7_75t_L g2595 ( 
.A(n_2270),
.B(n_1819),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2284),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2060),
.A2(n_1743),
.B1(n_1793),
.B2(n_1789),
.Y(n_2597)
);

INVxp33_ASAP7_75t_L g2598 ( 
.A(n_2138),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2070),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2044),
.Y(n_2600)
);

CKINVDCx16_ASAP7_75t_R g2601 ( 
.A(n_2002),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2044),
.B(n_1772),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2246),
.B(n_1773),
.Y(n_2603)
);

AO22x2_ASAP7_75t_L g2604 ( 
.A1(n_2249),
.A2(n_52),
.B1(n_53),
.B2(n_51),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2270),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2272),
.B(n_1793),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2070),
.Y(n_2607)
);

INVx4_ASAP7_75t_L g2608 ( 
.A(n_2087),
.Y(n_2608)
);

AND2x6_ASAP7_75t_L g2609 ( 
.A(n_2292),
.B(n_1793),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2277),
.B(n_1793),
.Y(n_2610)
);

AND2x2_ASAP7_75t_SL g2611 ( 
.A(n_2282),
.B(n_1794),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2087),
.Y(n_2612)
);

INVx5_ASAP7_75t_L g2613 ( 
.A(n_2221),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2001),
.A2(n_1743),
.B1(n_1716),
.B2(n_1794),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2302),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2302),
.Y(n_2616)
);

OAI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2287),
.A2(n_1812),
.B1(n_1784),
.B2(n_1801),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2152),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2221),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2290),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2045),
.B(n_1784),
.Y(n_2621)
);

XOR2xp5_ASAP7_75t_L g2622 ( 
.A(n_2144),
.B(n_1794),
.Y(n_2622)
);

OR2x6_ASAP7_75t_L g2623 ( 
.A(n_2163),
.B(n_1743),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2256),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_SL g2625 ( 
.A(n_2232),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2054),
.B(n_1812),
.Y(n_2626)
);

INVx4_ASAP7_75t_L g2627 ( 
.A(n_2232),
.Y(n_2627)
);

XNOR2xp5_ASAP7_75t_L g2628 ( 
.A(n_2154),
.B(n_177),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2305),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2307),
.A2(n_1810),
.B1(n_1801),
.B2(n_1794),
.Y(n_2630)
);

OAI22xp33_ASAP7_75t_SL g2631 ( 
.A1(n_2299),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2152),
.Y(n_2632)
);

NOR2x1p5_ASAP7_75t_L g2633 ( 
.A(n_2180),
.B(n_1716),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2080),
.B(n_1801),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2037),
.B(n_1801),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2299),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2153),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2008),
.B(n_1810),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2153),
.Y(n_2639)
);

OR2x6_ASAP7_75t_L g2640 ( 
.A(n_2166),
.B(n_1810),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2005),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2300),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2166),
.B(n_1810),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_2074),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2197),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2008),
.B(n_2022),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2018),
.B(n_1700),
.Y(n_2647)
);

AND3x2_ASAP7_75t_L g2648 ( 
.A(n_2197),
.B(n_52),
.C(n_53),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2308),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2206),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2206),
.Y(n_2651)
);

XNOR2xp5_ASAP7_75t_L g2652 ( 
.A(n_2156),
.B(n_54),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2158),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2031),
.B(n_1700),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2229),
.Y(n_2655)
);

OAI21xp33_ASAP7_75t_SL g2656 ( 
.A1(n_2200),
.A2(n_2209),
.B(n_2207),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2229),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2245),
.Y(n_2658)
);

NAND2xp33_ASAP7_75t_L g2659 ( 
.A(n_2212),
.B(n_1700),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2245),
.Y(n_2660)
);

INVxp67_ASAP7_75t_L g2661 ( 
.A(n_2167),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2103),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2103),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2104),
.Y(n_2664)
);

BUFx3_ASAP7_75t_L g2665 ( 
.A(n_2619),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2318),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2318),
.Y(n_2667)
);

BUFx3_ASAP7_75t_L g2668 ( 
.A(n_2619),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2404),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2319),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2544),
.B(n_2239),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2328),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2441),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2582),
.B(n_2035),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2404),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2407),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2395),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2454),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2598),
.B(n_2168),
.Y(n_2679)
);

BUFx3_ASAP7_75t_L g2680 ( 
.A(n_2587),
.Y(n_2680)
);

AND2x4_ASAP7_75t_L g2681 ( 
.A(n_2373),
.B(n_2394),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2381),
.B(n_2142),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2407),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2408),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2587),
.Y(n_2685)
);

BUFx6f_ASAP7_75t_L g2686 ( 
.A(n_2424),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2408),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_L g2688 ( 
.A(n_2424),
.Y(n_2688)
);

AOI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2414),
.A2(n_2193),
.B1(n_2194),
.B2(n_2171),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2319),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2323),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2411),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2424),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2598),
.B(n_2196),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2411),
.Y(n_2695)
);

AND2x6_ASAP7_75t_L g2696 ( 
.A(n_2469),
.B(n_2213),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2381),
.B(n_2042),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2328),
.Y(n_2698)
);

INVx4_ASAP7_75t_L g2699 ( 
.A(n_2424),
.Y(n_2699)
);

AND2x4_ASAP7_75t_L g2700 ( 
.A(n_2373),
.B(n_2222),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2420),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2420),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2544),
.B(n_2545),
.Y(n_2703)
);

INVx4_ASAP7_75t_L g2704 ( 
.A(n_2410),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2423),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_2373),
.B(n_2227),
.Y(n_2706)
);

OAI221xp5_ASAP7_75t_L g2707 ( 
.A1(n_2656),
.A2(n_2237),
.B1(n_2250),
.B2(n_2242),
.C(n_2228),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2323),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2545),
.B(n_2215),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2325),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2338),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2338),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2394),
.B(n_2251),
.Y(n_2713)
);

INVx4_ASAP7_75t_L g2714 ( 
.A(n_2410),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2454),
.Y(n_2715)
);

HB1xp67_ASAP7_75t_L g2716 ( 
.A(n_2441),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2423),
.Y(n_2717)
);

INVxp67_ASAP7_75t_L g2718 ( 
.A(n_2473),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2341),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2433),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2325),
.Y(n_2721)
);

NAND2x1p5_ASAP7_75t_L g2722 ( 
.A(n_2445),
.B(n_1700),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2341),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2394),
.B(n_1842),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2342),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2342),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2410),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2325),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2473),
.Y(n_2729)
);

NAND2x1p5_ASAP7_75t_L g2730 ( 
.A(n_2445),
.B(n_1708),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2395),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2636),
.A2(n_2252),
.B1(n_2226),
.B2(n_2104),
.Y(n_2732)
);

INVx3_ASAP7_75t_L g2733 ( 
.A(n_2395),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2433),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2388),
.B(n_2243),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2438),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2438),
.Y(n_2737)
);

BUFx10_ASAP7_75t_L g2738 ( 
.A(n_2549),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2343),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2442),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2625),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2337),
.B(n_2260),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2442),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2339),
.B(n_2263),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2403),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2446),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2625),
.Y(n_2747)
);

BUFx3_ASAP7_75t_L g2748 ( 
.A(n_2406),
.Y(n_2748)
);

OA21x2_ASAP7_75t_L g2749 ( 
.A1(n_2320),
.A2(n_2049),
.B(n_2038),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2446),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2554),
.B(n_2273),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2447),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2447),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2343),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2350),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2357),
.B(n_2095),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2450),
.Y(n_2757)
);

INVx3_ASAP7_75t_L g2758 ( 
.A(n_2403),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2350),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2661),
.B(n_2244),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2366),
.B(n_2059),
.Y(n_2761)
);

HB1xp67_ASAP7_75t_L g2762 ( 
.A(n_2414),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2353),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2406),
.B(n_1842),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2359),
.B(n_2271),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2450),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2625),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2406),
.B(n_2312),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2422),
.A2(n_2297),
.B1(n_2137),
.B2(n_2191),
.Y(n_2769)
);

AO22x2_ASAP7_75t_L g2770 ( 
.A1(n_2570),
.A2(n_2040),
.B1(n_2068),
.B2(n_2177),
.Y(n_2770)
);

OAI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2570),
.A2(n_2134),
.B1(n_2130),
.B2(n_2126),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2353),
.Y(n_2772)
);

AND2x4_ASAP7_75t_L g2773 ( 
.A(n_2312),
.B(n_1842),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2517),
.B(n_2081),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2354),
.Y(n_2775)
);

OR2x6_ASAP7_75t_L g2776 ( 
.A(n_2574),
.B(n_1708),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2403),
.Y(n_2777)
);

CKINVDCx20_ASAP7_75t_R g2778 ( 
.A(n_2507),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2453),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2416),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2409),
.Y(n_2781)
);

AND2x6_ASAP7_75t_L g2782 ( 
.A(n_2469),
.B(n_2224),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2359),
.B(n_2098),
.Y(n_2783)
);

AO22x2_ASAP7_75t_L g2784 ( 
.A1(n_2570),
.A2(n_2268),
.B1(n_2257),
.B2(n_2125),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2354),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2364),
.B(n_2370),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2453),
.Y(n_2787)
);

NAND2x1p5_ASAP7_75t_L g2788 ( 
.A(n_2445),
.B(n_1720),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2477),
.B(n_2084),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2356),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2498),
.B(n_2128),
.Y(n_2791)
);

AND2x4_ASAP7_75t_L g2792 ( 
.A(n_2312),
.B(n_1842),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_2560),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2356),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2494),
.B(n_2108),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2448),
.B(n_1708),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2494),
.B(n_54),
.Y(n_2797)
);

AND2x4_ASAP7_75t_L g2798 ( 
.A(n_2448),
.B(n_2351),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_2560),
.Y(n_2799)
);

INVx4_ASAP7_75t_L g2800 ( 
.A(n_2410),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2417),
.Y(n_2801)
);

INVx3_ASAP7_75t_L g2802 ( 
.A(n_2417),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2425),
.B(n_179),
.Y(n_2803)
);

INVx4_ASAP7_75t_L g2804 ( 
.A(n_2410),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2399),
.B(n_55),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2351),
.B(n_1708),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2477),
.B(n_688),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2512),
.Y(n_2808)
);

OAI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2640),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2417),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2358),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2325),
.Y(n_2812)
);

OR2x2_ASAP7_75t_SL g2813 ( 
.A(n_2601),
.B(n_55),
.Y(n_2813)
);

NAND2x1p5_ASAP7_75t_L g2814 ( 
.A(n_2445),
.B(n_1709),
.Y(n_2814)
);

AND2x6_ASAP7_75t_L g2815 ( 
.A(n_2472),
.B(n_1709),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_L g2816 ( 
.A(n_2352),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2506),
.Y(n_2817)
);

INVxp67_ASAP7_75t_L g2818 ( 
.A(n_2324),
.Y(n_2818)
);

INVx4_ASAP7_75t_L g2819 ( 
.A(n_2352),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2358),
.Y(n_2820)
);

INVxp67_ASAP7_75t_L g2821 ( 
.A(n_2324),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2371),
.B(n_56),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2379),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2383),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2364),
.B(n_1709),
.Y(n_2825)
);

INVx2_ASAP7_75t_SL g2826 ( 
.A(n_2574),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2384),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2370),
.B(n_1709),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2492),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2492),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2430),
.B(n_58),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2390),
.Y(n_2832)
);

BUFx2_ASAP7_75t_L g2833 ( 
.A(n_2572),
.Y(n_2833)
);

OR2x6_ASAP7_75t_L g2834 ( 
.A(n_2574),
.B(n_1719),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2391),
.Y(n_2835)
);

BUFx3_ASAP7_75t_L g2836 ( 
.A(n_2416),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2430),
.B(n_58),
.Y(n_2837)
);

AND2x6_ASAP7_75t_L g2838 ( 
.A(n_2472),
.B(n_1719),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2397),
.Y(n_2839)
);

NAND3xp33_ASAP7_75t_L g2840 ( 
.A(n_2412),
.B(n_2419),
.C(n_2474),
.Y(n_2840)
);

BUFx3_ASAP7_75t_L g2841 ( 
.A(n_2443),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2352),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2497),
.Y(n_2843)
);

INVxp67_ASAP7_75t_L g2844 ( 
.A(n_2330),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2402),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2431),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2497),
.Y(n_2847)
);

OR2x2_ASAP7_75t_L g2848 ( 
.A(n_2314),
.B(n_180),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2444),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2490),
.B(n_181),
.Y(n_2850)
);

AO22x2_ASAP7_75t_L g2851 ( 
.A1(n_2615),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2451),
.Y(n_2852)
);

INVx1_ASAP7_75t_SL g2853 ( 
.A(n_2562),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2382),
.B(n_2316),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2456),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2352),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2459),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2351),
.B(n_1719),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2560),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2466),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2393),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2443),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2382),
.Y(n_2863)
);

BUFx2_ASAP7_75t_L g2864 ( 
.A(n_2595),
.Y(n_2864)
);

AND2x6_ASAP7_75t_L g2865 ( 
.A(n_2475),
.B(n_1719),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2393),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2501),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2393),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2498),
.B(n_1720),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2501),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2498),
.B(n_1720),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2502),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2330),
.B(n_674),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2481),
.B(n_1720),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2317),
.A2(n_1729),
.B1(n_1707),
.B2(n_183),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2502),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2508),
.Y(n_2877)
);

BUFx2_ASAP7_75t_L g2878 ( 
.A(n_2595),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2508),
.Y(n_2879)
);

BUFx4f_ASAP7_75t_L g2880 ( 
.A(n_2574),
.Y(n_2880)
);

INVx3_ASAP7_75t_L g2881 ( 
.A(n_2393),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2387),
.B(n_59),
.Y(n_2882)
);

NAND3xp33_ASAP7_75t_L g2883 ( 
.A(n_2317),
.B(n_1729),
.C(n_1707),
.Y(n_2883)
);

AND2x6_ASAP7_75t_L g2884 ( 
.A(n_2475),
.B(n_1729),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2515),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2455),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2387),
.B(n_59),
.Y(n_2887)
);

AND2x6_ASAP7_75t_L g2888 ( 
.A(n_2488),
.B(n_1729),
.Y(n_2888)
);

INVx4_ASAP7_75t_L g2889 ( 
.A(n_2493),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2488),
.B(n_60),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2608),
.B(n_60),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2515),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2518),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_2498),
.B(n_1707),
.Y(n_2894)
);

BUFx2_ASAP7_75t_L g2895 ( 
.A(n_2595),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2518),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2460),
.B(n_61),
.Y(n_2897)
);

BUFx3_ASAP7_75t_L g2898 ( 
.A(n_2455),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2467),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_2481),
.B(n_1707),
.Y(n_2900)
);

AND2x6_ASAP7_75t_L g2901 ( 
.A(n_2583),
.B(n_2594),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2471),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2481),
.B(n_182),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2428),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2608),
.B(n_61),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2332),
.B(n_679),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2457),
.B(n_182),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2489),
.Y(n_2908)
);

AOI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2413),
.A2(n_184),
.B1(n_185),
.B2(n_183),
.Y(n_2909)
);

INVx4_ASAP7_75t_L g2910 ( 
.A(n_2493),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2479),
.Y(n_2911)
);

BUFx6f_ASAP7_75t_L g2912 ( 
.A(n_2489),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2493),
.Y(n_2913)
);

BUFx6f_ASAP7_75t_L g2914 ( 
.A(n_2542),
.Y(n_2914)
);

AND2x4_ASAP7_75t_L g2915 ( 
.A(n_2340),
.B(n_185),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2482),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2608),
.B(n_62),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2483),
.Y(n_2918)
);

AND2x6_ASAP7_75t_L g2919 ( 
.A(n_2583),
.B(n_62),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2380),
.B(n_62),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2607),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2495),
.Y(n_2922)
);

BUFx3_ASAP7_75t_L g2923 ( 
.A(n_2507),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2380),
.B(n_63),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2332),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2428),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2499),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2504),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2428),
.Y(n_2929)
);

AND2x4_ASAP7_75t_L g2930 ( 
.A(n_2340),
.B(n_186),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2380),
.B(n_63),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2439),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2514),
.Y(n_2933)
);

OR2x2_ASAP7_75t_SL g2934 ( 
.A(n_2511),
.B(n_2605),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2605),
.Y(n_2935)
);

INVx1_ASAP7_75t_SL g2936 ( 
.A(n_2562),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2543),
.B(n_63),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2624),
.B(n_64),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2484),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2543),
.B(n_65),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2439),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2413),
.A2(n_188),
.B1(n_189),
.B2(n_187),
.Y(n_2942)
);

A2O1A1Ixp33_ASAP7_75t_L g2943 ( 
.A1(n_2491),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2520),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2527),
.Y(n_2945)
);

INVx3_ASAP7_75t_L g2946 ( 
.A(n_2311),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2542),
.Y(n_2947)
);

BUFx3_ASAP7_75t_L g2948 ( 
.A(n_2605),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2439),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2458),
.Y(n_2950)
);

AO22x2_ASAP7_75t_L g2951 ( 
.A1(n_2615),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2951)
);

BUFx3_ASAP7_75t_L g2952 ( 
.A(n_2605),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2331),
.B(n_187),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2458),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2604),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2458),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2542),
.Y(n_2957)
);

AND2x2_ASAP7_75t_SL g2958 ( 
.A(n_2831),
.B(n_2440),
.Y(n_2958)
);

OR2x2_ASAP7_75t_L g2959 ( 
.A(n_2698),
.B(n_2653),
.Y(n_2959)
);

INVx2_ASAP7_75t_SL g2960 ( 
.A(n_2880),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_2778),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2817),
.B(n_2679),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2880),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2831),
.A2(n_2604),
.B1(n_2649),
.B2(n_2631),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2678),
.B(n_2715),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2837),
.A2(n_2604),
.B1(n_2629),
.B2(n_2620),
.Y(n_2966)
);

NOR2x2_ASAP7_75t_L g2967 ( 
.A(n_2776),
.B(n_2640),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2694),
.B(n_2369),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2704),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2678),
.B(n_2369),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2704),
.Y(n_2971)
);

O2A1O1Ixp33_ASAP7_75t_L g2972 ( 
.A1(n_2822),
.A2(n_2334),
.B(n_2435),
.C(n_2485),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2666),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_2741),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2840),
.A2(n_2334),
.B1(n_2310),
.B2(n_2405),
.Y(n_2975)
);

AO22x1_ASAP7_75t_L g2976 ( 
.A1(n_2822),
.A2(n_2542),
.B1(n_2486),
.B2(n_2360),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2715),
.B(n_2576),
.Y(n_2977)
);

OAI22xp33_ASAP7_75t_SL g2978 ( 
.A1(n_2682),
.A2(n_2640),
.B1(n_2643),
.B2(n_2435),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2714),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2921),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2718),
.B(n_2576),
.Y(n_2981)
);

OR2x2_ASAP7_75t_SL g2982 ( 
.A(n_2803),
.B(n_2616),
.Y(n_2982)
);

NAND2x1_ASAP7_75t_L g2983 ( 
.A(n_2714),
.B(n_2374),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2679),
.A2(n_2486),
.B1(n_2327),
.B2(n_2347),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2718),
.B(n_2576),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2921),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2694),
.B(n_2653),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2729),
.B(n_2586),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2729),
.B(n_2762),
.Y(n_2989)
);

AO22x1_ASAP7_75t_L g2990 ( 
.A1(n_2732),
.A2(n_2542),
.B1(n_2360),
.B2(n_2613),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2762),
.B(n_2586),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2667),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2823),
.Y(n_2993)
);

NOR2xp33_ASAP7_75t_SL g2994 ( 
.A(n_2923),
.B(n_2627),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2840),
.B(n_2445),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2824),
.Y(n_2996)
);

AOI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2854),
.A2(n_2519),
.B(n_2478),
.Y(n_2997)
);

AOI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2760),
.A2(n_2682),
.B1(n_2795),
.B2(n_2774),
.Y(n_2998)
);

OR2x6_ASAP7_75t_L g2999 ( 
.A(n_2914),
.B(n_2627),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2914),
.Y(n_3000)
);

NAND2x1p5_ASAP7_75t_L g3001 ( 
.A(n_2914),
.B(n_2957),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2703),
.B(n_2355),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2817),
.B(n_2427),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2670),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2853),
.B(n_2646),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2837),
.A2(n_2604),
.B1(n_2643),
.B2(n_2640),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2827),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2760),
.B(n_2484),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2832),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2672),
.B(n_2427),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2835),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2703),
.B(n_2355),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2735),
.B(n_2744),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2735),
.B(n_2375),
.Y(n_3014)
);

OR2x6_ASAP7_75t_L g3015 ( 
.A(n_2947),
.B(n_2627),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2768),
.B(n_2375),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2744),
.B(n_2487),
.Y(n_3017)
);

INVx4_ASAP7_75t_L g3018 ( 
.A(n_2913),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2853),
.B(n_2427),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2818),
.B(n_2386),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2839),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2690),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2742),
.B(n_2487),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2691),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_2936),
.B(n_2513),
.Y(n_3025)
);

NOR2x1p5_ASAP7_75t_L g3026 ( 
.A(n_2748),
.B(n_2641),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2727),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2818),
.B(n_2386),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2708),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2845),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2936),
.B(n_2646),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2698),
.B(n_2513),
.Y(n_3032)
);

BUFx3_ASAP7_75t_L g3033 ( 
.A(n_2886),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2711),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2821),
.B(n_2513),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2789),
.B(n_2526),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2712),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2665),
.Y(n_3038)
);

A2O1A1Ixp33_ASAP7_75t_L g3039 ( 
.A1(n_2707),
.A2(n_2327),
.B(n_2491),
.C(n_2470),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_L g3040 ( 
.A(n_2821),
.B(n_2565),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2844),
.B(n_2526),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2844),
.B(n_2510),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2719),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2925),
.B(n_2510),
.Y(n_3044)
);

BUFx3_ASAP7_75t_L g3045 ( 
.A(n_2886),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2925),
.B(n_2599),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_2781),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2798),
.B(n_2565),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2886),
.Y(n_3049)
);

INVxp67_ASAP7_75t_L g3050 ( 
.A(n_2808),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2798),
.B(n_2565),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2756),
.B(n_2612),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2756),
.B(n_2555),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2795),
.A2(n_2633),
.B1(n_2421),
.B2(n_2580),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2707),
.A2(n_2563),
.B1(n_2429),
.B2(n_2426),
.Y(n_3055)
);

INVxp67_ASAP7_75t_L g3056 ( 
.A(n_2673),
.Y(n_3056)
);

INVx2_ASAP7_75t_SL g3057 ( 
.A(n_2668),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2751),
.B(n_2553),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_2727),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2751),
.B(n_2546),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_2761),
.B(n_2421),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2846),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2723),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2938),
.B(n_2546),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2725),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2849),
.Y(n_3066)
);

NOR2xp67_ASAP7_75t_L g3067 ( 
.A(n_2699),
.B(n_2613),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2938),
.B(n_2547),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2761),
.B(n_2547),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2689),
.B(n_2616),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2742),
.B(n_2561),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2697),
.B(n_2600),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2671),
.B(n_2561),
.Y(n_3073)
);

BUFx8_ASAP7_75t_L g3074 ( 
.A(n_2908),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2697),
.B(n_2600),
.Y(n_3075)
);

INVx2_ASAP7_75t_SL g3076 ( 
.A(n_2908),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2671),
.B(n_2577),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2852),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2807),
.B(n_2623),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2774),
.A2(n_2706),
.B1(n_2713),
.B2(n_2700),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2850),
.B(n_2577),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2709),
.B(n_2596),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2709),
.B(n_2596),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2769),
.B(n_2396),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_2908),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2681),
.B(n_2613),
.Y(n_3086)
);

NOR2xp67_ASAP7_75t_L g3087 ( 
.A(n_2699),
.B(n_2613),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2769),
.B(n_2607),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_SL g3089 ( 
.A(n_2780),
.Y(n_3089)
);

INVx2_ASAP7_75t_SL g3090 ( 
.A(n_2912),
.Y(n_3090)
);

INVx3_ASAP7_75t_L g3091 ( 
.A(n_2800),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_L g3092 ( 
.A(n_2732),
.B(n_2622),
.Y(n_3092)
);

BUFx3_ASAP7_75t_L g3093 ( 
.A(n_2912),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2674),
.B(n_2623),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2681),
.B(n_2607),
.Y(n_3095)
);

NAND2xp33_ASAP7_75t_SL g3096 ( 
.A(n_2947),
.B(n_2372),
.Y(n_3096)
);

AOI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_2700),
.A2(n_2644),
.B1(n_2642),
.B2(n_2434),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2706),
.B(n_2641),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2873),
.B(n_2623),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2747),
.Y(n_3100)
);

NAND3xp33_ASAP7_75t_L g3101 ( 
.A(n_2909),
.B(n_2628),
.C(n_2652),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2713),
.B(n_2641),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2906),
.B(n_2623),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2939),
.A2(n_2643),
.B1(n_2594),
.B2(n_2583),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2726),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2739),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2768),
.B(n_2613),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2791),
.A2(n_2642),
.B1(n_2537),
.B2(n_2566),
.Y(n_3108)
);

INVx8_ASAP7_75t_L g3109 ( 
.A(n_2776),
.Y(n_3109)
);

OAI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_2855),
.A2(n_2385),
.B1(n_2468),
.B2(n_2480),
.Y(n_3110)
);

AOI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_2791),
.A2(n_2537),
.B1(n_2566),
.B2(n_2907),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2696),
.B(n_2594),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2800),
.Y(n_3113)
);

AOI221xp5_ASAP7_75t_L g3114 ( 
.A1(n_2809),
.A2(n_2652),
.B1(n_2593),
.B2(n_2662),
.C(n_2567),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2947),
.B(n_2541),
.Y(n_3115)
);

INVx3_ASAP7_75t_L g3116 ( 
.A(n_2804),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2696),
.B(n_2618),
.Y(n_3117)
);

OAI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2953),
.A2(n_2320),
.B(n_2539),
.Y(n_3118)
);

BUFx6f_ASAP7_75t_L g3119 ( 
.A(n_2957),
.Y(n_3119)
);

NOR2xp67_ASAP7_75t_L g3120 ( 
.A(n_2889),
.B(n_2533),
.Y(n_3120)
);

OAI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2953),
.A2(n_2485),
.B(n_2470),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2854),
.A2(n_2519),
.B(n_2478),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2754),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2955),
.A2(n_2643),
.B1(n_2632),
.B2(n_2637),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2857),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_2673),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2957),
.B(n_2541),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2860),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2955),
.A2(n_2632),
.B1(n_2637),
.B2(n_2618),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_2767),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2783),
.A2(n_2487),
.B1(n_2611),
.B2(n_2566),
.Y(n_3131)
);

NAND3xp33_ASAP7_75t_L g3132 ( 
.A(n_2942),
.B(n_2556),
.C(n_2579),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2696),
.B(n_2639),
.Y(n_3133)
);

INVx4_ASAP7_75t_L g3134 ( 
.A(n_2913),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_SL g3135 ( 
.A(n_2793),
.B(n_2571),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2897),
.B(n_2487),
.Y(n_3136)
);

A2O1A1Ixp33_ASAP7_75t_L g3137 ( 
.A1(n_2875),
.A2(n_2537),
.B(n_2591),
.C(n_2440),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2696),
.B(n_2639),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2851),
.A2(n_2650),
.B1(n_2651),
.B2(n_2645),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2716),
.B(n_2645),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2716),
.B(n_2650),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_2833),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2755),
.Y(n_3143)
);

HB1xp67_ASAP7_75t_L g3144 ( 
.A(n_2786),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2759),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2863),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2797),
.B(n_2651),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2797),
.B(n_2655),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2771),
.B(n_2557),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2882),
.B(n_2638),
.Y(n_3150)
);

INVx8_ASAP7_75t_L g3151 ( 
.A(n_2776),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2851),
.A2(n_2657),
.B1(n_2658),
.B2(n_2655),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2897),
.B(n_2487),
.Y(n_3153)
);

NOR2xp67_ASAP7_75t_L g3154 ( 
.A(n_2889),
.B(n_2575),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2782),
.B(n_2657),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2782),
.B(n_2658),
.Y(n_3156)
);

NOR2xp67_ASAP7_75t_L g3157 ( 
.A(n_2910),
.B(n_2365),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2669),
.Y(n_3158)
);

INVx8_ASAP7_75t_L g3159 ( 
.A(n_2834),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2763),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2882),
.B(n_2638),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2772),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2782),
.B(n_2660),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2782),
.B(n_2901),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_2912),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2675),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2775),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_2935),
.Y(n_3168)
);

NOR3xp33_ASAP7_75t_SL g3169 ( 
.A(n_2809),
.B(n_2532),
.C(n_2635),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2887),
.B(n_2903),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2901),
.B(n_2660),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2903),
.B(n_2541),
.Y(n_3172)
);

OAI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_2891),
.A2(n_2664),
.B1(n_2663),
.B2(n_2595),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2901),
.B(n_2664),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2785),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_SL g3176 ( 
.A(n_2764),
.B(n_2496),
.Y(n_3176)
);

NAND3xp33_ASAP7_75t_SL g3177 ( 
.A(n_2891),
.B(n_2349),
.C(n_2335),
.Y(n_3177)
);

OR2x6_ASAP7_75t_L g3178 ( 
.A(n_2864),
.B(n_2578),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2794),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2901),
.B(n_2663),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2783),
.B(n_2558),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_3000),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2993),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2996),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2987),
.B(n_2905),
.Y(n_3185)
);

NAND2xp33_ASAP7_75t_L g3186 ( 
.A(n_3026),
.B(n_2913),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_3047),
.Y(n_3187)
);

BUFx6f_ASAP7_75t_L g3188 ( 
.A(n_3033),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3007),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3009),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2973),
.Y(n_3191)
);

OR2x2_ASAP7_75t_SL g3192 ( 
.A(n_3101),
.B(n_2848),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3061),
.B(n_3144),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_3074),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3061),
.B(n_2937),
.Y(n_3195)
);

INVxp67_ASAP7_75t_L g3196 ( 
.A(n_3126),
.Y(n_3196)
);

OR2x2_ASAP7_75t_L g3197 ( 
.A(n_2959),
.B(n_2937),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3011),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_3016),
.B(n_2878),
.Y(n_3199)
);

INVxp33_ASAP7_75t_L g3200 ( 
.A(n_2987),
.Y(n_3200)
);

AND2x4_ASAP7_75t_L g3201 ( 
.A(n_3016),
.B(n_2895),
.Y(n_3201)
);

AND2x4_ASAP7_75t_L g3202 ( 
.A(n_3178),
.B(n_2948),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3006),
.A2(n_2951),
.B1(n_2851),
.B2(n_2917),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3021),
.Y(n_3204)
);

INVx3_ASAP7_75t_L g3205 ( 
.A(n_3000),
.Y(n_3205)
);

INVx4_ASAP7_75t_L g3206 ( 
.A(n_3109),
.Y(n_3206)
);

BUFx3_ASAP7_75t_L g3207 ( 
.A(n_3074),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3030),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3062),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2992),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_3045),
.Y(n_3211)
);

BUFx4f_ASAP7_75t_L g3212 ( 
.A(n_3109),
.Y(n_3212)
);

INVx4_ASAP7_75t_L g3213 ( 
.A(n_3109),
.Y(n_3213)
);

AOI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_2997),
.A2(n_3122),
.B(n_3121),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3066),
.Y(n_3215)
);

NOR2xp67_ASAP7_75t_L g3216 ( 
.A(n_3050),
.B(n_2826),
.Y(n_3216)
);

INVx3_ASAP7_75t_L g3217 ( 
.A(n_3000),
.Y(n_3217)
);

INVx2_ASAP7_75t_SL g3218 ( 
.A(n_3049),
.Y(n_3218)
);

AOI22xp5_ASAP7_75t_L g3219 ( 
.A1(n_2998),
.A2(n_3092),
.B1(n_3080),
.B2(n_2984),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3078),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3144),
.B(n_2940),
.Y(n_3221)
);

INVx5_ASAP7_75t_L g3222 ( 
.A(n_3151),
.Y(n_3222)
);

BUFx3_ASAP7_75t_L g3223 ( 
.A(n_3093),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3170),
.B(n_2784),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3013),
.B(n_2940),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3125),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_3150),
.B(n_2784),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_3126),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3004),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_3178),
.B(n_2952),
.Y(n_3230)
);

INVx3_ASAP7_75t_L g3231 ( 
.A(n_3000),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_3161),
.B(n_2784),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3128),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3140),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3022),
.Y(n_3235)
);

NAND2x1p5_ASAP7_75t_L g3236 ( 
.A(n_3086),
.B(n_2804),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_3038),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3141),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3024),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3146),
.Y(n_3240)
);

BUFx12f_ASAP7_75t_L g3241 ( 
.A(n_2961),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_3119),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3158),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3092),
.A2(n_2571),
.B1(n_2321),
.B2(n_2905),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3166),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_3029),
.Y(n_3246)
);

INVx2_ASAP7_75t_SL g3247 ( 
.A(n_3057),
.Y(n_3247)
);

INVx3_ASAP7_75t_L g3248 ( 
.A(n_3119),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2980),
.Y(n_3249)
);

INVx4_ASAP7_75t_L g3250 ( 
.A(n_3151),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3053),
.B(n_2786),
.Y(n_3251)
);

AND2x2_ASAP7_75t_SL g3252 ( 
.A(n_2958),
.B(n_2415),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3034),
.Y(n_3253)
);

HB1xp67_ASAP7_75t_L g3254 ( 
.A(n_2986),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3069),
.B(n_2676),
.Y(n_3255)
);

INVx3_ASAP7_75t_L g3256 ( 
.A(n_3119),
.Y(n_3256)
);

OR2x2_ASAP7_75t_L g3257 ( 
.A(n_3036),
.B(n_2962),
.Y(n_3257)
);

INVx2_ASAP7_75t_SL g3258 ( 
.A(n_3076),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3037),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3043),
.Y(n_3260)
);

INVx5_ASAP7_75t_L g3261 ( 
.A(n_3151),
.Y(n_3261)
);

AND2x6_ASAP7_75t_SL g3262 ( 
.A(n_3008),
.B(n_2887),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3063),
.Y(n_3263)
);

AOI22x1_ASAP7_75t_L g3264 ( 
.A1(n_2997),
.A2(n_2951),
.B1(n_2770),
.B2(n_2559),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_3168),
.Y(n_3265)
);

INVx3_ASAP7_75t_L g3266 ( 
.A(n_3119),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3065),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3058),
.B(n_2683),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_3132),
.A2(n_2917),
.B1(n_2951),
.B2(n_2770),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3105),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3178),
.B(n_2806),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_3054),
.B(n_2551),
.Y(n_3272)
);

CKINVDCx20_ASAP7_75t_R g3273 ( 
.A(n_2974),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_L g3274 ( 
.A(n_3008),
.B(n_2771),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_2968),
.B(n_2805),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3056),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3106),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3123),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3143),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3145),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3160),
.Y(n_3281)
);

INVx2_ASAP7_75t_SL g3282 ( 
.A(n_3085),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3162),
.Y(n_3283)
);

OR2x6_ASAP7_75t_L g3284 ( 
.A(n_3159),
.B(n_2552),
.Y(n_3284)
);

OAI22x1_ASAP7_75t_SL g3285 ( 
.A1(n_3100),
.A2(n_2799),
.B1(n_2859),
.B2(n_2813),
.Y(n_3285)
);

BUFx4f_ASAP7_75t_L g3286 ( 
.A(n_3159),
.Y(n_3286)
);

BUFx6f_ASAP7_75t_L g3287 ( 
.A(n_3159),
.Y(n_3287)
);

BUFx2_ASAP7_75t_L g3288 ( 
.A(n_3142),
.Y(n_3288)
);

BUFx6f_ASAP7_75t_L g3289 ( 
.A(n_3090),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_3114),
.A2(n_2770),
.B1(n_2648),
.B2(n_2919),
.Y(n_3290)
);

AND2x6_ASAP7_75t_L g3291 ( 
.A(n_3164),
.B(n_2389),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3084),
.B(n_2684),
.Y(n_3292)
);

INVx2_ASAP7_75t_SL g3293 ( 
.A(n_3165),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3071),
.B(n_2687),
.Y(n_3294)
);

AND2x4_ASAP7_75t_L g3295 ( 
.A(n_2960),
.B(n_2806),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3167),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_2958),
.B(n_2611),
.Y(n_3297)
);

INVxp67_ASAP7_75t_SL g3298 ( 
.A(n_2989),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3175),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_3108),
.B(n_2532),
.Y(n_3300)
);

OAI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_3114),
.A2(n_2765),
.B1(n_2902),
.B2(n_2899),
.Y(n_3301)
);

BUFx3_ASAP7_75t_L g3302 ( 
.A(n_3142),
.Y(n_3302)
);

AOI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3102),
.A2(n_2321),
.B1(n_2432),
.B2(n_2805),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_3018),
.Y(n_3304)
);

INVx3_ASAP7_75t_L g3305 ( 
.A(n_3018),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3052),
.B(n_2692),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3179),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3149),
.B(n_3070),
.Y(n_3308)
);

INVx3_ASAP7_75t_L g3309 ( 
.A(n_3134),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2977),
.Y(n_3310)
);

INVx2_ASAP7_75t_SL g3311 ( 
.A(n_3130),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3098),
.B(n_2432),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_3102),
.B(n_3070),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_3005),
.B(n_2915),
.Y(n_3314)
);

AOI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_3072),
.A2(n_2321),
.B1(n_2578),
.B2(n_2415),
.Y(n_3315)
);

BUFx6f_ASAP7_75t_L g3316 ( 
.A(n_2963),
.Y(n_3316)
);

INVx2_ASAP7_75t_SL g3317 ( 
.A(n_3031),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3046),
.Y(n_3318)
);

O2A1O1Ixp33_ASAP7_75t_L g3319 ( 
.A1(n_3039),
.A2(n_2943),
.B(n_2589),
.C(n_2635),
.Y(n_3319)
);

BUFx3_ASAP7_75t_L g3320 ( 
.A(n_2999),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3094),
.B(n_3079),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2981),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_3089),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_2985),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2965),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_3089),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2991),
.Y(n_3327)
);

INVx2_ASAP7_75t_SL g3328 ( 
.A(n_2999),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3002),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3149),
.B(n_2695),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2988),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3012),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3020),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3117),
.Y(n_3334)
);

BUFx3_ASAP7_75t_L g3335 ( 
.A(n_2999),
.Y(n_3335)
);

OR2x6_ASAP7_75t_L g3336 ( 
.A(n_2976),
.B(n_2552),
.Y(n_3336)
);

BUFx2_ASAP7_75t_L g3337 ( 
.A(n_3050),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_3134),
.Y(n_3338)
);

CKINVDCx5p33_ASAP7_75t_R g3339 ( 
.A(n_3097),
.Y(n_3339)
);

BUFx2_ASAP7_75t_L g3340 ( 
.A(n_2982),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3028),
.Y(n_3341)
);

INVx2_ASAP7_75t_SL g3342 ( 
.A(n_3015),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3133),
.Y(n_3343)
);

BUFx12f_ASAP7_75t_L g3344 ( 
.A(n_3015),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3181),
.B(n_2701),
.Y(n_3345)
);

AND2x6_ASAP7_75t_L g3346 ( 
.A(n_3112),
.B(n_2389),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_2966),
.A2(n_2919),
.B1(n_2749),
.B2(n_2609),
.Y(n_3347)
);

AND2x4_ASAP7_75t_SL g3348 ( 
.A(n_3015),
.B(n_2686),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3072),
.A2(n_2321),
.B1(n_2578),
.B2(n_2749),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2970),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3073),
.B(n_2702),
.Y(n_3351)
);

BUFx3_ASAP7_75t_L g3352 ( 
.A(n_3001),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3138),
.Y(n_3353)
);

INVx1_ASAP7_75t_SL g3354 ( 
.A(n_3095),
.Y(n_3354)
);

AND2x4_ASAP7_75t_L g3355 ( 
.A(n_3172),
.B(n_2858),
.Y(n_3355)
);

INVxp67_ASAP7_75t_L g3356 ( 
.A(n_3155),
.Y(n_3356)
);

NAND2x1p5_ASAP7_75t_L g3357 ( 
.A(n_3107),
.B(n_2677),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3156),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3163),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3077),
.B(n_2705),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3056),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3014),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3041),
.Y(n_3363)
);

HB1xp67_ASAP7_75t_L g3364 ( 
.A(n_3023),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3171),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3042),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3174),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3044),
.Y(n_3368)
);

INVxp67_ASAP7_75t_SL g3369 ( 
.A(n_2995),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3082),
.B(n_3083),
.Y(n_3370)
);

AND2x4_ASAP7_75t_L g3371 ( 
.A(n_3120),
.B(n_2858),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3088),
.B(n_2717),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3001),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_3003),
.Y(n_3374)
);

INVx2_ASAP7_75t_SL g3375 ( 
.A(n_3010),
.Y(n_3375)
);

INVx4_ASAP7_75t_L g3376 ( 
.A(n_2969),
.Y(n_3376)
);

INVx2_ASAP7_75t_SL g3377 ( 
.A(n_3032),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3060),
.B(n_2966),
.Y(n_3378)
);

BUFx8_ASAP7_75t_L g3379 ( 
.A(n_3099),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3180),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3147),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3081),
.Y(n_3382)
);

INVx5_ASAP7_75t_L g3383 ( 
.A(n_2969),
.Y(n_3383)
);

NOR2xp67_ASAP7_75t_L g3384 ( 
.A(n_3019),
.B(n_2910),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3148),
.Y(n_3385)
);

OR2x6_ASAP7_75t_L g3386 ( 
.A(n_2990),
.B(n_2552),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_3064),
.B(n_2392),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3103),
.B(n_2915),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_SL g3389 ( 
.A(n_2994),
.B(n_2321),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_2967),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3118),
.B(n_2720),
.Y(n_3391)
);

O2A1O1Ixp5_ASAP7_75t_L g3392 ( 
.A1(n_3300),
.A2(n_2995),
.B(n_3023),
.C(n_3017),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_3219),
.B(n_3035),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3362),
.B(n_3068),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3200),
.B(n_3135),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3214),
.A2(n_3122),
.B(n_2975),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_3274),
.A2(n_3055),
.B(n_3137),
.C(n_3173),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3350),
.B(n_3075),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3214),
.A2(n_3017),
.B(n_3136),
.Y(n_3399)
);

OAI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3185),
.A2(n_2972),
.B(n_3177),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3274),
.A2(n_3177),
.B1(n_3006),
.B2(n_2964),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3389),
.A2(n_3153),
.B(n_3136),
.Y(n_3402)
);

AND2x6_ASAP7_75t_SL g3403 ( 
.A(n_3312),
.B(n_3035),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3254),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3363),
.B(n_3366),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3368),
.B(n_3075),
.Y(n_3406)
);

O2A1O1Ixp33_ASAP7_75t_L g3407 ( 
.A1(n_3185),
.A2(n_3301),
.B(n_3308),
.C(n_3272),
.Y(n_3407)
);

AO32x2_ASAP7_75t_L g3408 ( 
.A1(n_3203),
.A2(n_3131),
.A3(n_3110),
.B1(n_3173),
.B2(n_3169),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3200),
.B(n_3040),
.Y(n_3409)
);

O2A1O1Ixp33_ASAP7_75t_L g3410 ( 
.A1(n_3301),
.A2(n_3025),
.B(n_2978),
.C(n_2972),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3389),
.A2(n_3153),
.B(n_2345),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3252),
.A2(n_2345),
.B(n_2535),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_3313),
.B(n_3176),
.Y(n_3413)
);

AOI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3244),
.A2(n_3051),
.B1(n_3048),
.B2(n_3111),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3329),
.B(n_2964),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_3252),
.A2(n_2550),
.B(n_2535),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3272),
.A2(n_2550),
.B(n_2883),
.Y(n_3417)
);

OAI22x1_ASAP7_75t_L g3418 ( 
.A1(n_3340),
.A2(n_3040),
.B1(n_2930),
.B2(n_2589),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_3222),
.B(n_2680),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_3288),
.Y(n_3420)
);

AO221x2_ASAP7_75t_L g3421 ( 
.A1(n_3203),
.A2(n_3169),
.B1(n_3104),
.B2(n_2934),
.C(n_70),
.Y(n_3421)
);

AOI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3300),
.A2(n_2552),
.B(n_2603),
.Y(n_3422)
);

A2O1A1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3308),
.A2(n_3104),
.B(n_3124),
.C(n_3154),
.Y(n_3423)
);

NOR2xp33_ASAP7_75t_L g3424 ( 
.A(n_3313),
.B(n_2685),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3191),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3321),
.B(n_2930),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3332),
.B(n_3124),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3331),
.B(n_3139),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_3188),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3297),
.A2(n_2883),
.B(n_2610),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3210),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3224),
.B(n_3139),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3314),
.B(n_3152),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3297),
.A2(n_2610),
.B(n_2606),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_3251),
.A2(n_2606),
.B(n_2365),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_3251),
.A2(n_2659),
.B(n_2536),
.Y(n_3436)
);

A2O1A1Ixp33_ASAP7_75t_L g3437 ( 
.A1(n_3319),
.A2(n_3096),
.B(n_2659),
.C(n_3129),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3333),
.B(n_3152),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3339),
.B(n_2738),
.Y(n_3439)
);

AOI22x1_ASAP7_75t_L g3440 ( 
.A1(n_3298),
.A2(n_2911),
.B1(n_2918),
.B2(n_2916),
.Y(n_3440)
);

NOR2xp67_ASAP7_75t_SL g3441 ( 
.A(n_3194),
.B(n_2686),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3229),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3225),
.A2(n_2392),
.B(n_2516),
.Y(n_3443)
);

INVx2_ASAP7_75t_SL g3444 ( 
.A(n_3188),
.Y(n_3444)
);

O2A1O1Ixp33_ASAP7_75t_SL g3445 ( 
.A1(n_3330),
.A2(n_3127),
.B(n_3115),
.C(n_2654),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_3312),
.B(n_3195),
.Y(n_3446)
);

NAND2x1p5_ASAP7_75t_L g3447 ( 
.A(n_3222),
.B(n_3261),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_SL g3448 ( 
.A(n_3195),
.B(n_2738),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3257),
.B(n_2578),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3303),
.B(n_3157),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3341),
.B(n_3129),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3225),
.A2(n_2516),
.B(n_2869),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3254),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3327),
.B(n_2919),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_3275),
.B(n_2836),
.Y(n_3455)
);

AOI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3275),
.A2(n_2321),
.B1(n_2919),
.B2(n_2792),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3370),
.A2(n_2871),
.B(n_2869),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3188),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3382),
.B(n_2922),
.Y(n_3459)
);

NOR2xp33_ASAP7_75t_SL g3460 ( 
.A(n_3273),
.B(n_2841),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3375),
.B(n_3067),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3235),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3388),
.B(n_2602),
.Y(n_3463)
);

AOI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3390),
.A2(n_3290),
.B1(n_3269),
.B2(n_3355),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3262),
.B(n_2862),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3228),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3370),
.A2(n_2871),
.B(n_2630),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3228),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3290),
.A2(n_2531),
.B1(n_2522),
.B2(n_2765),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3391),
.A2(n_2654),
.B(n_2647),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3391),
.A2(n_2647),
.B(n_2722),
.Y(n_3471)
);

O2A1O1Ixp33_ASAP7_75t_L g3472 ( 
.A1(n_3319),
.A2(n_2634),
.B(n_2626),
.C(n_2621),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3317),
.B(n_2602),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3223),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_3199),
.B(n_2898),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3239),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3249),
.Y(n_3477)
);

NOR2xp67_ASAP7_75t_L g3478 ( 
.A(n_3311),
.B(n_2945),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3268),
.A2(n_2730),
.B(n_2722),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3310),
.B(n_2927),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3269),
.A2(n_2609),
.B1(n_2796),
.B2(n_2592),
.Y(n_3481)
);

A2O1A1Ixp33_ASAP7_75t_L g3482 ( 
.A1(n_3315),
.A2(n_2928),
.B(n_2944),
.C(n_2933),
.Y(n_3482)
);

NOR3xp33_ASAP7_75t_L g3483 ( 
.A(n_3186),
.B(n_2569),
.C(n_2521),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_3268),
.A2(n_2788),
.B(n_2730),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3192),
.A2(n_2834),
.B1(n_2581),
.B2(n_2597),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3374),
.B(n_3087),
.Y(n_3486)
);

OAI21xp33_ASAP7_75t_SL g3487 ( 
.A1(n_3347),
.A2(n_2890),
.B(n_2920),
.Y(n_3487)
);

AOI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_3355),
.A2(n_2792),
.B1(n_2773),
.B2(n_2764),
.Y(n_3488)
);

OAI21xp33_ASAP7_75t_L g3489 ( 
.A1(n_3387),
.A2(n_2890),
.B(n_2920),
.Y(n_3489)
);

BUFx4f_ASAP7_75t_L g3490 ( 
.A(n_3287),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3322),
.B(n_3324),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3330),
.A2(n_2814),
.B(n_2788),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3347),
.A2(n_2814),
.B(n_2564),
.Y(n_3493)
);

AO21x1_ASAP7_75t_L g3494 ( 
.A1(n_3387),
.A2(n_2931),
.B(n_2924),
.Y(n_3494)
);

INVxp67_ASAP7_75t_L g3495 ( 
.A(n_3337),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_SL g3496 ( 
.A(n_3241),
.B(n_2686),
.Y(n_3496)
);

AO21x2_ASAP7_75t_L g3497 ( 
.A1(n_3349),
.A2(n_2931),
.B(n_2924),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3183),
.Y(n_3498)
);

INVx3_ASAP7_75t_L g3499 ( 
.A(n_3287),
.Y(n_3499)
);

BUFx8_ASAP7_75t_L g3500 ( 
.A(n_3187),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3381),
.B(n_2734),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_SL g3502 ( 
.A1(n_3292),
.A2(n_2894),
.B(n_2529),
.C(n_2524),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3385),
.B(n_2736),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3369),
.A2(n_2894),
.B(n_2509),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3298),
.B(n_2737),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3369),
.A2(n_2509),
.B(n_2538),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_3306),
.A2(n_2538),
.B(n_2367),
.Y(n_3507)
);

INVxp67_ASAP7_75t_SL g3508 ( 
.A(n_3276),
.Y(n_3508)
);

AO32x2_ASAP7_75t_L g3509 ( 
.A1(n_3377),
.A2(n_2617),
.A3(n_2503),
.B1(n_2819),
.B2(n_2812),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_3354),
.B(n_2740),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3227),
.B(n_2796),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3325),
.B(n_2743),
.Y(n_3512)
);

A2O1A1Ixp33_ASAP7_75t_L g3513 ( 
.A1(n_3378),
.A2(n_2573),
.B(n_2548),
.C(n_2452),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3354),
.B(n_2746),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3306),
.A2(n_2529),
.B(n_2524),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3197),
.B(n_2750),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3345),
.A2(n_2463),
.B(n_2462),
.Y(n_3517)
);

BUFx4f_ASAP7_75t_L g3518 ( 
.A(n_3287),
.Y(n_3518)
);

NAND3xp33_ASAP7_75t_L g3519 ( 
.A(n_3264),
.B(n_2614),
.C(n_2867),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3193),
.B(n_2752),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3345),
.A2(n_2463),
.B(n_2462),
.Y(n_3521)
);

O2A1O1Ixp33_ASAP7_75t_SL g3522 ( 
.A1(n_3292),
.A2(n_2983),
.B(n_2757),
.C(n_2766),
.Y(n_3522)
);

BUFx6f_ASAP7_75t_L g3523 ( 
.A(n_3211),
.Y(n_3523)
);

A2O1A1Ixp33_ASAP7_75t_L g3524 ( 
.A1(n_3378),
.A2(n_2568),
.B(n_2588),
.C(n_2585),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3199),
.B(n_2773),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3193),
.B(n_3318),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3232),
.A2(n_2609),
.B1(n_2530),
.B2(n_2590),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3201),
.B(n_2688),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3201),
.B(n_3285),
.Y(n_3529)
);

OAI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3212),
.A2(n_2834),
.B1(n_2329),
.B2(n_2333),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3212),
.A2(n_2336),
.B1(n_2344),
.B2(n_2326),
.Y(n_3531)
);

BUFx2_ASAP7_75t_L g3532 ( 
.A(n_3302),
.Y(n_3532)
);

OA22x2_ASAP7_75t_L g3533 ( 
.A1(n_3234),
.A2(n_2877),
.B1(n_2879),
.B2(n_2876),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3358),
.B(n_2753),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3184),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3294),
.A2(n_2463),
.B(n_2462),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3359),
.B(n_2779),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3384),
.B(n_2787),
.Y(n_3538)
);

OAI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_3286),
.A2(n_3356),
.B1(n_3216),
.B2(n_3238),
.Y(n_3539)
);

OAI21xp33_ASAP7_75t_SL g3540 ( 
.A1(n_3255),
.A2(n_2811),
.B(n_2790),
.Y(n_3540)
);

INVx2_ASAP7_75t_SL g3541 ( 
.A(n_3211),
.Y(n_3541)
);

BUFx6f_ASAP7_75t_L g3542 ( 
.A(n_3211),
.Y(n_3542)
);

BUFx12f_ASAP7_75t_L g3543 ( 
.A(n_3323),
.Y(n_3543)
);

CKINVDCx10_ASAP7_75t_R g3544 ( 
.A(n_3207),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3356),
.B(n_2820),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3294),
.A2(n_2731),
.B(n_2677),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3255),
.A2(n_3221),
.B(n_3351),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3380),
.B(n_2904),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3334),
.B(n_2885),
.Y(n_3549)
);

OAI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_3286),
.A2(n_2348),
.B1(n_2362),
.B2(n_2346),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3343),
.B(n_2892),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3221),
.A2(n_2733),
.B(n_2731),
.Y(n_3552)
);

AOI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3336),
.A2(n_2401),
.B(n_2400),
.Y(n_3553)
);

BUFx10_ASAP7_75t_L g3554 ( 
.A(n_3326),
.Y(n_3554)
);

NAND2xp33_ASAP7_75t_L g3555 ( 
.A(n_3316),
.B(n_2688),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_L g3556 ( 
.A(n_3265),
.B(n_2688),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3372),
.A2(n_2401),
.B(n_2400),
.Y(n_3557)
);

O2A1O1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3276),
.A2(n_2500),
.B(n_2368),
.C(n_2376),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3353),
.B(n_2893),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_SL g3560 ( 
.A(n_3371),
.B(n_2724),
.Y(n_3560)
);

AO32x2_ASAP7_75t_L g3561 ( 
.A1(n_3328),
.A2(n_2503),
.A3(n_2866),
.B1(n_2819),
.B2(n_2812),
.Y(n_3561)
);

O2A1O1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_3196),
.A2(n_2378),
.B(n_2363),
.C(n_2584),
.Y(n_3562)
);

BUFx8_ASAP7_75t_L g3563 ( 
.A(n_3316),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_3351),
.A2(n_2745),
.B(n_2733),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3365),
.B(n_3367),
.Y(n_3565)
);

AO21x1_ASAP7_75t_L g3566 ( 
.A1(n_3372),
.A2(n_3360),
.B(n_3357),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3246),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3386),
.A2(n_2874),
.B1(n_2313),
.B2(n_2322),
.Y(n_3568)
);

NOR2x1_ASAP7_75t_R g3569 ( 
.A(n_3222),
.B(n_2693),
.Y(n_3569)
);

BUFx3_ASAP7_75t_L g3570 ( 
.A(n_3237),
.Y(n_3570)
);

AOI21x1_ASAP7_75t_L g3571 ( 
.A1(n_3336),
.A2(n_2418),
.B(n_2398),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3189),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3386),
.A2(n_2874),
.B1(n_2693),
.B2(n_2315),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3196),
.B(n_2829),
.Y(n_3574)
);

AOI33xp33_ASAP7_75t_L g3575 ( 
.A1(n_3361),
.A2(n_92),
.A3(n_76),
.B1(n_100),
.B2(n_84),
.B3(n_68),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3360),
.A2(n_2758),
.B(n_2745),
.Y(n_3576)
);

O2A1O1Ixp33_ASAP7_75t_L g3577 ( 
.A1(n_3247),
.A2(n_2315),
.B(n_2946),
.C(n_2437),
.Y(n_3577)
);

BUFx2_ASAP7_75t_L g3578 ( 
.A(n_3379),
.Y(n_3578)
);

OAI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3357),
.A2(n_2449),
.B(n_2436),
.Y(n_3579)
);

AOI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3271),
.A2(n_2724),
.B1(n_2530),
.B2(n_2609),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_L g3581 ( 
.A(n_3202),
.B(n_2693),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3371),
.B(n_2971),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3263),
.B(n_2830),
.Y(n_3583)
);

BUFx6f_ASAP7_75t_L g3584 ( 
.A(n_3289),
.Y(n_3584)
);

NAND2x1p5_ASAP7_75t_L g3585 ( 
.A(n_3222),
.B(n_3261),
.Y(n_3585)
);

A2O1A1Ixp33_ASAP7_75t_L g3586 ( 
.A1(n_3190),
.A2(n_2801),
.B(n_2777),
.C(n_2758),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3386),
.A2(n_2801),
.B1(n_2802),
.B2(n_2777),
.Y(n_3587)
);

NOR2xp67_ASAP7_75t_L g3588 ( 
.A(n_3364),
.B(n_2971),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3284),
.A2(n_2810),
.B(n_2802),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3271),
.A2(n_2530),
.B1(n_2609),
.B2(n_2900),
.Y(n_3590)
);

OAI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3336),
.A2(n_2810),
.B1(n_2374),
.B2(n_2377),
.Y(n_3591)
);

NOR2xp67_ASAP7_75t_SL g3592 ( 
.A(n_3261),
.B(n_3344),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3198),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3267),
.B(n_2843),
.Y(n_3594)
);

BUFx6f_ASAP7_75t_L g3595 ( 
.A(n_3289),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3277),
.B(n_2847),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3278),
.B(n_2870),
.Y(n_3597)
);

BUFx3_ASAP7_75t_L g3598 ( 
.A(n_3218),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3280),
.B(n_2872),
.Y(n_3599)
);

INVxp67_ASAP7_75t_L g3600 ( 
.A(n_3258),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3284),
.A2(n_2534),
.B(n_2465),
.Y(n_3601)
);

AND2x2_ASAP7_75t_SL g3602 ( 
.A(n_3206),
.B(n_2866),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3364),
.A2(n_3346),
.B1(n_3291),
.B2(n_3202),
.Y(n_3603)
);

AOI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3230),
.A2(n_2609),
.B1(n_2900),
.B2(n_2590),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_3584),
.Y(n_3605)
);

NOR3xp33_ASAP7_75t_L g3606 ( 
.A(n_3407),
.B(n_3342),
.C(n_3213),
.Y(n_3606)
);

OA21x2_ASAP7_75t_L g3607 ( 
.A1(n_3400),
.A2(n_3243),
.B(n_3240),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3404),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3396),
.A2(n_3245),
.B(n_3236),
.Y(n_3609)
);

INVx1_ASAP7_75t_SL g3610 ( 
.A(n_3448),
.Y(n_3610)
);

OAI21x1_ASAP7_75t_L g3611 ( 
.A1(n_3571),
.A2(n_3236),
.B(n_3208),
.Y(n_3611)
);

OAI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3397),
.A2(n_3346),
.B(n_3291),
.Y(n_3612)
);

OAI21x1_ASAP7_75t_L g3613 ( 
.A1(n_3422),
.A2(n_3209),
.B(n_3204),
.Y(n_3613)
);

OAI21x1_ASAP7_75t_L g3614 ( 
.A1(n_3506),
.A2(n_3220),
.B(n_3215),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_3511),
.B(n_3226),
.Y(n_3615)
);

INVx3_ASAP7_75t_L g3616 ( 
.A(n_3584),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3436),
.A2(n_3284),
.B(n_3383),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3401),
.A2(n_3233),
.B1(n_3261),
.B2(n_3281),
.Y(n_3618)
);

AOI21xp33_ASAP7_75t_L g3619 ( 
.A1(n_3410),
.A2(n_3296),
.B(n_3283),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3426),
.B(n_3230),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3453),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3526),
.B(n_3299),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3466),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3553),
.A2(n_2828),
.B(n_2825),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3557),
.A2(n_3507),
.B(n_3417),
.Y(n_3625)
);

A2O1A1Ixp33_ASAP7_75t_L g3626 ( 
.A1(n_3437),
.A2(n_3320),
.B(n_3335),
.C(n_3348),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3393),
.A2(n_3346),
.B(n_3291),
.Y(n_3627)
);

O2A1O1Ixp5_ASAP7_75t_SL g3628 ( 
.A1(n_3446),
.A2(n_3205),
.B(n_3217),
.C(n_3182),
.Y(n_3628)
);

NOR3xp33_ASAP7_75t_L g3629 ( 
.A(n_3539),
.B(n_3213),
.C(n_3206),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3508),
.B(n_3250),
.Y(n_3630)
);

BUFx4_ASAP7_75t_SL g3631 ( 
.A(n_3578),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_3478),
.B(n_3250),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3504),
.A2(n_2828),
.B(n_2825),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3532),
.B(n_3432),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3522),
.A2(n_3383),
.B(n_3376),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3477),
.Y(n_3636)
);

BUFx3_ASAP7_75t_L g3637 ( 
.A(n_3474),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3547),
.B(n_3253),
.Y(n_3638)
);

OAI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3423),
.A2(n_3259),
.B1(n_3270),
.B2(n_3260),
.Y(n_3639)
);

AND2x4_ASAP7_75t_L g3640 ( 
.A(n_3468),
.B(n_3182),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3445),
.A2(n_3399),
.B(n_3467),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3584),
.Y(n_3642)
);

INVx2_ASAP7_75t_SL g3643 ( 
.A(n_3429),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3565),
.B(n_3307),
.Y(n_3644)
);

NOR2x1_ASAP7_75t_SL g3645 ( 
.A(n_3587),
.B(n_3383),
.Y(n_3645)
);

INVx1_ASAP7_75t_SL g3646 ( 
.A(n_3420),
.Y(n_3646)
);

AO32x2_ASAP7_75t_L g3647 ( 
.A1(n_3591),
.A2(n_3293),
.A3(n_3282),
.B1(n_3376),
.B2(n_3291),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3411),
.A2(n_3383),
.B(n_2476),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3601),
.A2(n_3373),
.B(n_3027),
.Y(n_3649)
);

INVx2_ASAP7_75t_SL g3650 ( 
.A(n_3429),
.Y(n_3650)
);

OAI21x1_ASAP7_75t_L g3651 ( 
.A1(n_3471),
.A2(n_3027),
.B(n_2979),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3500),
.Y(n_3652)
);

O2A1O1Ixp5_ASAP7_75t_SL g3653 ( 
.A1(n_3409),
.A2(n_3217),
.B(n_3231),
.C(n_3205),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3412),
.A2(n_2464),
.B(n_2979),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3430),
.A2(n_3434),
.B(n_3492),
.Y(n_3655)
);

AOI21xp33_ASAP7_75t_L g3656 ( 
.A1(n_3489),
.A2(n_3279),
.B(n_3379),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3540),
.A2(n_3091),
.B(n_3059),
.Y(n_3657)
);

AO31x2_ASAP7_75t_L g3658 ( 
.A1(n_3494),
.A2(n_2503),
.A3(n_2929),
.B(n_2926),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3552),
.A2(n_3470),
.B(n_3546),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3487),
.A2(n_3346),
.B(n_3291),
.Y(n_3660)
);

OAI21x1_ASAP7_75t_L g3661 ( 
.A1(n_3564),
.A2(n_3091),
.B(n_3059),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3575),
.A2(n_3295),
.B(n_3352),
.C(n_3305),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3398),
.B(n_3346),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3406),
.B(n_3266),
.Y(n_3664)
);

XOR2xp5_ASAP7_75t_L g3665 ( 
.A(n_3488),
.B(n_3295),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3413),
.B(n_3304),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3502),
.A2(n_3116),
.B(n_3113),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3576),
.A2(n_3116),
.B(n_3113),
.Y(n_3668)
);

OAI21x1_ASAP7_75t_SL g3669 ( 
.A1(n_3566),
.A2(n_2941),
.B(n_2932),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3498),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3416),
.A2(n_3338),
.B(n_3309),
.Y(n_3671)
);

INVx4_ASAP7_75t_L g3672 ( 
.A(n_3595),
.Y(n_3672)
);

OAI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3435),
.A2(n_3242),
.B(n_3231),
.Y(n_3673)
);

HB1xp67_ASAP7_75t_L g3674 ( 
.A(n_3588),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3491),
.B(n_3242),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3405),
.B(n_3248),
.Y(n_3676)
);

AO31x2_ASAP7_75t_L g3677 ( 
.A1(n_3418),
.A2(n_2949),
.A3(n_2954),
.B(n_2950),
.Y(n_3677)
);

OAI21x1_ASAP7_75t_L g3678 ( 
.A1(n_3536),
.A2(n_3256),
.B(n_3248),
.Y(n_3678)
);

NAND2x1_ASAP7_75t_L g3679 ( 
.A(n_3592),
.B(n_3304),
.Y(n_3679)
);

OAI21xp5_ASAP7_75t_L g3680 ( 
.A1(n_3472),
.A2(n_2590),
.B(n_2540),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3429),
.Y(n_3681)
);

OAI21x1_ASAP7_75t_L g3682 ( 
.A1(n_3517),
.A2(n_3266),
.B(n_3256),
.Y(n_3682)
);

OAI21x1_ASAP7_75t_L g3683 ( 
.A1(n_3521),
.A2(n_2946),
.B(n_2523),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3433),
.B(n_3289),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3500),
.Y(n_3685)
);

OA21x2_ASAP7_75t_L g3686 ( 
.A1(n_3392),
.A2(n_2896),
.B(n_2956),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3535),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3395),
.B(n_3316),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3394),
.B(n_3305),
.Y(n_3689)
);

BUFx3_ASAP7_75t_L g3690 ( 
.A(n_3570),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3424),
.B(n_3455),
.Y(n_3691)
);

A2O1A1Ixp33_ASAP7_75t_L g3692 ( 
.A1(n_3414),
.A2(n_3338),
.B(n_3309),
.C(n_2868),
.Y(n_3692)
);

BUFx8_ASAP7_75t_L g3693 ( 
.A(n_3543),
.Y(n_3693)
);

OAI21x1_ASAP7_75t_L g3694 ( 
.A1(n_3493),
.A2(n_3515),
.B(n_3457),
.Y(n_3694)
);

BUFx2_ASAP7_75t_L g3695 ( 
.A(n_3563),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3460),
.B(n_189),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3569),
.A2(n_2361),
.B(n_2311),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3469),
.A2(n_2590),
.B(n_2540),
.Y(n_3698)
);

AND2x4_ASAP7_75t_L g3699 ( 
.A(n_3588),
.B(n_2842),
.Y(n_3699)
);

OAI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3440),
.A2(n_2523),
.B(n_2505),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3520),
.B(n_190),
.Y(n_3701)
);

INVx3_ASAP7_75t_L g3702 ( 
.A(n_3595),
.Y(n_3702)
);

OAI21x1_ASAP7_75t_L g3703 ( 
.A1(n_3479),
.A2(n_2523),
.B(n_2505),
.Y(n_3703)
);

INVxp67_ASAP7_75t_L g3704 ( 
.A(n_3598),
.Y(n_3704)
);

OAI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3519),
.A2(n_2590),
.B(n_2540),
.Y(n_3705)
);

OAI21x1_ASAP7_75t_L g3706 ( 
.A1(n_3484),
.A2(n_2525),
.B(n_2505),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3572),
.B(n_2540),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3505),
.B(n_190),
.Y(n_3708)
);

AOI21x1_ASAP7_75t_SL g3709 ( 
.A1(n_3454),
.A2(n_2528),
.B(n_192),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_3439),
.B(n_2710),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3415),
.B(n_191),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3593),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3569),
.A2(n_2361),
.B(n_2311),
.Y(n_3713)
);

OA22x2_ASAP7_75t_L g3714 ( 
.A1(n_3464),
.A2(n_2868),
.B1(n_2881),
.B2(n_2842),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_SL g3715 ( 
.A(n_3602),
.B(n_2710),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_3475),
.B(n_191),
.Y(n_3716)
);

AND2x4_ASAP7_75t_L g3717 ( 
.A(n_3495),
.B(n_2881),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3465),
.B(n_3403),
.Y(n_3718)
);

INVx2_ASAP7_75t_SL g3719 ( 
.A(n_3458),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3427),
.B(n_192),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3516),
.B(n_193),
.Y(n_3721)
);

AO21x1_ASAP7_75t_L g3722 ( 
.A1(n_3510),
.A2(n_3450),
.B(n_3503),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3425),
.B(n_193),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3533),
.Y(n_3724)
);

BUFx2_ASAP7_75t_L g3725 ( 
.A(n_3563),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3431),
.B(n_194),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3419),
.B(n_2710),
.Y(n_3727)
);

OAI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3482),
.A2(n_2590),
.B(n_2540),
.Y(n_3728)
);

A2O1A1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_3456),
.A2(n_2377),
.B(n_2374),
.C(n_2525),
.Y(n_3729)
);

OAI21x1_ASAP7_75t_L g3730 ( 
.A1(n_3402),
.A2(n_2525),
.B(n_2461),
.Y(n_3730)
);

BUFx6f_ASAP7_75t_L g3731 ( 
.A(n_3458),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3442),
.B(n_196),
.Y(n_3732)
);

AOI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3538),
.A2(n_3486),
.B(n_3461),
.Y(n_3733)
);

AND3x4_ASAP7_75t_L g3734 ( 
.A(n_3544),
.B(n_69),
.C(n_70),
.Y(n_3734)
);

AOI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3568),
.A2(n_2361),
.B(n_2540),
.Y(n_3735)
);

A2O1A1Ixp33_ASAP7_75t_L g3736 ( 
.A1(n_3481),
.A2(n_2377),
.B(n_2461),
.C(n_2721),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3462),
.Y(n_3737)
);

OAI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3513),
.A2(n_2838),
.B(n_2815),
.Y(n_3738)
);

AOI21xp33_ASAP7_75t_L g3739 ( 
.A1(n_3497),
.A2(n_3577),
.B(n_3558),
.Y(n_3739)
);

A2O1A1Ixp33_ASAP7_75t_L g3740 ( 
.A1(n_3604),
.A2(n_2461),
.B(n_2728),
.C(n_2721),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3476),
.B(n_196),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3567),
.B(n_197),
.Y(n_3742)
);

OAI21xp33_ASAP7_75t_L g3743 ( 
.A1(n_3451),
.A2(n_70),
.B(n_71),
.Y(n_3743)
);

OAI21x1_ASAP7_75t_L g3744 ( 
.A1(n_3589),
.A2(n_3443),
.B(n_3452),
.Y(n_3744)
);

CKINVDCx5p33_ASAP7_75t_R g3745 ( 
.A(n_3554),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3514),
.B(n_197),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3586),
.A2(n_2728),
.B(n_2721),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3497),
.A2(n_2816),
.B(n_2728),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_SL g3749 ( 
.A1(n_3524),
.A2(n_2856),
.B(n_2816),
.Y(n_3749)
);

OAI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3483),
.A2(n_2838),
.B(n_2815),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3545),
.B(n_198),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3574),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3447),
.A2(n_2838),
.B(n_2815),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3548),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3512),
.Y(n_3755)
);

OAI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3585),
.A2(n_2838),
.B(n_2815),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3579),
.A2(n_2884),
.B(n_2865),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3473),
.Y(n_3758)
);

BUFx2_ASAP7_75t_L g3759 ( 
.A(n_3499),
.Y(n_3759)
);

AOI221x1_ASAP7_75t_L g3760 ( 
.A1(n_3485),
.A2(n_2856),
.B1(n_2816),
.B2(n_2861),
.C(n_73),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3421),
.A2(n_2861),
.B(n_2856),
.Y(n_3761)
);

OAI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_3562),
.A2(n_2884),
.B(n_2865),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3421),
.A2(n_2861),
.B(n_2884),
.Y(n_3763)
);

OAI21x1_ASAP7_75t_L g3764 ( 
.A1(n_3603),
.A2(n_2884),
.B(n_2865),
.Y(n_3764)
);

AOI31xp67_ASAP7_75t_L g3765 ( 
.A1(n_3590),
.A2(n_2888),
.A3(n_2865),
.B(n_73),
.Y(n_3765)
);

AO22x2_ASAP7_75t_L g3766 ( 
.A1(n_3573),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3428),
.B(n_199),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3438),
.B(n_199),
.Y(n_3768)
);

OAI21xp33_ASAP7_75t_L g3769 ( 
.A1(n_3459),
.A2(n_71),
.B(n_72),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3449),
.B(n_200),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3480),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3582),
.A2(n_2888),
.B(n_72),
.Y(n_3772)
);

BUFx3_ASAP7_75t_L g3773 ( 
.A(n_3458),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_3419),
.B(n_2888),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3501),
.B(n_200),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3534),
.A2(n_2888),
.B(n_74),
.Y(n_3776)
);

INVx3_ASAP7_75t_L g3777 ( 
.A(n_3595),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3537),
.A2(n_74),
.B(n_75),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3549),
.B(n_201),
.Y(n_3779)
);

OAI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3531),
.A2(n_82),
.B(n_74),
.Y(n_3780)
);

AND2x6_ASAP7_75t_L g3781 ( 
.A(n_3580),
.B(n_75),
.Y(n_3781)
);

A2O1A1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_3529),
.A2(n_203),
.B(n_205),
.C(n_202),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3551),
.B(n_205),
.Y(n_3783)
);

OAI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3550),
.A2(n_83),
.B(n_75),
.Y(n_3784)
);

AOI211x1_ASAP7_75t_L g3785 ( 
.A1(n_3441),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3559),
.B(n_208),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3530),
.A2(n_3555),
.B(n_3560),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3463),
.B(n_208),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3527),
.A2(n_77),
.B(n_79),
.Y(n_3789)
);

OAI21x1_ASAP7_75t_L g3790 ( 
.A1(n_3583),
.A2(n_77),
.B(n_79),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3490),
.A2(n_79),
.B(n_80),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3594),
.B(n_3596),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3528),
.B(n_209),
.Y(n_3793)
);

OAI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3597),
.A2(n_80),
.B(n_81),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3525),
.B(n_209),
.Y(n_3795)
);

AO21x2_ASAP7_75t_L g3796 ( 
.A1(n_3599),
.A2(n_80),
.B(n_81),
.Y(n_3796)
);

CKINVDCx5p33_ASAP7_75t_R g3797 ( 
.A(n_3554),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3499),
.A2(n_82),
.B(n_83),
.Y(n_3798)
);

CKINVDCx5p33_ASAP7_75t_R g3799 ( 
.A(n_3523),
.Y(n_3799)
);

INVx5_ASAP7_75t_L g3800 ( 
.A(n_3523),
.Y(n_3800)
);

INVx1_ASAP7_75t_SL g3801 ( 
.A(n_3523),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3600),
.B(n_211),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3581),
.A2(n_82),
.B(n_84),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3408),
.B(n_692),
.Y(n_3804)
);

OAI21x1_ASAP7_75t_L g3805 ( 
.A1(n_3509),
.A2(n_84),
.B(n_85),
.Y(n_3805)
);

OA21x2_ASAP7_75t_L g3806 ( 
.A1(n_3509),
.A2(n_3556),
.B(n_3408),
.Y(n_3806)
);

OAI21xp33_ASAP7_75t_L g3807 ( 
.A1(n_3496),
.A2(n_85),
.B(n_86),
.Y(n_3807)
);

NOR2xp67_ASAP7_75t_L g3808 ( 
.A(n_3444),
.B(n_85),
.Y(n_3808)
);

BUFx3_ASAP7_75t_L g3809 ( 
.A(n_3542),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3541),
.B(n_211),
.Y(n_3810)
);

INVx5_ASAP7_75t_L g3811 ( 
.A(n_3542),
.Y(n_3811)
);

AOI21x1_ASAP7_75t_SL g3812 ( 
.A1(n_3490),
.A2(n_213),
.B(n_212),
.Y(n_3812)
);

NOR2xp33_ASAP7_75t_L g3813 ( 
.A(n_3542),
.B(n_212),
.Y(n_3813)
);

OAI21xp5_ASAP7_75t_L g3814 ( 
.A1(n_3518),
.A2(n_86),
.B(n_87),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3518),
.A2(n_86),
.B(n_87),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_L g3816 ( 
.A1(n_3408),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3816)
);

INVx3_ASAP7_75t_L g3817 ( 
.A(n_3561),
.Y(n_3817)
);

OAI21x1_ASAP7_75t_L g3818 ( 
.A1(n_3509),
.A2(n_88),
.B(n_89),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3561),
.B(n_213),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3561),
.B(n_88),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3526),
.B(n_215),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_SL g3822 ( 
.A1(n_3397),
.A2(n_90),
.B(n_91),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3526),
.B(n_215),
.Y(n_3823)
);

NAND2x1_ASAP7_75t_L g3824 ( 
.A(n_3592),
.B(n_216),
.Y(n_3824)
);

OR2x6_ASAP7_75t_L g3825 ( 
.A(n_3399),
.B(n_217),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3526),
.B(n_217),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3511),
.B(n_692),
.Y(n_3827)
);

HB1xp67_ASAP7_75t_L g3828 ( 
.A(n_3420),
.Y(n_3828)
);

AOI21xp33_ASAP7_75t_L g3829 ( 
.A1(n_3407),
.A2(n_90),
.B(n_91),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3404),
.Y(n_3830)
);

NOR2x1_ASAP7_75t_L g3831 ( 
.A(n_3448),
.B(n_218),
.Y(n_3831)
);

OAI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3396),
.A2(n_92),
.B(n_93),
.Y(n_3832)
);

OAI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3400),
.A2(n_92),
.B(n_93),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3728),
.A2(n_93),
.B(n_94),
.Y(n_3834)
);

A2O1A1Ixp33_ASAP7_75t_L g3835 ( 
.A1(n_3833),
.A2(n_219),
.B(n_220),
.C(n_218),
.Y(n_3835)
);

O2A1O1Ixp33_ASAP7_75t_L g3836 ( 
.A1(n_3782),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_3836)
);

AOI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3728),
.A2(n_94),
.B(n_96),
.Y(n_3837)
);

OAI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3833),
.A2(n_96),
.B(n_97),
.Y(n_3838)
);

AOI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3820),
.A2(n_97),
.B(n_98),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3636),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3752),
.B(n_220),
.Y(n_3841)
);

OAI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3791),
.A2(n_3815),
.B(n_3829),
.Y(n_3842)
);

NOR2x1_ASAP7_75t_L g3843 ( 
.A(n_3749),
.B(n_97),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3687),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3641),
.A2(n_98),
.B(n_99),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3670),
.Y(n_3846)
);

O2A1O1Ixp33_ASAP7_75t_L g3847 ( 
.A1(n_3829),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_3847)
);

AO31x2_ASAP7_75t_L g3848 ( 
.A1(n_3617),
.A2(n_102),
.A3(n_99),
.B(n_101),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3712),
.Y(n_3849)
);

NAND2x1_ASAP7_75t_L g3850 ( 
.A(n_3607),
.B(n_221),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3674),
.B(n_3828),
.Y(n_3851)
);

INVx3_ASAP7_75t_L g3852 ( 
.A(n_3637),
.Y(n_3852)
);

OAI21x1_ASAP7_75t_L g3853 ( 
.A1(n_3625),
.A2(n_102),
.B(n_103),
.Y(n_3853)
);

INVx3_ASAP7_75t_L g3854 ( 
.A(n_3690),
.Y(n_3854)
);

AOI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_3680),
.A2(n_3698),
.B(n_3635),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3680),
.A2(n_102),
.B(n_103),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_SL g3857 ( 
.A(n_3745),
.B(n_3797),
.Y(n_3857)
);

A2O1A1Ixp33_ASAP7_75t_L g3858 ( 
.A1(n_3807),
.A2(n_222),
.B(n_223),
.C(n_221),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3659),
.A2(n_104),
.B(n_105),
.Y(n_3859)
);

INVx3_ASAP7_75t_L g3860 ( 
.A(n_3731),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3698),
.A2(n_104),
.B(n_105),
.Y(n_3861)
);

AO32x2_ASAP7_75t_L g3862 ( 
.A1(n_3618),
.A2(n_106),
.A3(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_3862)
);

AO31x2_ASAP7_75t_L g3863 ( 
.A1(n_3722),
.A2(n_109),
.A3(n_106),
.B(n_107),
.Y(n_3863)
);

O2A1O1Ixp5_ASAP7_75t_L g3864 ( 
.A1(n_3814),
.A2(n_110),
.B(n_107),
.C(n_109),
.Y(n_3864)
);

AO21x1_ASAP7_75t_L g3865 ( 
.A1(n_3820),
.A2(n_110),
.B(n_111),
.Y(n_3865)
);

AOI21x1_ASAP7_75t_L g3866 ( 
.A1(n_3819),
.A2(n_111),
.B(n_112),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3705),
.A2(n_112),
.B(n_113),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3646),
.B(n_224),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3634),
.B(n_224),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3608),
.Y(n_3870)
);

A2O1A1Ixp33_ASAP7_75t_L g3871 ( 
.A1(n_3807),
.A2(n_3743),
.B(n_3769),
.C(n_3814),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3621),
.Y(n_3872)
);

HB1xp67_ASAP7_75t_L g3873 ( 
.A(n_3646),
.Y(n_3873)
);

O2A1O1Ixp33_ASAP7_75t_L g3874 ( 
.A1(n_3743),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3816),
.A2(n_3662),
.B1(n_3825),
.B2(n_3626),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3830),
.Y(n_3876)
);

AND2x6_ASAP7_75t_SL g3877 ( 
.A(n_3718),
.B(n_3716),
.Y(n_3877)
);

A2O1A1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_3769),
.A2(n_3784),
.B(n_3780),
.C(n_3696),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3771),
.B(n_225),
.Y(n_3879)
);

AO31x2_ASAP7_75t_L g3880 ( 
.A1(n_3645),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_3880)
);

OAI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3744),
.A2(n_114),
.B(n_115),
.Y(n_3881)
);

INVx1_ASAP7_75t_SL g3882 ( 
.A(n_3631),
.Y(n_3882)
);

BUFx2_ASAP7_75t_L g3883 ( 
.A(n_3759),
.Y(n_3883)
);

OAI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3778),
.A2(n_115),
.B(n_116),
.Y(n_3884)
);

OAI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3776),
.A2(n_116),
.B(n_117),
.Y(n_3885)
);

HB1xp67_ASAP7_75t_L g3886 ( 
.A(n_3607),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3623),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3737),
.Y(n_3888)
);

O2A1O1Ixp33_ASAP7_75t_L g3889 ( 
.A1(n_3780),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_3889)
);

INVx2_ASAP7_75t_SL g3890 ( 
.A(n_3799),
.Y(n_3890)
);

INVxp67_ASAP7_75t_L g3891 ( 
.A(n_3691),
.Y(n_3891)
);

OAI21x1_ASAP7_75t_L g3892 ( 
.A1(n_3655),
.A2(n_117),
.B(n_118),
.Y(n_3892)
);

AO31x2_ASAP7_75t_L g3893 ( 
.A1(n_3760),
.A2(n_120),
.A3(n_118),
.B(n_119),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3705),
.A2(n_119),
.B(n_120),
.Y(n_3894)
);

AOI221x1_ASAP7_75t_L g3895 ( 
.A1(n_3766),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3614),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3613),
.Y(n_3897)
);

O2A1O1Ixp33_ASAP7_75t_L g3898 ( 
.A1(n_3784),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_3898)
);

AO31x2_ASAP7_75t_L g3899 ( 
.A1(n_3618),
.A2(n_125),
.A3(n_121),
.B(n_124),
.Y(n_3899)
);

OAI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_3825),
.A2(n_124),
.B(n_125),
.Y(n_3900)
);

BUFx6f_ASAP7_75t_L g3901 ( 
.A(n_3731),
.Y(n_3901)
);

AOI21x1_ASAP7_75t_L g3902 ( 
.A1(n_3679),
.A2(n_124),
.B(n_125),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3663),
.B(n_225),
.Y(n_3903)
);

NOR2xp33_ASAP7_75t_L g3904 ( 
.A(n_3610),
.B(n_3666),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3638),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3755),
.B(n_226),
.Y(n_3906)
);

BUFx6f_ASAP7_75t_L g3907 ( 
.A(n_3731),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3758),
.Y(n_3908)
);

BUFx10_ASAP7_75t_L g3909 ( 
.A(n_3813),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3694),
.A2(n_126),
.B(n_127),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3754),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3825),
.A2(n_126),
.B(n_128),
.Y(n_3912)
);

OAI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3787),
.A2(n_126),
.B(n_128),
.Y(n_3913)
);

AOI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_3648),
.A2(n_129),
.B(n_130),
.Y(n_3914)
);

AND2x4_ASAP7_75t_L g3915 ( 
.A(n_3640),
.B(n_226),
.Y(n_3915)
);

BUFx3_ASAP7_75t_L g3916 ( 
.A(n_3693),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3610),
.B(n_228),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3612),
.A2(n_129),
.B(n_130),
.Y(n_3918)
);

BUFx12f_ASAP7_75t_L g3919 ( 
.A(n_3693),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_3688),
.B(n_229),
.Y(n_3920)
);

AO31x2_ASAP7_75t_L g3921 ( 
.A1(n_3740),
.A2(n_132),
.A3(n_129),
.B(n_131),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3664),
.B(n_230),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3689),
.B(n_230),
.Y(n_3923)
);

BUFx12f_ASAP7_75t_L g3924 ( 
.A(n_3652),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3789),
.A2(n_232),
.B(n_233),
.C(n_231),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3612),
.A2(n_131),
.B(n_132),
.Y(n_3926)
);

NOR2xp67_ASAP7_75t_L g3927 ( 
.A(n_3704),
.B(n_3817),
.Y(n_3927)
);

INVx4_ASAP7_75t_L g3928 ( 
.A(n_3605),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3640),
.Y(n_3929)
);

INVx3_ASAP7_75t_L g3930 ( 
.A(n_3773),
.Y(n_3930)
);

OR2x2_ASAP7_75t_L g3931 ( 
.A(n_3615),
.B(n_233),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3735),
.A2(n_131),
.B(n_132),
.Y(n_3932)
);

OAI21x1_ASAP7_75t_L g3933 ( 
.A1(n_3669),
.A2(n_133),
.B(n_134),
.Y(n_3933)
);

BUFx6f_ASAP7_75t_L g3934 ( 
.A(n_3809),
.Y(n_3934)
);

OAI21x1_ASAP7_75t_L g3935 ( 
.A1(n_3703),
.A2(n_133),
.B(n_134),
.Y(n_3935)
);

OR2x2_ASAP7_75t_L g3936 ( 
.A(n_3644),
.B(n_234),
.Y(n_3936)
);

BUFx10_ASAP7_75t_L g3937 ( 
.A(n_3795),
.Y(n_3937)
);

AO31x2_ASAP7_75t_L g3938 ( 
.A1(n_3747),
.A2(n_135),
.A3(n_133),
.B(n_134),
.Y(n_3938)
);

AND2x2_ASAP7_75t_L g3939 ( 
.A(n_3684),
.B(n_234),
.Y(n_3939)
);

CKINVDCx20_ASAP7_75t_R g3940 ( 
.A(n_3685),
.Y(n_3940)
);

AOI21xp5_ASAP7_75t_L g3941 ( 
.A1(n_3739),
.A2(n_135),
.B(n_235),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3739),
.A2(n_135),
.B(n_236),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3622),
.B(n_236),
.Y(n_3943)
);

INVxp67_ASAP7_75t_L g3944 ( 
.A(n_3802),
.Y(n_3944)
);

INVx3_ASAP7_75t_SL g3945 ( 
.A(n_3643),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3675),
.B(n_237),
.Y(n_3946)
);

AOI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3738),
.A2(n_237),
.B(n_238),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3781),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.Y(n_3948)
);

CKINVDCx5p33_ASAP7_75t_R g3949 ( 
.A(n_3695),
.Y(n_3949)
);

INVx2_ASAP7_75t_SL g3950 ( 
.A(n_3800),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3676),
.B(n_239),
.Y(n_3951)
);

NOR2xp67_ASAP7_75t_L g3952 ( 
.A(n_3817),
.B(n_241),
.Y(n_3952)
);

AOI22xp5_ASAP7_75t_L g3953 ( 
.A1(n_3781),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_3953)
);

AOI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3738),
.A2(n_3660),
.B(n_3657),
.Y(n_3954)
);

AO31x2_ASAP7_75t_L g3955 ( 
.A1(n_3667),
.A2(n_246),
.A3(n_244),
.B(n_245),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3660),
.A2(n_3692),
.B(n_3762),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_3770),
.B(n_247),
.Y(n_3957)
);

A2O1A1Ixp33_ASAP7_75t_L g3958 ( 
.A1(n_3772),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_3958)
);

AO31x2_ASAP7_75t_L g3959 ( 
.A1(n_3697),
.A2(n_254),
.A3(n_252),
.B(n_253),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3724),
.Y(n_3960)
);

OAI21x1_ASAP7_75t_L g3961 ( 
.A1(n_3706),
.A2(n_252),
.B(n_255),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3762),
.A2(n_255),
.B(n_257),
.Y(n_3962)
);

NOR2xp33_ASAP7_75t_L g3963 ( 
.A(n_3720),
.B(n_259),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3609),
.Y(n_3964)
);

AOI22xp5_ASAP7_75t_L g3965 ( 
.A1(n_3781),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_3965)
);

OAI21x1_ASAP7_75t_SL g3966 ( 
.A1(n_3733),
.A2(n_260),
.B(n_261),
.Y(n_3966)
);

OAI21x1_ASAP7_75t_L g3967 ( 
.A1(n_3611),
.A2(n_262),
.B(n_263),
.Y(n_3967)
);

INVx1_ASAP7_75t_SL g3968 ( 
.A(n_3801),
.Y(n_3968)
);

A2O1A1Ixp33_ASAP7_75t_L g3969 ( 
.A1(n_3831),
.A2(n_3627),
.B(n_3656),
.C(n_3824),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3620),
.B(n_264),
.Y(n_3970)
);

INVxp67_ASAP7_75t_SL g3971 ( 
.A(n_3673),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3630),
.Y(n_3972)
);

BUFx6f_ASAP7_75t_L g3973 ( 
.A(n_3800),
.Y(n_3973)
);

OAI21x1_ASAP7_75t_L g3974 ( 
.A1(n_3730),
.A2(n_265),
.B(n_266),
.Y(n_3974)
);

AO31x2_ASAP7_75t_L g3975 ( 
.A1(n_3713),
.A2(n_3748),
.A3(n_3639),
.B(n_3671),
.Y(n_3975)
);

OAI21x1_ASAP7_75t_L g3976 ( 
.A1(n_3757),
.A2(n_265),
.B(n_267),
.Y(n_3976)
);

OAI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3714),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_3977)
);

BUFx3_ASAP7_75t_L g3978 ( 
.A(n_3725),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3806),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3792),
.B(n_268),
.Y(n_3980)
);

AO31x2_ASAP7_75t_L g3981 ( 
.A1(n_3639),
.A2(n_272),
.A3(n_270),
.B(n_271),
.Y(n_3981)
);

OAI22x1_ASAP7_75t_L g3982 ( 
.A1(n_3734),
.A2(n_273),
.B1(n_270),
.B2(n_271),
.Y(n_3982)
);

OAI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3651),
.A2(n_274),
.B(n_276),
.Y(n_3983)
);

BUFx4_ASAP7_75t_SL g3984 ( 
.A(n_3808),
.Y(n_3984)
);

HB1xp67_ASAP7_75t_L g3985 ( 
.A(n_3677),
.Y(n_3985)
);

NOR2xp67_ASAP7_75t_SL g3986 ( 
.A(n_3800),
.B(n_274),
.Y(n_3986)
);

O2A1O1Ixp33_ASAP7_75t_SL g3987 ( 
.A1(n_3632),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3654),
.A2(n_277),
.B(n_278),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3630),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3677),
.Y(n_3990)
);

OAI22xp5_ASAP7_75t_L g3991 ( 
.A1(n_3785),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3806),
.Y(n_3992)
);

AO31x2_ASAP7_75t_L g3993 ( 
.A1(n_3736),
.A2(n_284),
.A3(n_282),
.B(n_283),
.Y(n_3993)
);

AO31x2_ASAP7_75t_L g3994 ( 
.A1(n_3729),
.A2(n_3707),
.A3(n_3763),
.B(n_3761),
.Y(n_3994)
);

OAI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3832),
.A2(n_3656),
.B(n_3606),
.Y(n_3995)
);

CKINVDCx8_ASAP7_75t_R g3996 ( 
.A(n_3811),
.Y(n_3996)
);

OAI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3619),
.A2(n_285),
.B(n_286),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3707),
.B(n_3804),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3801),
.B(n_3827),
.Y(n_3999)
);

BUFx2_ASAP7_75t_L g4000 ( 
.A(n_3605),
.Y(n_4000)
);

OAI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_3619),
.A2(n_285),
.B(n_286),
.Y(n_4001)
);

HB1xp67_ASAP7_75t_L g4002 ( 
.A(n_3677),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3796),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3796),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3750),
.A2(n_287),
.B(n_288),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3750),
.A2(n_3627),
.B(n_3715),
.Y(n_4006)
);

AOI21x1_ASAP7_75t_L g4007 ( 
.A1(n_3767),
.A2(n_290),
.B(n_291),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_SL g4008 ( 
.A(n_3642),
.B(n_292),
.Y(n_4008)
);

OAI21x1_ASAP7_75t_L g4009 ( 
.A1(n_3624),
.A2(n_3628),
.B(n_3633),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3711),
.B(n_293),
.Y(n_4010)
);

AO21x2_ASAP7_75t_L g4011 ( 
.A1(n_3629),
.A2(n_293),
.B(n_294),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3616),
.Y(n_4012)
);

OAI22x1_ASAP7_75t_L g4013 ( 
.A1(n_3710),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3708),
.B(n_295),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3653),
.A2(n_297),
.B(n_298),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3871),
.A2(n_3701),
.B(n_3775),
.Y(n_4016)
);

BUFx6f_ASAP7_75t_SL g4017 ( 
.A(n_3916),
.Y(n_4017)
);

OAI21x1_ASAP7_75t_L g4018 ( 
.A1(n_4009),
.A2(n_3818),
.B(n_3805),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3851),
.Y(n_4019)
);

BUFx6f_ASAP7_75t_L g4020 ( 
.A(n_3973),
.Y(n_4020)
);

AND2x4_ASAP7_75t_L g4021 ( 
.A(n_3960),
.B(n_3650),
.Y(n_4021)
);

OAI21x1_ASAP7_75t_L g4022 ( 
.A1(n_3850),
.A2(n_3682),
.B(n_3678),
.Y(n_4022)
);

HB1xp67_ASAP7_75t_L g4023 ( 
.A(n_3873),
.Y(n_4023)
);

INVxp67_ASAP7_75t_L g4024 ( 
.A(n_3851),
.Y(n_4024)
);

OAI21x1_ASAP7_75t_L g4025 ( 
.A1(n_3932),
.A2(n_3764),
.B(n_3649),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3954),
.A2(n_3709),
.B(n_3668),
.Y(n_4026)
);

AO31x2_ASAP7_75t_L g4027 ( 
.A1(n_3895),
.A2(n_3642),
.A3(n_3672),
.B(n_3768),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3883),
.B(n_3647),
.Y(n_4028)
);

HB1xp67_ASAP7_75t_L g4029 ( 
.A(n_3905),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3842),
.A2(n_3781),
.B1(n_3822),
.B2(n_3766),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_4003),
.B(n_3658),
.Y(n_4031)
);

AND2x4_ASAP7_75t_L g4032 ( 
.A(n_3929),
.B(n_3681),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3844),
.Y(n_4033)
);

OAI21x1_ASAP7_75t_L g4034 ( 
.A1(n_3855),
.A2(n_3661),
.B(n_3790),
.Y(n_4034)
);

INVx4_ASAP7_75t_L g4035 ( 
.A(n_3919),
.Y(n_4035)
);

NAND3x1_ASAP7_75t_L g4036 ( 
.A(n_3852),
.B(n_3746),
.C(n_3821),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3878),
.A2(n_3783),
.B(n_3779),
.Y(n_4037)
);

AO21x2_ASAP7_75t_L g4038 ( 
.A1(n_4004),
.A2(n_3751),
.B(n_3786),
.Y(n_4038)
);

INVx6_ASAP7_75t_L g4039 ( 
.A(n_3924),
.Y(n_4039)
);

CKINVDCx20_ASAP7_75t_R g4040 ( 
.A(n_3940),
.Y(n_4040)
);

OR2x2_ASAP7_75t_L g4041 ( 
.A(n_3998),
.B(n_3658),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3849),
.Y(n_4042)
);

OA21x2_ASAP7_75t_L g4043 ( 
.A1(n_3979),
.A2(n_3794),
.B(n_3798),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3918),
.A2(n_3803),
.B(n_3721),
.Y(n_4044)
);

OAI21x1_ASAP7_75t_L g4045 ( 
.A1(n_3995),
.A2(n_3683),
.B(n_3686),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3990),
.A2(n_3686),
.B(n_3753),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_SL g4047 ( 
.A1(n_3838),
.A2(n_3793),
.B1(n_3826),
.B2(n_3823),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3892),
.A2(n_3756),
.B(n_3812),
.Y(n_4048)
);

OAI21x1_ASAP7_75t_L g4049 ( 
.A1(n_3881),
.A2(n_3700),
.B(n_3727),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3870),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3840),
.Y(n_4051)
);

OA21x2_ASAP7_75t_L g4052 ( 
.A1(n_3992),
.A2(n_3726),
.B(n_3723),
.Y(n_4052)
);

CKINVDCx16_ASAP7_75t_R g4053 ( 
.A(n_3857),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3872),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3853),
.A2(n_3741),
.B(n_3732),
.Y(n_4055)
);

AND2x4_ASAP7_75t_L g4056 ( 
.A(n_3972),
.B(n_3719),
.Y(n_4056)
);

INVxp67_ASAP7_75t_SL g4057 ( 
.A(n_3886),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3846),
.B(n_3658),
.Y(n_4058)
);

NOR2x1_ASAP7_75t_SL g4059 ( 
.A(n_3973),
.B(n_3811),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3876),
.Y(n_4060)
);

NAND2x1p5_ASAP7_75t_L g4061 ( 
.A(n_3843),
.B(n_3811),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3887),
.Y(n_4062)
);

NOR2x1_ASAP7_75t_L g4063 ( 
.A(n_3964),
.B(n_3672),
.Y(n_4063)
);

BUFx6f_ASAP7_75t_SL g4064 ( 
.A(n_3909),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_SL g4065 ( 
.A(n_3996),
.B(n_3699),
.Y(n_4065)
);

AOI21xp5_ASAP7_75t_L g4066 ( 
.A1(n_3988),
.A2(n_3774),
.B(n_3742),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3989),
.B(n_3616),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3888),
.Y(n_4068)
);

BUFx2_ASAP7_75t_L g4069 ( 
.A(n_4000),
.Y(n_4069)
);

OAI21x1_ASAP7_75t_L g4070 ( 
.A1(n_3910),
.A2(n_3777),
.B(n_3702),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3911),
.Y(n_4071)
);

AOI221xp5_ASAP7_75t_L g4072 ( 
.A1(n_3913),
.A2(n_3788),
.B1(n_3810),
.B2(n_3717),
.C(n_3665),
.Y(n_4072)
);

AND2x4_ASAP7_75t_L g4073 ( 
.A(n_3927),
.B(n_3702),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3908),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3897),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3891),
.B(n_3647),
.Y(n_4076)
);

CKINVDCx16_ASAP7_75t_R g4077 ( 
.A(n_3978),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3896),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3968),
.Y(n_4079)
);

AO21x2_ASAP7_75t_L g4080 ( 
.A1(n_3971),
.A2(n_3717),
.B(n_3699),
.Y(n_4080)
);

AOI21xp33_ASAP7_75t_L g4081 ( 
.A1(n_3889),
.A2(n_3777),
.B(n_297),
.Y(n_4081)
);

OA21x2_ASAP7_75t_L g4082 ( 
.A1(n_3941),
.A2(n_3647),
.B(n_3765),
.Y(n_4082)
);

NAND3xp33_ASAP7_75t_L g4083 ( 
.A(n_3898),
.B(n_298),
.C(n_299),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3999),
.B(n_299),
.Y(n_4084)
);

NOR2xp67_ASAP7_75t_L g4085 ( 
.A(n_3985),
.B(n_4002),
.Y(n_4085)
);

O2A1O1Ixp33_ASAP7_75t_SL g4086 ( 
.A1(n_3858),
.A2(n_3835),
.B(n_3882),
.C(n_3900),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3848),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_3904),
.B(n_300),
.Y(n_4088)
);

AND2x6_ASAP7_75t_L g4089 ( 
.A(n_3953),
.B(n_300),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3926),
.A2(n_304),
.B1(n_301),
.B2(n_302),
.Y(n_4090)
);

INVx1_ASAP7_75t_SL g4091 ( 
.A(n_3868),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_4012),
.B(n_302),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3930),
.Y(n_4093)
);

AND2x4_ASAP7_75t_L g4094 ( 
.A(n_3928),
.B(n_304),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3848),
.Y(n_4095)
);

OAI211xp5_ASAP7_75t_L g4096 ( 
.A1(n_3965),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3854),
.B(n_305),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3875),
.A2(n_688),
.B1(n_308),
.B2(n_306),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3950),
.B(n_307),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3934),
.Y(n_4100)
);

INVx4_ASAP7_75t_L g4101 ( 
.A(n_3949),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_L g4102 ( 
.A1(n_3861),
.A2(n_3856),
.B1(n_3837),
.B2(n_3834),
.Y(n_4102)
);

OAI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_3947),
.A2(n_4005),
.B(n_3894),
.Y(n_4103)
);

CKINVDCx8_ASAP7_75t_R g4104 ( 
.A(n_3877),
.Y(n_4104)
);

AND2x2_ASAP7_75t_SL g4105 ( 
.A(n_4008),
.B(n_308),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_SL g4106 ( 
.A1(n_3969),
.A2(n_309),
.B(n_310),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3845),
.A2(n_309),
.B(n_311),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3859),
.A2(n_313),
.B(n_315),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3934),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3914),
.A2(n_313),
.B(n_315),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3934),
.Y(n_4111)
);

CKINVDCx20_ASAP7_75t_R g4112 ( 
.A(n_3945),
.Y(n_4112)
);

OAI21x1_ASAP7_75t_L g4113 ( 
.A1(n_3956),
.A2(n_317),
.B(n_319),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3975),
.B(n_317),
.Y(n_4114)
);

AOI21xp33_ASAP7_75t_SL g4115 ( 
.A1(n_3982),
.A2(n_3836),
.B(n_3874),
.Y(n_4115)
);

O2A1O1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_3925),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_4116)
);

OAI21x1_ASAP7_75t_L g4117 ( 
.A1(n_3935),
.A2(n_322),
.B(n_323),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3944),
.B(n_3903),
.Y(n_4118)
);

NAND2x1_ASAP7_75t_L g4119 ( 
.A(n_3973),
.B(n_3860),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3975),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3867),
.A2(n_325),
.B1(n_322),
.B2(n_324),
.Y(n_4121)
);

OR2x6_ASAP7_75t_L g4122 ( 
.A(n_4006),
.B(n_324),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3962),
.A2(n_686),
.B(n_325),
.Y(n_4123)
);

OAI21x1_ASAP7_75t_L g4124 ( 
.A1(n_3974),
.A2(n_326),
.B(n_327),
.Y(n_4124)
);

BUFx3_ASAP7_75t_L g4125 ( 
.A(n_3890),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3885),
.A2(n_331),
.B1(n_326),
.B2(n_328),
.Y(n_4126)
);

OAI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_3948),
.A2(n_332),
.B1(n_328),
.B2(n_331),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3923),
.B(n_686),
.Y(n_4128)
);

NOR2x1_ASAP7_75t_SL g4129 ( 
.A(n_4011),
.B(n_333),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_3909),
.B(n_333),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_3937),
.B(n_334),
.Y(n_4131)
);

AOI22xp33_ASAP7_75t_L g4132 ( 
.A1(n_3884),
.A2(n_338),
.B1(n_335),
.B2(n_336),
.Y(n_4132)
);

INVx3_ASAP7_75t_SL g4133 ( 
.A(n_3915),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3848),
.Y(n_4134)
);

CKINVDCx14_ASAP7_75t_R g4135 ( 
.A(n_3937),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3880),
.Y(n_4136)
);

OAI21x1_ASAP7_75t_L g4137 ( 
.A1(n_3961),
.A2(n_336),
.B(n_338),
.Y(n_4137)
);

HB1xp67_ASAP7_75t_L g4138 ( 
.A(n_3880),
.Y(n_4138)
);

OA21x2_ASAP7_75t_L g4139 ( 
.A1(n_3942),
.A2(n_3967),
.B(n_3865),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3864),
.A2(n_339),
.B(n_340),
.Y(n_4140)
);

CKINVDCx11_ASAP7_75t_R g4141 ( 
.A(n_3901),
.Y(n_4141)
);

HB1xp67_ASAP7_75t_L g4142 ( 
.A(n_3880),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_SL g4143 ( 
.A1(n_3839),
.A2(n_3866),
.B(n_3966),
.Y(n_4143)
);

BUFx4f_ASAP7_75t_L g4144 ( 
.A(n_3915),
.Y(n_4144)
);

AOI21xp5_ASAP7_75t_L g4145 ( 
.A1(n_3847),
.A2(n_4001),
.B(n_3997),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3959),
.Y(n_4146)
);

AND2x4_ASAP7_75t_L g4147 ( 
.A(n_3994),
.B(n_339),
.Y(n_4147)
);

O2A1O1Ixp33_ASAP7_75t_L g4148 ( 
.A1(n_3958),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_4148)
);

INVx3_ASAP7_75t_L g4149 ( 
.A(n_3901),
.Y(n_4149)
);

HB1xp67_ASAP7_75t_L g4150 ( 
.A(n_3994),
.Y(n_4150)
);

OAI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3912),
.A2(n_341),
.B(n_342),
.Y(n_4151)
);

OA21x2_ASAP7_75t_L g4152 ( 
.A1(n_3983),
.A2(n_344),
.B(n_345),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3922),
.B(n_685),
.Y(n_4153)
);

AND2x4_ASAP7_75t_L g4154 ( 
.A(n_3994),
.B(n_344),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3959),
.Y(n_4155)
);

OAI21x1_ASAP7_75t_L g4156 ( 
.A1(n_3933),
.A2(n_346),
.B(n_347),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_SL g4157 ( 
.A1(n_3991),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3959),
.Y(n_4158)
);

OAI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_3977),
.A2(n_349),
.B(n_350),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_3984),
.Y(n_4160)
);

AO31x2_ASAP7_75t_L g4161 ( 
.A1(n_4013),
.A2(n_353),
.A3(n_351),
.B(n_352),
.Y(n_4161)
);

OR2x2_ASAP7_75t_L g4162 ( 
.A(n_3931),
.B(n_351),
.Y(n_4162)
);

BUFx2_ASAP7_75t_L g4163 ( 
.A(n_3901),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3975),
.Y(n_4164)
);

BUFx2_ASAP7_75t_L g4165 ( 
.A(n_3907),
.Y(n_4165)
);

OR2x6_ASAP7_75t_L g4166 ( 
.A(n_3976),
.B(n_352),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_3907),
.Y(n_4167)
);

INVx3_ASAP7_75t_L g4168 ( 
.A(n_3907),
.Y(n_4168)
);

AO21x2_ASAP7_75t_L g4169 ( 
.A1(n_3952),
.A2(n_3902),
.B(n_3841),
.Y(n_4169)
);

CKINVDCx20_ASAP7_75t_R g4170 ( 
.A(n_4040),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_4030),
.A2(n_3917),
.B1(n_3957),
.B2(n_3963),
.Y(n_4171)
);

OAI21x1_ASAP7_75t_SL g4172 ( 
.A1(n_4059),
.A2(n_4007),
.B(n_3906),
.Y(n_4172)
);

OAI21x1_ASAP7_75t_L g4173 ( 
.A1(n_4063),
.A2(n_4015),
.B(n_3879),
.Y(n_4173)
);

AOI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_4098),
.A2(n_4010),
.B1(n_3986),
.B2(n_3920),
.Y(n_4174)
);

BUFx8_ASAP7_75t_SL g4175 ( 
.A(n_4017),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4069),
.Y(n_4176)
);

OAI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_4103),
.A2(n_4014),
.B(n_3980),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4029),
.Y(n_4178)
);

NOR2xp33_ASAP7_75t_L g4179 ( 
.A(n_4035),
.B(n_3936),
.Y(n_4179)
);

OA21x2_ASAP7_75t_L g4180 ( 
.A1(n_4057),
.A2(n_3951),
.B(n_3946),
.Y(n_4180)
);

AO21x2_ASAP7_75t_L g4181 ( 
.A1(n_4114),
.A2(n_3943),
.B(n_3869),
.Y(n_4181)
);

AO21x2_ASAP7_75t_L g4182 ( 
.A1(n_4114),
.A2(n_3987),
.B(n_3862),
.Y(n_4182)
);

AO21x2_ASAP7_75t_L g4183 ( 
.A1(n_4085),
.A2(n_3862),
.B(n_3939),
.Y(n_4183)
);

OAI21x1_ASAP7_75t_L g4184 ( 
.A1(n_4063),
.A2(n_3970),
.B(n_3863),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4021),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_SL g4186 ( 
.A(n_4053),
.B(n_3862),
.Y(n_4186)
);

BUFx3_ASAP7_75t_L g4187 ( 
.A(n_4112),
.Y(n_4187)
);

BUFx8_ASAP7_75t_L g4188 ( 
.A(n_4017),
.Y(n_4188)
);

AOI21xp33_ASAP7_75t_SL g4189 ( 
.A1(n_4105),
.A2(n_353),
.B(n_354),
.Y(n_4189)
);

AND2x6_ASAP7_75t_L g4190 ( 
.A(n_4098),
.B(n_3893),
.Y(n_4190)
);

AO21x2_ASAP7_75t_L g4191 ( 
.A1(n_4085),
.A2(n_4164),
.B(n_4120),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4075),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_4019),
.B(n_4024),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_4103),
.A2(n_3893),
.B(n_3899),
.Y(n_4194)
);

AO31x2_ASAP7_75t_L g4195 ( 
.A1(n_4136),
.A2(n_3863),
.A3(n_3899),
.B(n_3981),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_4106),
.A2(n_3893),
.B(n_3899),
.Y(n_4196)
);

OAI21x1_ASAP7_75t_L g4197 ( 
.A1(n_4022),
.A2(n_3863),
.B(n_3955),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4033),
.Y(n_4198)
);

OAI21x1_ASAP7_75t_L g4199 ( 
.A1(n_4031),
.A2(n_3955),
.B(n_3981),
.Y(n_4199)
);

AOI21x1_ASAP7_75t_L g4200 ( 
.A1(n_4119),
.A2(n_3955),
.B(n_3981),
.Y(n_4200)
);

OAI21x1_ASAP7_75t_L g4201 ( 
.A1(n_4031),
.A2(n_3938),
.B(n_3921),
.Y(n_4201)
);

A2O1A1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4115),
.A2(n_3938),
.B(n_3921),
.C(n_3993),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4050),
.Y(n_4203)
);

OAI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_4104),
.A2(n_3938),
.B1(n_3921),
.B2(n_3993),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4054),
.Y(n_4205)
);

OA21x2_ASAP7_75t_L g4206 ( 
.A1(n_4078),
.A2(n_3993),
.B(n_355),
.Y(n_4206)
);

OAI21x1_ASAP7_75t_SL g4207 ( 
.A1(n_4129),
.A2(n_355),
.B(n_356),
.Y(n_4207)
);

OR2x2_ASAP7_75t_L g4208 ( 
.A(n_4041),
.B(n_683),
.Y(n_4208)
);

OAI21x1_ASAP7_75t_L g4209 ( 
.A1(n_4058),
.A2(n_356),
.B(n_357),
.Y(n_4209)
);

CKINVDCx20_ASAP7_75t_R g4210 ( 
.A(n_4077),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4060),
.Y(n_4211)
);

OAI21x1_ASAP7_75t_L g4212 ( 
.A1(n_4058),
.A2(n_357),
.B(n_358),
.Y(n_4212)
);

AO21x2_ASAP7_75t_L g4213 ( 
.A1(n_4138),
.A2(n_4142),
.B(n_4095),
.Y(n_4213)
);

BUFx6f_ASAP7_75t_L g4214 ( 
.A(n_4035),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4062),
.Y(n_4215)
);

AOI21x1_ASAP7_75t_L g4216 ( 
.A1(n_4037),
.A2(n_358),
.B(n_359),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4038),
.B(n_359),
.Y(n_4217)
);

OR2x2_ASAP7_75t_L g4218 ( 
.A(n_4023),
.B(n_4076),
.Y(n_4218)
);

AOI21xp5_ASAP7_75t_SL g4219 ( 
.A1(n_4147),
.A2(n_360),
.B(n_361),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4042),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4093),
.B(n_4073),
.Y(n_4221)
);

AO21x2_ASAP7_75t_L g4222 ( 
.A1(n_4087),
.A2(n_360),
.B(n_362),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_4073),
.B(n_362),
.Y(n_4223)
);

AND2x4_ASAP7_75t_L g4224 ( 
.A(n_4147),
.B(n_363),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4068),
.Y(n_4225)
);

A2O1A1Ixp33_ASAP7_75t_L g4226 ( 
.A1(n_4115),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_4226)
);

OAI22xp5_ASAP7_75t_L g4227 ( 
.A1(n_4102),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_4227)
);

NOR2x1_ASAP7_75t_L g4228 ( 
.A(n_4038),
.B(n_366),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4071),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4021),
.Y(n_4230)
);

CKINVDCx14_ASAP7_75t_R g4231 ( 
.A(n_4135),
.Y(n_4231)
);

A2O1A1Ixp33_ASAP7_75t_L g4232 ( 
.A1(n_4148),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_4232)
);

BUFx8_ASAP7_75t_L g4233 ( 
.A(n_4064),
.Y(n_4233)
);

INVx3_ASAP7_75t_L g4234 ( 
.A(n_4020),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4080),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4074),
.Y(n_4236)
);

OA21x2_ASAP7_75t_L g4237 ( 
.A1(n_4134),
.A2(n_367),
.B(n_368),
.Y(n_4237)
);

OAI21x1_ASAP7_75t_SL g4238 ( 
.A1(n_4143),
.A2(n_370),
.B(n_371),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_4145),
.A2(n_373),
.B(n_374),
.Y(n_4239)
);

NOR2x1_ASAP7_75t_SL g4240 ( 
.A(n_4080),
.B(n_373),
.Y(n_4240)
);

OA21x2_ASAP7_75t_L g4241 ( 
.A1(n_4146),
.A2(n_4158),
.B(n_4155),
.Y(n_4241)
);

OAI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_4083),
.A2(n_375),
.B(n_376),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4052),
.B(n_375),
.Y(n_4243)
);

OR2x2_ASAP7_75t_L g4244 ( 
.A(n_4091),
.B(n_682),
.Y(n_4244)
);

BUFx2_ASAP7_75t_L g4245 ( 
.A(n_4020),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4091),
.B(n_4079),
.Y(n_4246)
);

INVx2_ASAP7_75t_L g4247 ( 
.A(n_4051),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4067),
.B(n_376),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_SL g4249 ( 
.A1(n_4089),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_4249)
);

OA21x2_ASAP7_75t_L g4250 ( 
.A1(n_4070),
.A2(n_377),
.B(n_379),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4052),
.B(n_4028),
.Y(n_4251)
);

OAI22xp5_ASAP7_75t_L g4252 ( 
.A1(n_4083),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4043),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_4039),
.B(n_4064),
.Y(n_4254)
);

CKINVDCx8_ASAP7_75t_R g4255 ( 
.A(n_4160),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4043),
.Y(n_4256)
);

INVx3_ASAP7_75t_L g4257 ( 
.A(n_4020),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4118),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4163),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4165),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4150),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4154),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_4123),
.A2(n_380),
.B(n_381),
.Y(n_4263)
);

CKINVDCx20_ASAP7_75t_R g4264 ( 
.A(n_4141),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4154),
.B(n_382),
.Y(n_4265)
);

BUFx12f_ASAP7_75t_L g4266 ( 
.A(n_4101),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4067),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4149),
.Y(n_4268)
);

CKINVDCx5p33_ASAP7_75t_R g4269 ( 
.A(n_4167),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4100),
.B(n_384),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4082),
.B(n_385),
.Y(n_4271)
);

OAI21x1_ASAP7_75t_L g4272 ( 
.A1(n_4045),
.A2(n_386),
.B(n_387),
.Y(n_4272)
);

OR2x6_ASAP7_75t_L g4273 ( 
.A(n_4061),
.B(n_387),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4149),
.Y(n_4274)
);

BUFx6f_ASAP7_75t_L g4275 ( 
.A(n_4094),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4168),
.Y(n_4276)
);

OAI21x1_ASAP7_75t_L g4277 ( 
.A1(n_4046),
.A2(n_388),
.B(n_389),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4168),
.Y(n_4278)
);

OAI21x1_ASAP7_75t_L g4279 ( 
.A1(n_4026),
.A2(n_390),
.B(n_391),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4032),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4082),
.B(n_392),
.Y(n_4281)
);

AOI22xp33_ASAP7_75t_L g4282 ( 
.A1(n_4089),
.A2(n_681),
.B1(n_394),
.B2(n_392),
.Y(n_4282)
);

NAND2x1_ASAP7_75t_L g4283 ( 
.A(n_4039),
.B(n_393),
.Y(n_4283)
);

AO31x2_ASAP7_75t_L g4284 ( 
.A1(n_4109),
.A2(n_397),
.A3(n_395),
.B(n_396),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_4139),
.B(n_395),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4111),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4032),
.Y(n_4287)
);

OA21x2_ASAP7_75t_L g4288 ( 
.A1(n_4034),
.A2(n_396),
.B(n_397),
.Y(n_4288)
);

OAI21x1_ASAP7_75t_L g4289 ( 
.A1(n_4025),
.A2(n_398),
.B(n_399),
.Y(n_4289)
);

INVx2_ASAP7_75t_SL g4290 ( 
.A(n_4125),
.Y(n_4290)
);

NOR2xp33_ASAP7_75t_L g4291 ( 
.A(n_4101),
.B(n_398),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4056),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4056),
.Y(n_4293)
);

OAI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_4036),
.A2(n_400),
.B(n_401),
.Y(n_4294)
);

AO21x2_ASAP7_75t_L g4295 ( 
.A1(n_4081),
.A2(n_400),
.B(n_401),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_4055),
.B(n_402),
.Y(n_4296)
);

AO31x2_ASAP7_75t_L g4297 ( 
.A1(n_4016),
.A2(n_405),
.A3(n_403),
.B(n_404),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4169),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4018),
.A2(n_403),
.B(n_404),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4169),
.Y(n_4300)
);

HB1xp67_ASAP7_75t_L g4301 ( 
.A(n_4139),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4094),
.Y(n_4302)
);

INVx3_ASAP7_75t_L g4303 ( 
.A(n_4144),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4133),
.B(n_405),
.Y(n_4304)
);

BUFx4f_ASAP7_75t_L g4305 ( 
.A(n_4122),
.Y(n_4305)
);

OAI21x1_ASAP7_75t_L g4306 ( 
.A1(n_4049),
.A2(n_406),
.B(n_407),
.Y(n_4306)
);

HB1xp67_ASAP7_75t_L g4307 ( 
.A(n_4152),
.Y(n_4307)
);

OAI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_4122),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4081),
.A2(n_408),
.B(n_409),
.Y(n_4309)
);

OAI21x1_ASAP7_75t_L g4310 ( 
.A1(n_4048),
.A2(n_410),
.B(n_411),
.Y(n_4310)
);

OA21x2_ASAP7_75t_L g4311 ( 
.A1(n_4044),
.A2(n_411),
.B(n_412),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4152),
.Y(n_4312)
);

O2A1O1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_4086),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_4313)
);

AND2x4_ASAP7_75t_SL g4314 ( 
.A(n_4092),
.B(n_413),
.Y(n_4314)
);

NAND3xp33_ASAP7_75t_L g4315 ( 
.A(n_4151),
.B(n_414),
.C(n_415),
.Y(n_4315)
);

BUFx12f_ASAP7_75t_L g4316 ( 
.A(n_4131),
.Y(n_4316)
);

BUFx2_ASAP7_75t_SL g4317 ( 
.A(n_4099),
.Y(n_4317)
);

AOI211xp5_ASAP7_75t_L g4318 ( 
.A1(n_4151),
.A2(n_419),
.B(n_416),
.C(n_418),
.Y(n_4318)
);

BUFx8_ASAP7_75t_L g4319 ( 
.A(n_4097),
.Y(n_4319)
);

OAI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4122),
.A2(n_4140),
.B(n_4044),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_4116),
.A2(n_419),
.B(n_420),
.Y(n_4321)
);

INVx5_ASAP7_75t_L g4322 ( 
.A(n_4175),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4234),
.Y(n_4323)
);

OAI22xp5_ASAP7_75t_L g4324 ( 
.A1(n_4305),
.A2(n_4090),
.B1(n_4047),
.B2(n_4121),
.Y(n_4324)
);

BUFx2_ASAP7_75t_L g4325 ( 
.A(n_4233),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_SL g4326 ( 
.A1(n_4305),
.A2(n_4089),
.B1(n_4096),
.B2(n_4159),
.Y(n_4326)
);

OAI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4318),
.A2(n_4132),
.B1(n_4126),
.B2(n_4072),
.Y(n_4327)
);

BUFx3_ASAP7_75t_L g4328 ( 
.A(n_4188),
.Y(n_4328)
);

CKINVDCx5p33_ASAP7_75t_R g4329 ( 
.A(n_4170),
.Y(n_4329)
);

AOI22xp33_ASAP7_75t_L g4330 ( 
.A1(n_4190),
.A2(n_4089),
.B1(n_4159),
.B2(n_4157),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4229),
.Y(n_4331)
);

AOI22xp33_ASAP7_75t_L g4332 ( 
.A1(n_4190),
.A2(n_4140),
.B1(n_4127),
.B2(n_4107),
.Y(n_4332)
);

OAI211xp5_ASAP7_75t_L g4333 ( 
.A1(n_4313),
.A2(n_4130),
.B(n_4110),
.C(n_4088),
.Y(n_4333)
);

OAI222xp33_ASAP7_75t_L g4334 ( 
.A1(n_4186),
.A2(n_4166),
.B1(n_4127),
.B2(n_4162),
.C1(n_4066),
.C2(n_4084),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_L g4335 ( 
.A1(n_4190),
.A2(n_4166),
.B1(n_4144),
.B2(n_4113),
.Y(n_4335)
);

BUFx4f_ASAP7_75t_SL g4336 ( 
.A(n_4188),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4190),
.A2(n_4166),
.B1(n_4065),
.B2(n_4153),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4236),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4234),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_4214),
.B(n_4128),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4257),
.Y(n_4341)
);

BUFx12f_ASAP7_75t_L g4342 ( 
.A(n_4233),
.Y(n_4342)
);

AOI22xp33_ASAP7_75t_L g4343 ( 
.A1(n_4320),
.A2(n_4065),
.B1(n_4092),
.B2(n_4156),
.Y(n_4343)
);

AOI22xp33_ASAP7_75t_L g4344 ( 
.A1(n_4320),
.A2(n_4137),
.B1(n_4124),
.B2(n_4099),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4257),
.Y(n_4345)
);

OAI22xp5_ASAP7_75t_L g4346 ( 
.A1(n_4315),
.A2(n_4027),
.B1(n_4161),
.B2(n_4108),
.Y(n_4346)
);

INVxp67_ASAP7_75t_L g4347 ( 
.A(n_4240),
.Y(n_4347)
);

INVx1_ASAP7_75t_SL g4348 ( 
.A(n_4210),
.Y(n_4348)
);

OAI21xp33_ASAP7_75t_L g4349 ( 
.A1(n_4226),
.A2(n_4117),
.B(n_4027),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4194),
.A2(n_4027),
.B1(n_4161),
.B2(n_422),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_4315),
.A2(n_4161),
.B1(n_422),
.B2(n_420),
.Y(n_4351)
);

OAI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_4294),
.A2(n_421),
.B(n_423),
.Y(n_4352)
);

AND2x2_ASAP7_75t_L g4353 ( 
.A(n_4221),
.B(n_421),
.Y(n_4353)
);

AOI22xp33_ASAP7_75t_L g4354 ( 
.A1(n_4242),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_4354)
);

AOI22xp33_ASAP7_75t_L g4355 ( 
.A1(n_4242),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_4355)
);

BUFx3_ASAP7_75t_L g4356 ( 
.A(n_4264),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4252),
.A2(n_4204),
.B1(n_4318),
.B2(n_4227),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_4214),
.B(n_427),
.Y(n_4358)
);

HB1xp67_ASAP7_75t_L g4359 ( 
.A(n_4250),
.Y(n_4359)
);

AOI22xp33_ASAP7_75t_L g4360 ( 
.A1(n_4239),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_4360)
);

HB1xp67_ASAP7_75t_L g4361 ( 
.A(n_4250),
.Y(n_4361)
);

INVx2_ASAP7_75t_SL g4362 ( 
.A(n_4214),
.Y(n_4362)
);

BUFx8_ASAP7_75t_SL g4363 ( 
.A(n_4266),
.Y(n_4363)
);

OAI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4196),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4245),
.Y(n_4365)
);

OAI22xp5_ASAP7_75t_L g4366 ( 
.A1(n_4249),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_4366)
);

AOI22xp33_ASAP7_75t_L g4367 ( 
.A1(n_4252),
.A2(n_435),
.B1(n_432),
.B2(n_434),
.Y(n_4367)
);

OAI22xp5_ASAP7_75t_L g4368 ( 
.A1(n_4249),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_4368)
);

INVx4_ASAP7_75t_L g4369 ( 
.A(n_4273),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4198),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4203),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4260),
.B(n_436),
.Y(n_4372)
);

OAI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_4294),
.A2(n_4174),
.B1(n_4228),
.B2(n_4282),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_4268),
.Y(n_4374)
);

BUFx2_ASAP7_75t_L g4375 ( 
.A(n_4231),
.Y(n_4375)
);

INVx5_ASAP7_75t_SL g4376 ( 
.A(n_4273),
.Y(n_4376)
);

BUFx4f_ASAP7_75t_SL g4377 ( 
.A(n_4187),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4274),
.Y(n_4378)
);

CKINVDCx20_ASAP7_75t_R g4379 ( 
.A(n_4255),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4181),
.B(n_438),
.Y(n_4380)
);

INVx3_ASAP7_75t_L g4381 ( 
.A(n_4275),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4181),
.B(n_438),
.Y(n_4382)
);

BUFx6f_ASAP7_75t_L g4383 ( 
.A(n_4273),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4311),
.A2(n_442),
.B1(n_439),
.B2(n_440),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_SL g4385 ( 
.A1(n_4171),
.A2(n_4183),
.B1(n_4311),
.B2(n_4177),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4180),
.B(n_439),
.Y(n_4386)
);

OAI222xp33_ASAP7_75t_L g4387 ( 
.A1(n_4228),
.A2(n_440),
.B1(n_443),
.B2(n_444),
.C1(n_445),
.C2(n_446),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_4321),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4174),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4276),
.Y(n_4390)
);

AOI22xp33_ASAP7_75t_L g4391 ( 
.A1(n_4295),
.A2(n_4309),
.B1(n_4227),
.B2(n_4171),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_4202),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_L g4393 ( 
.A(n_4254),
.B(n_451),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_4269),
.Y(n_4394)
);

AOI22xp33_ASAP7_75t_SL g4395 ( 
.A1(n_4183),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4285),
.A2(n_456),
.B1(n_453),
.B2(n_455),
.Y(n_4396)
);

HB1xp67_ASAP7_75t_L g4397 ( 
.A(n_4307),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4205),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4180),
.B(n_455),
.Y(n_4399)
);

AOI22xp33_ASAP7_75t_L g4400 ( 
.A1(n_4295),
.A2(n_4177),
.B1(n_4258),
.B2(n_4301),
.Y(n_4400)
);

AOI22xp33_ASAP7_75t_SL g4401 ( 
.A1(n_4317),
.A2(n_459),
.B1(n_456),
.B2(n_457),
.Y(n_4401)
);

AOI22xp33_ASAP7_75t_SL g4402 ( 
.A1(n_4308),
.A2(n_462),
.B1(n_459),
.B2(n_461),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4278),
.Y(n_4403)
);

OAI22xp5_ASAP7_75t_L g4404 ( 
.A1(n_4232),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_4404)
);

INVx4_ASAP7_75t_SL g4405 ( 
.A(n_4297),
.Y(n_4405)
);

AOI22xp33_ASAP7_75t_L g4406 ( 
.A1(n_4182),
.A2(n_466),
.B1(n_463),
.B2(n_465),
.Y(n_4406)
);

BUFx6f_ASAP7_75t_L g4407 ( 
.A(n_4299),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_4182),
.A2(n_468),
.B1(n_465),
.B2(n_467),
.Y(n_4408)
);

AOI22xp33_ASAP7_75t_L g4409 ( 
.A1(n_4263),
.A2(n_470),
.B1(n_467),
.B2(n_468),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4267),
.B(n_471),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4303),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4211),
.Y(n_4412)
);

HB1xp67_ASAP7_75t_L g4413 ( 
.A(n_4312),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4280),
.B(n_472),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4308),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_4415)
);

AOI22xp33_ASAP7_75t_L g4416 ( 
.A1(n_4303),
.A2(n_4296),
.B1(n_4285),
.B2(n_4179),
.Y(n_4416)
);

AOI22xp33_ASAP7_75t_L g4417 ( 
.A1(n_4296),
.A2(n_478),
.B1(n_475),
.B2(n_477),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4292),
.B(n_4262),
.Y(n_4418)
);

AOI222xp33_ASAP7_75t_L g4419 ( 
.A1(n_4271),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.C1(n_481),
.C2(n_482),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4193),
.B(n_479),
.Y(n_4420)
);

AOI22xp5_ASAP7_75t_L g4421 ( 
.A1(n_4271),
.A2(n_484),
.B1(n_481),
.B2(n_483),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4172),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4215),
.Y(n_4423)
);

OAI22xp5_ASAP7_75t_L g4424 ( 
.A1(n_4281),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4192),
.Y(n_4425)
);

OAI22xp5_ASAP7_75t_L g4426 ( 
.A1(n_4281),
.A2(n_489),
.B1(n_486),
.B2(n_488),
.Y(n_4426)
);

OAI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_4217),
.A2(n_4243),
.B1(n_4275),
.B2(n_4208),
.Y(n_4427)
);

AOI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4316),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4241),
.Y(n_4429)
);

OAI22xp33_ASAP7_75t_L g4430 ( 
.A1(n_4243),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4291),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4241),
.Y(n_4432)
);

AOI22xp33_ASAP7_75t_L g4433 ( 
.A1(n_4238),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_4433)
);

AOI22xp33_ASAP7_75t_L g4434 ( 
.A1(n_4288),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_4434)
);

OAI22xp33_ASAP7_75t_L g4435 ( 
.A1(n_4217),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_4435)
);

AOI22xp5_ASAP7_75t_L g4436 ( 
.A1(n_4224),
.A2(n_499),
.B1(n_501),
.B2(n_502),
.Y(n_4436)
);

OAI21xp5_ASAP7_75t_SL g4437 ( 
.A1(n_4189),
.A2(n_501),
.B(n_502),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4178),
.Y(n_4438)
);

INVx4_ASAP7_75t_L g4439 ( 
.A(n_4224),
.Y(n_4439)
);

AND2x2_ASAP7_75t_L g4440 ( 
.A(n_4176),
.B(n_503),
.Y(n_4440)
);

OAI22xp5_ASAP7_75t_L g4441 ( 
.A1(n_4189),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_4441)
);

AOI22xp33_ASAP7_75t_L g4442 ( 
.A1(n_4288),
.A2(n_504),
.B1(n_505),
.B2(n_507),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_4246),
.A2(n_4206),
.B1(n_4275),
.B2(n_4302),
.Y(n_4443)
);

NAND2xp33_ASAP7_75t_SL g4444 ( 
.A(n_4283),
.B(n_507),
.Y(n_4444)
);

BUFx6f_ASAP7_75t_L g4445 ( 
.A(n_4289),
.Y(n_4445)
);

AOI22xp33_ASAP7_75t_L g4446 ( 
.A1(n_4206),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_4446)
);

BUFx3_ASAP7_75t_L g4447 ( 
.A(n_4319),
.Y(n_4447)
);

OAI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_4251),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_4448)
);

AOI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4287),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_4449)
);

HB1xp67_ASAP7_75t_L g4450 ( 
.A(n_4298),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4220),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_SL g4452 ( 
.A1(n_4222),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_4452)
);

BUFx2_ASAP7_75t_L g4453 ( 
.A(n_4319),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4185),
.Y(n_4454)
);

INVx6_ASAP7_75t_L g4455 ( 
.A(n_4304),
.Y(n_4455)
);

INVx2_ASAP7_75t_SL g4456 ( 
.A(n_4290),
.Y(n_4456)
);

OAI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_4219),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4293),
.B(n_516),
.Y(n_4458)
);

AOI22xp33_ASAP7_75t_SL g4459 ( 
.A1(n_4222),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_4459)
);

OAI21xp33_ASAP7_75t_L g4460 ( 
.A1(n_4216),
.A2(n_519),
.B(n_520),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4244),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4225),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4237),
.Y(n_4463)
);

OAI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_4237),
.A2(n_522),
.B1(n_523),
.B2(n_525),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4261),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_L g4466 ( 
.A1(n_4259),
.A2(n_525),
.B1(n_526),
.B2(n_527),
.Y(n_4466)
);

OAI22xp5_ASAP7_75t_L g4467 ( 
.A1(n_4265),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4265),
.A2(n_4251),
.B1(n_4200),
.B2(n_4314),
.Y(n_4468)
);

OAI22xp33_ASAP7_75t_L g4469 ( 
.A1(n_4218),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_SL g4470 ( 
.A1(n_4207),
.A2(n_677),
.B1(n_531),
.B2(n_532),
.Y(n_4470)
);

INVx2_ASAP7_75t_L g4471 ( 
.A(n_4230),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4286),
.B(n_529),
.Y(n_4472)
);

BUFx6f_ASAP7_75t_L g4473 ( 
.A(n_4342),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4413),
.Y(n_4474)
);

INVx3_ASAP7_75t_L g4475 ( 
.A(n_4369),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4383),
.Y(n_4476)
);

OR2x2_ASAP7_75t_L g4477 ( 
.A(n_4463),
.B(n_4300),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4331),
.Y(n_4478)
);

INVx2_ASAP7_75t_SL g4479 ( 
.A(n_4322),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4381),
.B(n_4213),
.Y(n_4480)
);

AO21x2_ASAP7_75t_L g4481 ( 
.A1(n_4380),
.A2(n_4256),
.B(n_4253),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4338),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4381),
.B(n_4213),
.Y(n_4483)
);

AO21x2_ASAP7_75t_L g4484 ( 
.A1(n_4382),
.A2(n_4235),
.B(n_4197),
.Y(n_4484)
);

OAI21x1_ASAP7_75t_L g4485 ( 
.A1(n_4468),
.A2(n_4199),
.B(n_4201),
.Y(n_4485)
);

AO21x2_ASAP7_75t_L g4486 ( 
.A1(n_4386),
.A2(n_4272),
.B(n_4279),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4370),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4383),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4383),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4391),
.B(n_4223),
.Y(n_4490)
);

INVx2_ASAP7_75t_SL g4491 ( 
.A(n_4322),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4371),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4439),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4439),
.Y(n_4494)
);

OAI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_4385),
.A2(n_4184),
.B(n_4209),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4429),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_4432),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4407),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4398),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4407),
.Y(n_4500)
);

OAI21xp5_ASAP7_75t_L g4501 ( 
.A1(n_4357),
.A2(n_4212),
.B(n_4310),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4407),
.Y(n_4502)
);

INVx3_ASAP7_75t_L g4503 ( 
.A(n_4369),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4412),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4365),
.B(n_4247),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_4445),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4375),
.B(n_4248),
.Y(n_4507)
);

BUFx2_ASAP7_75t_L g4508 ( 
.A(n_4397),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4423),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4373),
.B(n_4270),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4373),
.B(n_4297),
.Y(n_4511)
);

INVx2_ASAP7_75t_SL g4512 ( 
.A(n_4322),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4425),
.Y(n_4513)
);

OR2x2_ASAP7_75t_L g4514 ( 
.A(n_4359),
.B(n_4195),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4445),
.Y(n_4515)
);

INVx2_ASAP7_75t_SL g4516 ( 
.A(n_4322),
.Y(n_4516)
);

NOR2x1_ASAP7_75t_SL g4517 ( 
.A(n_4468),
.B(n_4191),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_4447),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4347),
.B(n_4297),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4445),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4405),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4405),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4465),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4323),
.B(n_4339),
.Y(n_4524)
);

INVx1_ASAP7_75t_SL g4525 ( 
.A(n_4453),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4341),
.B(n_4345),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4405),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4455),
.Y(n_4528)
);

INVx3_ASAP7_75t_L g4529 ( 
.A(n_4328),
.Y(n_4529)
);

INVx3_ASAP7_75t_L g4530 ( 
.A(n_4363),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_4361),
.B(n_4195),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_4455),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4451),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4462),
.Y(n_4534)
);

INVx1_ASAP7_75t_SL g4535 ( 
.A(n_4325),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4455),
.Y(n_4536)
);

INVxp67_ASAP7_75t_L g4537 ( 
.A(n_4340),
.Y(n_4537)
);

INVx3_ASAP7_75t_L g4538 ( 
.A(n_4376),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4443),
.B(n_4195),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4374),
.B(n_4191),
.Y(n_4540)
);

INVx3_ASAP7_75t_L g4541 ( 
.A(n_4376),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4438),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4399),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4418),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4378),
.B(n_4173),
.Y(n_4545)
);

BUFx4f_ASAP7_75t_SL g4546 ( 
.A(n_4379),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4390),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_4376),
.Y(n_4548)
);

OR2x2_ASAP7_75t_L g4549 ( 
.A(n_4427),
.B(n_4284),
.Y(n_4549)
);

BUFx6f_ASAP7_75t_L g4550 ( 
.A(n_4356),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4403),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4454),
.B(n_4277),
.Y(n_4552)
);

AOI21x1_ASAP7_75t_L g4553 ( 
.A1(n_4450),
.A2(n_4306),
.B(n_4284),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4471),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4456),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4362),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4372),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4410),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_4327),
.A2(n_4284),
.B1(n_534),
.B2(n_535),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4416),
.B(n_4337),
.Y(n_4560)
);

AO21x2_ASAP7_75t_L g4561 ( 
.A1(n_4448),
.A2(n_532),
.B(n_535),
.Y(n_4561)
);

INVx2_ASAP7_75t_SL g4562 ( 
.A(n_4336),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4464),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4464),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4472),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4349),
.B(n_536),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4414),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4353),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4440),
.Y(n_4569)
);

OR2x6_ASAP7_75t_L g4570 ( 
.A(n_4352),
.B(n_536),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4458),
.Y(n_4571)
);

BUFx3_ASAP7_75t_L g4572 ( 
.A(n_4377),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4420),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4348),
.Y(n_4574)
);

AO21x2_ASAP7_75t_L g4575 ( 
.A1(n_4435),
.A2(n_537),
.B(n_538),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4343),
.B(n_537),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4358),
.Y(n_4577)
);

AO21x2_ASAP7_75t_L g4578 ( 
.A1(n_4334),
.A2(n_538),
.B(n_539),
.Y(n_4578)
);

OR2x6_ASAP7_75t_L g4579 ( 
.A(n_4352),
.B(n_539),
.Y(n_4579)
);

BUFx4f_ASAP7_75t_SL g4580 ( 
.A(n_4329),
.Y(n_4580)
);

AOI221xp5_ASAP7_75t_L g4581 ( 
.A1(n_4389),
.A2(n_540),
.B1(n_541),
.B2(n_542),
.C(n_543),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4400),
.B(n_540),
.Y(n_4582)
);

OR2x6_ASAP7_75t_L g4583 ( 
.A(n_4457),
.B(n_541),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4346),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4424),
.Y(n_4585)
);

BUFx3_ASAP7_75t_L g4586 ( 
.A(n_4394),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4392),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_SL g4588 ( 
.A(n_4395),
.B(n_4330),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4457),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4426),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4389),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4335),
.B(n_542),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4396),
.Y(n_4593)
);

OR2x2_ASAP7_75t_L g4594 ( 
.A(n_4344),
.B(n_543),
.Y(n_4594)
);

AO21x2_ASAP7_75t_L g4595 ( 
.A1(n_4430),
.A2(n_544),
.B(n_545),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4421),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4467),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4350),
.B(n_545),
.Y(n_4598)
);

AND2x4_ASAP7_75t_L g4599 ( 
.A(n_4332),
.B(n_546),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4422),
.B(n_546),
.Y(n_4600)
);

OA21x2_ASAP7_75t_L g4601 ( 
.A1(n_4406),
.A2(n_547),
.B(n_548),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4393),
.B(n_549),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4467),
.Y(n_4603)
);

AOI21x1_ASAP7_75t_L g4604 ( 
.A1(n_4366),
.A2(n_550),
.B(n_551),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4333),
.B(n_550),
.Y(n_4605)
);

OAI21x1_ASAP7_75t_L g4606 ( 
.A1(n_4366),
.A2(n_4368),
.B(n_4364),
.Y(n_4606)
);

OR2x6_ASAP7_75t_L g4607 ( 
.A(n_4368),
.B(n_551),
.Y(n_4607)
);

OA21x2_ASAP7_75t_L g4608 ( 
.A1(n_4408),
.A2(n_552),
.B(n_553),
.Y(n_4608)
);

AND2x4_ASAP7_75t_L g4609 ( 
.A(n_4446),
.B(n_552),
.Y(n_4609)
);

AO31x2_ASAP7_75t_L g4610 ( 
.A1(n_4517),
.A2(n_4441),
.A3(n_4461),
.B(n_4404),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4525),
.B(n_4326),
.Y(n_4611)
);

AOI22xp33_ASAP7_75t_L g4612 ( 
.A1(n_4588),
.A2(n_4327),
.B1(n_4324),
.B2(n_4404),
.Y(n_4612)
);

INVx3_ASAP7_75t_L g4613 ( 
.A(n_4530),
.Y(n_4613)
);

AOI22xp33_ASAP7_75t_L g4614 ( 
.A1(n_4588),
.A2(n_4324),
.B1(n_4354),
.B2(n_4355),
.Y(n_4614)
);

OAI22xp5_ASAP7_75t_L g4615 ( 
.A1(n_4598),
.A2(n_4351),
.B1(n_4384),
.B2(n_4459),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4508),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4508),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4507),
.Y(n_4618)
);

OAI221xp5_ASAP7_75t_L g4619 ( 
.A1(n_4495),
.A2(n_4437),
.B1(n_4401),
.B2(n_4470),
.C(n_4431),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4496),
.Y(n_4620)
);

AND2x4_ASAP7_75t_L g4621 ( 
.A(n_4538),
.B(n_4415),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4496),
.Y(n_4622)
);

INVx2_ASAP7_75t_SL g4623 ( 
.A(n_4479),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4497),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4497),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4474),
.Y(n_4626)
);

AO21x2_ASAP7_75t_L g4627 ( 
.A1(n_4511),
.A2(n_4387),
.B(n_4469),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4478),
.Y(n_4628)
);

OR2x2_ASAP7_75t_L g4629 ( 
.A(n_4563),
.B(n_4564),
.Y(n_4629)
);

AND2x4_ASAP7_75t_L g4630 ( 
.A(n_4538),
.B(n_4436),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4535),
.B(n_4433),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4599),
.B(n_4419),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4482),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4507),
.Y(n_4634)
);

AO31x2_ASAP7_75t_L g4635 ( 
.A1(n_4582),
.A2(n_4441),
.A3(n_4461),
.B(n_4419),
.Y(n_4635)
);

INVx1_ASAP7_75t_SL g4636 ( 
.A(n_4546),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4538),
.B(n_4452),
.Y(n_4637)
);

BUFx2_ASAP7_75t_L g4638 ( 
.A(n_4518),
.Y(n_4638)
);

OR2x2_ASAP7_75t_L g4639 ( 
.A(n_4510),
.B(n_4434),
.Y(n_4639)
);

AOI22xp33_ASAP7_75t_L g4640 ( 
.A1(n_4578),
.A2(n_4460),
.B1(n_4367),
.B2(n_4388),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4541),
.B(n_4442),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4541),
.B(n_4417),
.Y(n_4642)
);

OR2x2_ASAP7_75t_L g4643 ( 
.A(n_4589),
.B(n_4466),
.Y(n_4643)
);

INVx1_ASAP7_75t_SL g4644 ( 
.A(n_4580),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4475),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4541),
.B(n_4402),
.Y(n_4646)
);

OR2x2_ASAP7_75t_L g4647 ( 
.A(n_4589),
.B(n_4444),
.Y(n_4647)
);

BUFx6f_ASAP7_75t_L g4648 ( 
.A(n_4473),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4548),
.B(n_4428),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4522),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4548),
.B(n_4360),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4475),
.Y(n_4652)
);

INVx1_ASAP7_75t_SL g4653 ( 
.A(n_4572),
.Y(n_4653)
);

AO31x2_ASAP7_75t_L g4654 ( 
.A1(n_4566),
.A2(n_4409),
.A3(n_4449),
.B(n_4411),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4487),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4475),
.Y(n_4656)
);

OAI21x1_ASAP7_75t_L g4657 ( 
.A1(n_4485),
.A2(n_553),
.B(n_554),
.Y(n_4657)
);

INVx3_ASAP7_75t_L g4658 ( 
.A(n_4530),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4548),
.B(n_554),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4476),
.B(n_555),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4492),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4499),
.Y(n_4662)
);

INVxp67_ASAP7_75t_L g4663 ( 
.A(n_4479),
.Y(n_4663)
);

INVx3_ASAP7_75t_L g4664 ( 
.A(n_4530),
.Y(n_4664)
);

OR2x2_ASAP7_75t_L g4665 ( 
.A(n_4597),
.B(n_555),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4503),
.Y(n_4666)
);

OR2x2_ASAP7_75t_L g4667 ( 
.A(n_4603),
.B(n_556),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4518),
.B(n_557),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4503),
.Y(n_4669)
);

INVx2_ASAP7_75t_SL g4670 ( 
.A(n_4491),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4518),
.B(n_558),
.Y(n_4671)
);

AND2x4_ASAP7_75t_L g4672 ( 
.A(n_4503),
.B(n_558),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4476),
.B(n_559),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4488),
.B(n_559),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4488),
.B(n_560),
.Y(n_4675)
);

BUFx2_ASAP7_75t_L g4676 ( 
.A(n_4529),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4504),
.Y(n_4677)
);

AOI22xp33_ASAP7_75t_SL g4678 ( 
.A1(n_4578),
.A2(n_560),
.B1(n_561),
.B2(n_562),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4509),
.Y(n_4679)
);

NAND2x1p5_ASAP7_75t_L g4680 ( 
.A(n_4604),
.B(n_561),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4491),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4513),
.Y(n_4682)
);

HB1xp67_ASAP7_75t_L g4683 ( 
.A(n_4578),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4533),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4512),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4489),
.B(n_562),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4534),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4489),
.B(n_563),
.Y(n_4688)
);

INVx3_ASAP7_75t_L g4689 ( 
.A(n_4473),
.Y(n_4689)
);

NOR2xp33_ASAP7_75t_SL g4690 ( 
.A(n_4512),
.B(n_564),
.Y(n_4690)
);

BUFx2_ASAP7_75t_L g4691 ( 
.A(n_4529),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4523),
.Y(n_4692)
);

INVx2_ASAP7_75t_SL g4693 ( 
.A(n_4516),
.Y(n_4693)
);

INVx1_ASAP7_75t_SL g4694 ( 
.A(n_4572),
.Y(n_4694)
);

OR2x2_ASAP7_75t_L g4695 ( 
.A(n_4573),
.B(n_564),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4516),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4550),
.Y(n_4697)
);

HB1xp67_ASAP7_75t_L g4698 ( 
.A(n_4514),
.Y(n_4698)
);

BUFx6f_ASAP7_75t_L g4699 ( 
.A(n_4473),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4529),
.B(n_565),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4550),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4599),
.B(n_567),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4550),
.Y(n_4703)
);

INVxp67_ASAP7_75t_SL g4704 ( 
.A(n_4550),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4574),
.B(n_567),
.Y(n_4705)
);

HB1xp67_ASAP7_75t_L g4706 ( 
.A(n_4514),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4542),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4574),
.B(n_568),
.Y(n_4708)
);

INVx2_ASAP7_75t_SL g4709 ( 
.A(n_4528),
.Y(n_4709)
);

INVxp33_ASAP7_75t_L g4710 ( 
.A(n_4473),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4573),
.B(n_568),
.Y(n_4711)
);

INVx3_ASAP7_75t_L g4712 ( 
.A(n_4473),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4528),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4477),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4532),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4532),
.Y(n_4716)
);

BUFx3_ASAP7_75t_L g4717 ( 
.A(n_4562),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4557),
.B(n_569),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4477),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4536),
.B(n_569),
.Y(n_4720)
);

INVxp67_ASAP7_75t_L g4721 ( 
.A(n_4638),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4613),
.B(n_4562),
.Y(n_4722)
);

NOR2x1_ASAP7_75t_L g4723 ( 
.A(n_4717),
.B(n_4605),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4650),
.Y(n_4724)
);

BUFx6f_ASAP7_75t_L g4725 ( 
.A(n_4648),
.Y(n_4725)
);

AND2x4_ASAP7_75t_L g4726 ( 
.A(n_4717),
.B(n_4536),
.Y(n_4726)
);

AND2x2_ASAP7_75t_L g4727 ( 
.A(n_4613),
.B(n_4555),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4650),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_4676),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4698),
.Y(n_4730)
);

HB1xp67_ASAP7_75t_L g4731 ( 
.A(n_4683),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4698),
.Y(n_4732)
);

AO21x2_ASAP7_75t_L g4733 ( 
.A1(n_4683),
.A2(n_4527),
.B(n_4521),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4691),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4613),
.B(n_4555),
.Y(n_4735)
);

HB1xp67_ASAP7_75t_L g4736 ( 
.A(n_4706),
.Y(n_4736)
);

HB1xp67_ASAP7_75t_L g4737 ( 
.A(n_4706),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4620),
.Y(n_4738)
);

BUFx6f_ASAP7_75t_L g4739 ( 
.A(n_4648),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4648),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4622),
.Y(n_4741)
);

AOI22xp33_ASAP7_75t_SL g4742 ( 
.A1(n_4627),
.A2(n_4560),
.B1(n_4606),
.B2(n_4584),
.Y(n_4742)
);

BUFx3_ASAP7_75t_L g4743 ( 
.A(n_4648),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4624),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4625),
.Y(n_4745)
);

NOR2xp33_ASAP7_75t_L g4746 ( 
.A(n_4710),
.B(n_4577),
.Y(n_4746)
);

INVx5_ASAP7_75t_L g4747 ( 
.A(n_4699),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4616),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4658),
.B(n_4493),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4704),
.B(n_4599),
.Y(n_4750)
);

INVx1_ASAP7_75t_SL g4751 ( 
.A(n_4653),
.Y(n_4751)
);

NOR2xp67_ASAP7_75t_L g4752 ( 
.A(n_4658),
.B(n_4537),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_L g4753 ( 
.A(n_4697),
.B(n_4568),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4617),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4658),
.B(n_4493),
.Y(n_4755)
);

BUFx6f_ASAP7_75t_L g4756 ( 
.A(n_4699),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4697),
.B(n_4568),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4664),
.B(n_4494),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4701),
.B(n_4557),
.Y(n_4759)
);

NOR2xp33_ASAP7_75t_L g4760 ( 
.A(n_4710),
.B(n_4577),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4701),
.B(n_4558),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4699),
.B(n_4490),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4629),
.B(n_4591),
.Y(n_4763)
);

NOR2xp33_ASAP7_75t_L g4764 ( 
.A(n_4699),
.B(n_4586),
.Y(n_4764)
);

INVx3_ASAP7_75t_L g4765 ( 
.A(n_4664),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_4689),
.Y(n_4766)
);

AND2x4_ASAP7_75t_SL g4767 ( 
.A(n_4664),
.B(n_4583),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4618),
.Y(n_4768)
);

INVx3_ASAP7_75t_L g4769 ( 
.A(n_4689),
.Y(n_4769)
);

INVx2_ASAP7_75t_SL g4770 ( 
.A(n_4689),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4618),
.B(n_4634),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4694),
.B(n_4494),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4703),
.B(n_4558),
.Y(n_4773)
);

INVxp67_ASAP7_75t_SL g4774 ( 
.A(n_4680),
.Y(n_4774)
);

AND2x4_ASAP7_75t_L g4775 ( 
.A(n_4623),
.B(n_4521),
.Y(n_4775)
);

INVx3_ASAP7_75t_L g4776 ( 
.A(n_4712),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4712),
.Y(n_4777)
);

INVx2_ASAP7_75t_SL g4778 ( 
.A(n_4712),
.Y(n_4778)
);

HB1xp67_ASAP7_75t_L g4779 ( 
.A(n_4634),
.Y(n_4779)
);

NOR2x1_ASAP7_75t_SL g4780 ( 
.A(n_4623),
.B(n_4607),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4670),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4660),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4670),
.Y(n_4783)
);

HB1xp67_ASAP7_75t_L g4784 ( 
.A(n_4610),
.Y(n_4784)
);

BUFx3_ASAP7_75t_L g4785 ( 
.A(n_4673),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4647),
.B(n_4591),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4736),
.Y(n_4787)
);

INVxp67_ASAP7_75t_SL g4788 ( 
.A(n_4752),
.Y(n_4788)
);

HB1xp67_ASAP7_75t_L g4789 ( 
.A(n_4736),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4765),
.Y(n_4790)
);

NOR2x1_ASAP7_75t_L g4791 ( 
.A(n_4765),
.B(n_4703),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4737),
.Y(n_4792)
);

OR2x6_ASAP7_75t_L g4793 ( 
.A(n_4725),
.B(n_4693),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4722),
.B(n_4637),
.Y(n_4794)
);

AND2x4_ASAP7_75t_L g4795 ( 
.A(n_4747),
.B(n_4693),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4751),
.B(n_4637),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4737),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4779),
.Y(n_4798)
);

OAI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4742),
.A2(n_4612),
.B(n_4614),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4779),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4729),
.B(n_4611),
.Y(n_4801)
);

AND2x2_ASAP7_75t_SL g4802 ( 
.A(n_4767),
.B(n_4612),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4750),
.B(n_4643),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4747),
.Y(n_4804)
);

AND2x4_ASAP7_75t_L g4805 ( 
.A(n_4747),
.B(n_4709),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4726),
.B(n_4646),
.Y(n_4806)
);

BUFx3_ASAP7_75t_L g4807 ( 
.A(n_4726),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4747),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4731),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4731),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4726),
.B(n_4646),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4734),
.B(n_4663),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_4723),
.B(n_4678),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4772),
.B(n_4641),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4724),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4734),
.B(n_4681),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4785),
.B(n_4681),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4728),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4727),
.B(n_4641),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4730),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4732),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_SL g4822 ( 
.A(n_4785),
.B(n_4632),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4725),
.Y(n_4823)
);

INVx3_ASAP7_75t_L g4824 ( 
.A(n_4725),
.Y(n_4824)
);

NOR2xp33_ASAP7_75t_L g4825 ( 
.A(n_4764),
.B(n_4644),
.Y(n_4825)
);

INVx2_ASAP7_75t_SL g4826 ( 
.A(n_4725),
.Y(n_4826)
);

AND2x4_ASAP7_75t_L g4827 ( 
.A(n_4778),
.B(n_4709),
.Y(n_4827)
);

OR2x2_ASAP7_75t_L g4828 ( 
.A(n_4786),
.B(n_4627),
.Y(n_4828)
);

INVx2_ASAP7_75t_L g4829 ( 
.A(n_4739),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4735),
.B(n_4649),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4721),
.B(n_4685),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4771),
.Y(n_4832)
);

OR2x2_ASAP7_75t_L g4833 ( 
.A(n_4763),
.B(n_4610),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4733),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4749),
.B(n_4649),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4739),
.Y(n_4836)
);

AND2x4_ASAP7_75t_SL g4837 ( 
.A(n_4739),
.B(n_4685),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4755),
.B(n_4630),
.Y(n_4838)
);

AND2x4_ASAP7_75t_SL g4839 ( 
.A(n_4739),
.B(n_4696),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4733),
.Y(n_4840)
);

INVx2_ASAP7_75t_L g4841 ( 
.A(n_4756),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4780),
.B(n_4630),
.Y(n_4842)
);

OR2x2_ASAP7_75t_L g4843 ( 
.A(n_4789),
.B(n_4784),
.Y(n_4843)
);

AND2x4_ASAP7_75t_SL g4844 ( 
.A(n_4838),
.B(n_4756),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4806),
.B(n_4767),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4798),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4800),
.Y(n_4847)
);

AOI22xp5_ASAP7_75t_L g4848 ( 
.A1(n_4799),
.A2(n_4614),
.B1(n_4560),
.B2(n_4619),
.Y(n_4848)
);

AND2x4_ASAP7_75t_L g4849 ( 
.A(n_4807),
.B(n_4778),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4806),
.B(n_4811),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4811),
.B(n_4758),
.Y(n_4851)
);

AND2x2_ASAP7_75t_L g4852 ( 
.A(n_4794),
.B(n_4758),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4794),
.B(n_4758),
.Y(n_4853)
);

INVx4_ASAP7_75t_L g4854 ( 
.A(n_4824),
.Y(n_4854)
);

NOR2xp67_ASAP7_75t_L g4855 ( 
.A(n_4842),
.B(n_4769),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4787),
.Y(n_4856)
);

AND2x4_ASAP7_75t_L g4857 ( 
.A(n_4807),
.B(n_4805),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4805),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4814),
.B(n_4774),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4834),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4814),
.B(n_4781),
.Y(n_4861)
);

INVxp67_ASAP7_75t_L g4862 ( 
.A(n_4842),
.Y(n_4862)
);

NAND4xp25_ASAP7_75t_L g4863 ( 
.A(n_4825),
.B(n_4762),
.C(n_4764),
.D(n_4760),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4840),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4792),
.Y(n_4865)
);

HB1xp67_ASAP7_75t_L g4866 ( 
.A(n_4805),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4838),
.B(n_4781),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4827),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4797),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4827),
.Y(n_4870)
);

AND2x4_ASAP7_75t_L g4871 ( 
.A(n_4827),
.B(n_4743),
.Y(n_4871)
);

AND2x4_ASAP7_75t_L g4872 ( 
.A(n_4795),
.B(n_4743),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4809),
.Y(n_4873)
);

OR2x6_ASAP7_75t_SL g4874 ( 
.A(n_4796),
.B(n_4740),
.Y(n_4874)
);

INVx2_ASAP7_75t_L g4875 ( 
.A(n_4795),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4835),
.B(n_4783),
.Y(n_4876)
);

INVxp67_ASAP7_75t_SL g4877 ( 
.A(n_4791),
.Y(n_4877)
);

OR2x2_ASAP7_75t_L g4878 ( 
.A(n_4828),
.B(n_4784),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4795),
.Y(n_4879)
);

INVx3_ASAP7_75t_L g4880 ( 
.A(n_4793),
.Y(n_4880)
);

BUFx2_ASAP7_75t_L g4881 ( 
.A(n_4793),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4835),
.B(n_4783),
.Y(n_4882)
);

NAND2x1p5_ASAP7_75t_L g4883 ( 
.A(n_4824),
.B(n_4756),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4819),
.B(n_4774),
.Y(n_4884)
);

INVx2_ASAP7_75t_SL g4885 ( 
.A(n_4837),
.Y(n_4885)
);

OR2x2_ASAP7_75t_L g4886 ( 
.A(n_4833),
.B(n_4782),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4819),
.B(n_4696),
.Y(n_4887)
);

AND2x4_ASAP7_75t_SL g4888 ( 
.A(n_4793),
.B(n_4756),
.Y(n_4888)
);

OR2x2_ASAP7_75t_L g4889 ( 
.A(n_4822),
.B(n_4753),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4830),
.B(n_4801),
.Y(n_4890)
);

BUFx3_ASAP7_75t_L g4891 ( 
.A(n_4837),
.Y(n_4891)
);

AOI22xp5_ASAP7_75t_L g4892 ( 
.A1(n_4848),
.A2(n_4813),
.B1(n_4822),
.B2(n_4802),
.Y(n_4892)
);

OR2x2_ASAP7_75t_L g4893 ( 
.A(n_4859),
.B(n_4817),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4890),
.B(n_4830),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4858),
.Y(n_4895)
);

OR2x2_ASAP7_75t_L g4896 ( 
.A(n_4884),
.B(n_4816),
.Y(n_4896)
);

INVx2_ASAP7_75t_L g4897 ( 
.A(n_4857),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4889),
.B(n_4831),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4890),
.B(n_4813),
.Y(n_4899)
);

OR2x2_ASAP7_75t_L g4900 ( 
.A(n_4861),
.B(n_4812),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4850),
.B(n_4801),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4850),
.B(n_4802),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4845),
.B(n_4825),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4845),
.B(n_4788),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4852),
.B(n_4630),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4861),
.B(n_4803),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4876),
.B(n_4833),
.Y(n_4907)
);

AND2x2_ASAP7_75t_SL g4908 ( 
.A(n_4844),
.B(n_4839),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_SL g4909 ( 
.A(n_4857),
.B(n_4690),
.Y(n_4909)
);

AND2x4_ASAP7_75t_L g4910 ( 
.A(n_4857),
.B(n_4839),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4871),
.B(n_4826),
.Y(n_4911)
);

INVx1_ASAP7_75t_SL g4912 ( 
.A(n_4852),
.Y(n_4912)
);

AND2x4_ASAP7_75t_L g4913 ( 
.A(n_4871),
.B(n_4826),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4866),
.B(n_4746),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4853),
.B(n_4636),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4853),
.B(n_4631),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4843),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4867),
.B(n_4642),
.Y(n_4918)
);

OR2x2_ASAP7_75t_L g4919 ( 
.A(n_4876),
.B(n_4757),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4882),
.B(n_4832),
.Y(n_4920)
);

NOR2xp33_ASAP7_75t_L g4921 ( 
.A(n_4874),
.B(n_4820),
.Y(n_4921)
);

OR2x2_ASAP7_75t_L g4922 ( 
.A(n_4882),
.B(n_4759),
.Y(n_4922)
);

OR2x2_ASAP7_75t_L g4923 ( 
.A(n_4863),
.B(n_4761),
.Y(n_4923)
);

INVx2_ASAP7_75t_SL g4924 ( 
.A(n_4844),
.Y(n_4924)
);

OR2x2_ASAP7_75t_L g4925 ( 
.A(n_4887),
.B(n_4773),
.Y(n_4925)
);

NAND2x1_ASAP7_75t_L g4926 ( 
.A(n_4871),
.B(n_4793),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4843),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4867),
.B(n_4642),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4883),
.Y(n_4929)
);

OR2x2_ASAP7_75t_L g4930 ( 
.A(n_4887),
.B(n_4748),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4912),
.B(n_4885),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4912),
.B(n_4874),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_SL g4933 ( 
.A(n_4910),
.B(n_4872),
.Y(n_4933)
);

OR2x2_ASAP7_75t_L g4934 ( 
.A(n_4914),
.B(n_4899),
.Y(n_4934)
);

AND2x2_ASAP7_75t_L g4935 ( 
.A(n_4901),
.B(n_4851),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4894),
.B(n_4868),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4904),
.B(n_4851),
.Y(n_4937)
);

INVx1_ASAP7_75t_SL g4938 ( 
.A(n_4908),
.Y(n_4938)
);

OAI22xp5_ASAP7_75t_L g4939 ( 
.A1(n_4892),
.A2(n_4877),
.B1(n_4639),
.B2(n_4621),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4897),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4918),
.B(n_4885),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4897),
.Y(n_4942)
);

HB1xp67_ASAP7_75t_L g4943 ( 
.A(n_4926),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4928),
.B(n_4862),
.Y(n_4944)
);

OR2x2_ASAP7_75t_L g4945 ( 
.A(n_4914),
.B(n_4870),
.Y(n_4945)
);

AND2x4_ASAP7_75t_L g4946 ( 
.A(n_4910),
.B(n_4872),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4920),
.Y(n_4947)
);

INVx1_ASAP7_75t_SL g4948 ( 
.A(n_4908),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4911),
.Y(n_4949)
);

HB1xp67_ASAP7_75t_L g4950 ( 
.A(n_4911),
.Y(n_4950)
);

NOR2x1_ASAP7_75t_L g4951 ( 
.A(n_4913),
.B(n_4891),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4907),
.Y(n_4952)
);

OR2x2_ASAP7_75t_L g4953 ( 
.A(n_4899),
.B(n_4868),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4895),
.B(n_4849),
.Y(n_4954)
);

OR2x2_ASAP7_75t_L g4955 ( 
.A(n_4906),
.B(n_4875),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_4913),
.B(n_4849),
.Y(n_4956)
);

OR2x2_ASAP7_75t_L g4957 ( 
.A(n_4900),
.B(n_4875),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4925),
.Y(n_4958)
);

AOI21xp5_ASAP7_75t_L g4959 ( 
.A1(n_4909),
.A2(n_4760),
.B(n_4746),
.Y(n_4959)
);

OR2x2_ASAP7_75t_L g4960 ( 
.A(n_4919),
.B(n_4879),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4915),
.B(n_4891),
.Y(n_4961)
);

AOI22xp5_ASAP7_75t_L g4962 ( 
.A1(n_4892),
.A2(n_4621),
.B1(n_4762),
.B2(n_4651),
.Y(n_4962)
);

OR2x2_ASAP7_75t_L g4963 ( 
.A(n_4922),
.B(n_4879),
.Y(n_4963)
);

NAND3xp33_ASAP7_75t_SL g4964 ( 
.A(n_4902),
.B(n_4881),
.C(n_4883),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4903),
.B(n_4855),
.Y(n_4965)
);

INVx2_ASAP7_75t_L g4966 ( 
.A(n_4905),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4916),
.B(n_4872),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4950),
.B(n_4849),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4949),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_L g4970 ( 
.A(n_4946),
.B(n_4924),
.Y(n_4970)
);

OAI22xp33_ASAP7_75t_L g4971 ( 
.A1(n_4962),
.A2(n_4549),
.B1(n_4607),
.B2(n_4579),
.Y(n_4971)
);

INVx3_ASAP7_75t_L g4972 ( 
.A(n_4946),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4931),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4954),
.Y(n_4974)
);

INVxp67_ASAP7_75t_L g4975 ( 
.A(n_4951),
.Y(n_4975)
);

NOR4xp25_ASAP7_75t_L g4976 ( 
.A(n_4932),
.B(n_4921),
.C(n_4927),
.D(n_4917),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4937),
.B(n_4967),
.Y(n_4977)
);

NOR2xp33_ASAP7_75t_L g4978 ( 
.A(n_4933),
.B(n_4909),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4961),
.B(n_4929),
.Y(n_4979)
);

OR2x2_ASAP7_75t_L g4980 ( 
.A(n_4932),
.B(n_4930),
.Y(n_4980)
);

O2A1O1Ixp33_ASAP7_75t_L g4981 ( 
.A1(n_4939),
.A2(n_4921),
.B(n_4878),
.C(n_4880),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4954),
.Y(n_4982)
);

AOI211xp5_ASAP7_75t_SL g4983 ( 
.A1(n_4939),
.A2(n_4880),
.B(n_4898),
.C(n_4893),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4936),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4936),
.Y(n_4985)
);

NAND4xp25_ASAP7_75t_L g4986 ( 
.A(n_4959),
.B(n_4923),
.C(n_4896),
.D(n_4865),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4935),
.B(n_4888),
.Y(n_4987)
);

INVxp67_ASAP7_75t_L g4988 ( 
.A(n_4943),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4955),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4965),
.B(n_4888),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4956),
.Y(n_4991)
);

AOI221xp5_ASAP7_75t_L g4992 ( 
.A1(n_4964),
.A2(n_4818),
.B1(n_4815),
.B2(n_4754),
.C(n_4821),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4953),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4944),
.B(n_4621),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4966),
.B(n_4880),
.Y(n_4995)
);

OR2x6_ASAP7_75t_L g4996 ( 
.A(n_4957),
.B(n_4854),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4938),
.B(n_4740),
.Y(n_4997)
);

INVxp67_ASAP7_75t_L g4998 ( 
.A(n_4972),
.Y(n_4998)
);

NAND2xp5_ASAP7_75t_L g4999 ( 
.A(n_4972),
.B(n_4938),
.Y(n_4999)
);

INVx1_ASAP7_75t_SL g5000 ( 
.A(n_4994),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4987),
.B(n_4948),
.Y(n_5001)
);

INVx1_ASAP7_75t_SL g5002 ( 
.A(n_4968),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4996),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4979),
.B(n_4948),
.Y(n_5004)
);

OR2x2_ASAP7_75t_L g5005 ( 
.A(n_4970),
.B(n_4941),
.Y(n_5005)
);

NAND2xp5_ASAP7_75t_L g5006 ( 
.A(n_4995),
.B(n_4940),
.Y(n_5006)
);

HB1xp67_ASAP7_75t_L g5007 ( 
.A(n_4996),
.Y(n_5007)
);

HB1xp67_ASAP7_75t_L g5008 ( 
.A(n_4996),
.Y(n_5008)
);

OR2x2_ASAP7_75t_L g5009 ( 
.A(n_4997),
.B(n_4963),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4975),
.B(n_4942),
.Y(n_5010)
);

HB1xp67_ASAP7_75t_L g5011 ( 
.A(n_4990),
.Y(n_5011)
);

NAND2x1p5_ASAP7_75t_L g5012 ( 
.A(n_4989),
.B(n_4854),
.Y(n_5012)
);

NAND2x1_ASAP7_75t_L g5013 ( 
.A(n_4993),
.B(n_4769),
.Y(n_5013)
);

AOI21xp33_ASAP7_75t_L g5014 ( 
.A1(n_4981),
.A2(n_4934),
.B(n_4960),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4980),
.Y(n_5015)
);

OAI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4988),
.A2(n_4947),
.B(n_4945),
.Y(n_5016)
);

INVx1_ASAP7_75t_SL g5017 ( 
.A(n_4977),
.Y(n_5017)
);

HB1xp67_ASAP7_75t_L g5018 ( 
.A(n_4973),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_5011),
.B(n_5000),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_5012),
.Y(n_5020)
);

OAI22xp33_ASAP7_75t_L g5021 ( 
.A1(n_4999),
.A2(n_4983),
.B1(n_4770),
.B2(n_4645),
.Y(n_5021)
);

O2A1O1Ixp33_ASAP7_75t_L g5022 ( 
.A1(n_5014),
.A2(n_4976),
.B(n_4878),
.C(n_4860),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_5012),
.Y(n_5023)
);

OAI221xp5_ASAP7_75t_L g5024 ( 
.A1(n_4998),
.A2(n_4992),
.B1(n_4976),
.B2(n_4978),
.C(n_4986),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_5007),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_5008),
.B(n_4823),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_5004),
.Y(n_5027)
);

OAI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_5001),
.A2(n_4969),
.B1(n_4645),
.B2(n_4656),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_5013),
.Y(n_5029)
);

OAI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_5016),
.A2(n_4952),
.B(n_4974),
.Y(n_5030)
);

OAI22xp33_ASAP7_75t_L g5031 ( 
.A1(n_5002),
.A2(n_4652),
.B1(n_4666),
.B2(n_4656),
.Y(n_5031)
);

AOI31xp33_ASAP7_75t_L g5032 ( 
.A1(n_5009),
.A2(n_4982),
.A3(n_4985),
.B(n_4984),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_5018),
.Y(n_5033)
);

INVxp67_ASAP7_75t_L g5034 ( 
.A(n_5006),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_5005),
.Y(n_5035)
);

NOR3xp33_ASAP7_75t_L g5036 ( 
.A(n_5024),
.B(n_4986),
.C(n_5015),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_5019),
.B(n_4856),
.Y(n_5037)
);

OAI22xp33_ASAP7_75t_L g5038 ( 
.A1(n_5032),
.A2(n_4652),
.B1(n_4669),
.B2(n_4666),
.Y(n_5038)
);

AOI21xp33_ASAP7_75t_SL g5039 ( 
.A1(n_5021),
.A2(n_4958),
.B(n_5003),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_5031),
.B(n_4869),
.Y(n_5040)
);

OAI22xp33_ASAP7_75t_L g5041 ( 
.A1(n_5032),
.A2(n_4669),
.B1(n_4776),
.B2(n_5017),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_5026),
.Y(n_5042)
);

AOI321xp33_ASAP7_75t_L g5043 ( 
.A1(n_5028),
.A2(n_4991),
.A3(n_5010),
.B1(n_4873),
.B2(n_4847),
.C(n_4846),
.Y(n_5043)
);

OR2x2_ASAP7_75t_L g5044 ( 
.A(n_5025),
.B(n_4886),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_5029),
.B(n_4854),
.Y(n_5045)
);

AND2x4_ASAP7_75t_L g5046 ( 
.A(n_5020),
.B(n_4823),
.Y(n_5046)
);

NOR2xp33_ASAP7_75t_L g5047 ( 
.A(n_5033),
.B(n_4971),
.Y(n_5047)
);

AOI22xp33_ASAP7_75t_L g5048 ( 
.A1(n_5035),
.A2(n_4775),
.B1(n_4776),
.B2(n_4790),
.Y(n_5048)
);

AOI21xp33_ASAP7_75t_L g5049 ( 
.A1(n_5022),
.A2(n_4808),
.B(n_4804),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_5023),
.Y(n_5050)
);

OR2x2_ASAP7_75t_L g5051 ( 
.A(n_5030),
.B(n_4886),
.Y(n_5051)
);

OAI221xp5_ASAP7_75t_L g5052 ( 
.A1(n_5034),
.A2(n_4790),
.B1(n_4808),
.B2(n_4804),
.C(n_4777),
.Y(n_5052)
);

NOR2x1_ASAP7_75t_L g5053 ( 
.A(n_5027),
.B(n_4824),
.Y(n_5053)
);

AOI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_5019),
.A2(n_4775),
.B1(n_4777),
.B2(n_4766),
.Y(n_5054)
);

INVx1_ASAP7_75t_SL g5055 ( 
.A(n_5019),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_5048),
.B(n_4829),
.Y(n_5056)
);

OR2x2_ASAP7_75t_L g5057 ( 
.A(n_5044),
.B(n_4829),
.Y(n_5057)
);

NOR2xp33_ASAP7_75t_L g5058 ( 
.A(n_5052),
.B(n_4836),
.Y(n_5058)
);

XNOR2x1_ASAP7_75t_L g5059 ( 
.A(n_5055),
.B(n_4860),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_5054),
.B(n_4836),
.Y(n_5060)
);

A2O1A1Ixp33_ASAP7_75t_L g5061 ( 
.A1(n_5049),
.A2(n_4841),
.B(n_4810),
.C(n_4766),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5038),
.B(n_4841),
.Y(n_5062)
);

NAND3xp33_ASAP7_75t_L g5063 ( 
.A(n_5043),
.B(n_4864),
.C(n_4768),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5051),
.Y(n_5064)
);

OAI221xp5_ASAP7_75t_L g5065 ( 
.A1(n_5036),
.A2(n_4864),
.B1(n_4738),
.B2(n_4745),
.C(n_4744),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_5046),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_5046),
.B(n_4626),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_SL g5068 ( 
.A(n_5041),
.B(n_4775),
.Y(n_5068)
);

OAI222xp33_ASAP7_75t_L g5069 ( 
.A1(n_5050),
.A2(n_4741),
.B1(n_4713),
.B2(n_4716),
.C1(n_4715),
.C2(n_4527),
.Y(n_5069)
);

INVxp67_ASAP7_75t_SL g5070 ( 
.A(n_5053),
.Y(n_5070)
);

AOI22xp33_ASAP7_75t_L g5071 ( 
.A1(n_5047),
.A2(n_5042),
.B1(n_4715),
.B2(n_4716),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_5037),
.B(n_4713),
.Y(n_5072)
);

NOR2xp33_ASAP7_75t_L g5073 ( 
.A(n_5039),
.B(n_4586),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5045),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_5040),
.B(n_4651),
.Y(n_5075)
);

INVx1_ASAP7_75t_SL g5076 ( 
.A(n_5044),
.Y(n_5076)
);

INVxp67_ASAP7_75t_L g5077 ( 
.A(n_5044),
.Y(n_5077)
);

OAI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_5048),
.A2(n_4500),
.B1(n_4502),
.B2(n_4498),
.Y(n_5078)
);

OAI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_5054),
.A2(n_4659),
.B(n_4668),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_5048),
.B(n_4543),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_5044),
.Y(n_5081)
);

INVx1_ASAP7_75t_SL g5082 ( 
.A(n_5044),
.Y(n_5082)
);

NOR2xp33_ASAP7_75t_SL g5083 ( 
.A(n_5055),
.B(n_4659),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5054),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_5083),
.B(n_4498),
.Y(n_5085)
);

OAI22xp5_ASAP7_75t_L g5086 ( 
.A1(n_5071),
.A2(n_4502),
.B1(n_4506),
.B2(n_4500),
.Y(n_5086)
);

OR2x2_ASAP7_75t_L g5087 ( 
.A(n_5057),
.B(n_5076),
.Y(n_5087)
);

OAI221xp5_ASAP7_75t_L g5088 ( 
.A1(n_5083),
.A2(n_5061),
.B1(n_5079),
.B2(n_5073),
.C(n_5076),
.Y(n_5088)
);

AOI22xp5_ASAP7_75t_L g5089 ( 
.A1(n_5082),
.A2(n_4672),
.B1(n_4700),
.B2(n_4671),
.Y(n_5089)
);

AOI221x1_ASAP7_75t_L g5090 ( 
.A1(n_5084),
.A2(n_4672),
.B1(n_4702),
.B2(n_4673),
.C(n_4714),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_5066),
.B(n_4506),
.Y(n_5091)
);

AOI211xp5_ASAP7_75t_L g5092 ( 
.A1(n_5065),
.A2(n_4674),
.B(n_4675),
.C(n_4660),
.Y(n_5092)
);

AOI22xp5_ASAP7_75t_L g5093 ( 
.A1(n_5082),
.A2(n_4672),
.B1(n_4673),
.B2(n_4720),
.Y(n_5093)
);

NAND2x1_ASAP7_75t_L g5094 ( 
.A(n_5067),
.B(n_4720),
.Y(n_5094)
);

OAI221xp5_ASAP7_75t_SL g5095 ( 
.A1(n_5077),
.A2(n_4667),
.B1(n_4665),
.B2(n_4718),
.C(n_4695),
.Y(n_5095)
);

OAI221xp5_ASAP7_75t_L g5096 ( 
.A1(n_5070),
.A2(n_4711),
.B1(n_4719),
.B2(n_4682),
.C(n_4707),
.Y(n_5096)
);

AOI22xp5_ASAP7_75t_L g5097 ( 
.A1(n_5081),
.A2(n_4708),
.B1(n_4705),
.B2(n_4675),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_L g5098 ( 
.A(n_5056),
.B(n_4515),
.Y(n_5098)
);

OAI221xp5_ASAP7_75t_L g5099 ( 
.A1(n_5063),
.A2(n_4692),
.B1(n_4628),
.B2(n_4687),
.C(n_4633),
.Y(n_5099)
);

OAI21xp33_ASAP7_75t_L g5100 ( 
.A1(n_5075),
.A2(n_4688),
.B(n_4686),
.Y(n_5100)
);

AOI221xp5_ASAP7_75t_L g5101 ( 
.A1(n_5078),
.A2(n_4688),
.B1(n_4686),
.B2(n_4674),
.C(n_4677),
.Y(n_5101)
);

AOI21xp5_ASAP7_75t_L g5102 ( 
.A1(n_5068),
.A2(n_5080),
.B(n_5064),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5062),
.Y(n_5103)
);

OAI221xp5_ASAP7_75t_L g5104 ( 
.A1(n_5058),
.A2(n_4684),
.B1(n_4655),
.B2(n_4679),
.C(n_4662),
.Y(n_5104)
);

AO21x1_ASAP7_75t_L g5105 ( 
.A1(n_5059),
.A2(n_4531),
.B(n_4520),
.Y(n_5105)
);

AOI221xp5_ASAP7_75t_L g5106 ( 
.A1(n_5069),
.A2(n_4661),
.B1(n_4615),
.B2(n_4515),
.C(n_4520),
.Y(n_5106)
);

AOI221xp5_ASAP7_75t_L g5107 ( 
.A1(n_5060),
.A2(n_4539),
.B1(n_4576),
.B2(n_4596),
.C(n_4602),
.Y(n_5107)
);

AOI222xp33_ASAP7_75t_L g5108 ( 
.A1(n_5072),
.A2(n_4576),
.B1(n_4602),
.B2(n_4592),
.C1(n_4539),
.C2(n_4587),
.Y(n_5108)
);

AOI21xp33_ASAP7_75t_SL g5109 ( 
.A1(n_5074),
.A2(n_4680),
.B(n_4657),
.Y(n_5109)
);

O2A1O1Ixp33_ASAP7_75t_L g5110 ( 
.A1(n_5068),
.A2(n_4531),
.B(n_4594),
.C(n_4583),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5057),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_5057),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_5083),
.B(n_4556),
.Y(n_5113)
);

AOI221xp5_ASAP7_75t_L g5114 ( 
.A1(n_5078),
.A2(n_4592),
.B1(n_4587),
.B2(n_4581),
.C(n_4590),
.Y(n_5114)
);

O2A1O1Ixp33_ASAP7_75t_L g5115 ( 
.A1(n_5068),
.A2(n_4594),
.B(n_4583),
.C(n_4607),
.Y(n_5115)
);

AOI311xp33_ASAP7_75t_L g5116 ( 
.A1(n_5088),
.A2(n_4565),
.A3(n_4593),
.B(n_4585),
.C(n_4519),
.Y(n_5116)
);

OAI21xp5_ASAP7_75t_L g5117 ( 
.A1(n_5102),
.A2(n_4657),
.B(n_4485),
.Y(n_5117)
);

O2A1O1Ixp33_ASAP7_75t_L g5118 ( 
.A1(n_5087),
.A2(n_4583),
.B(n_4607),
.C(n_4570),
.Y(n_5118)
);

AOI221x1_ASAP7_75t_L g5119 ( 
.A1(n_5111),
.A2(n_4556),
.B1(n_4483),
.B2(n_4480),
.C(n_4501),
.Y(n_5119)
);

NAND4xp25_ASAP7_75t_L g5120 ( 
.A(n_5089),
.B(n_4640),
.C(n_4559),
.D(n_4600),
.Y(n_5120)
);

NOR2xp33_ASAP7_75t_SL g5121 ( 
.A(n_5112),
.B(n_4569),
.Y(n_5121)
);

AOI221x1_ASAP7_75t_L g5122 ( 
.A1(n_5103),
.A2(n_4480),
.B1(n_4483),
.B2(n_4567),
.C(n_4540),
.Y(n_5122)
);

AOI221xp5_ASAP7_75t_L g5123 ( 
.A1(n_5086),
.A2(n_4640),
.B1(n_4481),
.B2(n_4549),
.C(n_4575),
.Y(n_5123)
);

OAI22xp5_ASAP7_75t_L g5124 ( 
.A1(n_5093),
.A2(n_4554),
.B1(n_4547),
.B2(n_4551),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_5097),
.B(n_4610),
.Y(n_5125)
);

NOR2x1_ASAP7_75t_L g5126 ( 
.A(n_5091),
.B(n_4481),
.Y(n_5126)
);

AOI21xp5_ASAP7_75t_SL g5127 ( 
.A1(n_5085),
.A2(n_4579),
.B(n_4570),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5113),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_5094),
.A2(n_4481),
.B(n_4484),
.Y(n_5129)
);

AOI221x1_ASAP7_75t_L g5130 ( 
.A1(n_5098),
.A2(n_5100),
.B1(n_5105),
.B2(n_5109),
.C(n_5090),
.Y(n_5130)
);

AOI221xp5_ASAP7_75t_L g5131 ( 
.A1(n_5110),
.A2(n_4575),
.B1(n_4595),
.B2(n_4561),
.C(n_4551),
.Y(n_5131)
);

NAND4xp75_ASAP7_75t_L g5132 ( 
.A(n_5106),
.B(n_5101),
.C(n_5107),
.D(n_5114),
.Y(n_5132)
);

NAND3xp33_ASAP7_75t_L g5133 ( 
.A(n_5092),
.B(n_4579),
.C(n_4570),
.Y(n_5133)
);

AOI211xp5_ASAP7_75t_L g5134 ( 
.A1(n_5096),
.A2(n_4606),
.B(n_4598),
.C(n_4545),
.Y(n_5134)
);

NOR3xp33_ASAP7_75t_L g5135 ( 
.A(n_5095),
.B(n_4604),
.C(n_4571),
.Y(n_5135)
);

NOR2xp33_ASAP7_75t_L g5136 ( 
.A(n_5099),
.B(n_4547),
.Y(n_5136)
);

AOI21xp33_ASAP7_75t_L g5137 ( 
.A1(n_5115),
.A2(n_4575),
.B(n_4595),
.Y(n_5137)
);

AOI22xp33_ASAP7_75t_SL g5138 ( 
.A1(n_5104),
.A2(n_5108),
.B1(n_4595),
.B2(n_4561),
.Y(n_5138)
);

AND2x2_ASAP7_75t_L g5139 ( 
.A(n_5093),
.B(n_4610),
.Y(n_5139)
);

O2A1O1Ixp33_ASAP7_75t_L g5140 ( 
.A1(n_5087),
.A2(n_4570),
.B(n_4579),
.C(n_4561),
.Y(n_5140)
);

AOI322xp5_ASAP7_75t_L g5141 ( 
.A1(n_5100),
.A2(n_4609),
.A3(n_4545),
.B1(n_4554),
.B2(n_4635),
.C1(n_4524),
.C2(n_4526),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5093),
.Y(n_5142)
);

OAI222xp33_ASAP7_75t_L g5143 ( 
.A1(n_5088),
.A2(n_4540),
.B1(n_4544),
.B2(n_4526),
.C1(n_4524),
.C2(n_4609),
.Y(n_5143)
);

AOI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_5102),
.A2(n_4484),
.B(n_4552),
.Y(n_5144)
);

NAND3xp33_ASAP7_75t_SL g5145 ( 
.A(n_5121),
.B(n_4552),
.C(n_4505),
.Y(n_5145)
);

NOR2xp33_ASAP7_75t_L g5146 ( 
.A(n_5139),
.B(n_4484),
.Y(n_5146)
);

OAI211xp5_ASAP7_75t_L g5147 ( 
.A1(n_5130),
.A2(n_4608),
.B(n_4601),
.C(n_4553),
.Y(n_5147)
);

AOI211xp5_ASAP7_75t_L g5148 ( 
.A1(n_5142),
.A2(n_4609),
.B(n_4505),
.C(n_573),
.Y(n_5148)
);

OAI22xp33_ASAP7_75t_L g5149 ( 
.A1(n_5133),
.A2(n_4608),
.B1(n_4601),
.B2(n_4553),
.Y(n_5149)
);

AOI211xp5_ASAP7_75t_L g5150 ( 
.A1(n_5136),
.A2(n_571),
.B(n_572),
.C(n_574),
.Y(n_5150)
);

OAI211xp5_ASAP7_75t_SL g5151 ( 
.A1(n_5128),
.A2(n_4635),
.B(n_572),
.C(n_574),
.Y(n_5151)
);

AOI21xp33_ASAP7_75t_L g5152 ( 
.A1(n_5118),
.A2(n_4486),
.B(n_575),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_5125),
.B(n_4635),
.Y(n_5153)
);

AOI221xp5_ASAP7_75t_L g5154 ( 
.A1(n_5137),
.A2(n_4486),
.B1(n_4635),
.B2(n_4654),
.C(n_577),
.Y(n_5154)
);

AOI22xp5_ASAP7_75t_L g5155 ( 
.A1(n_5135),
.A2(n_4486),
.B1(n_4608),
.B2(n_4601),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_5127),
.Y(n_5156)
);

OAI31xp33_ASAP7_75t_L g5157 ( 
.A1(n_5143),
.A2(n_4654),
.A3(n_575),
.B(n_576),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_5134),
.B(n_4654),
.Y(n_5158)
);

AOI21xp5_ASAP7_75t_L g5159 ( 
.A1(n_5126),
.A2(n_4654),
.B(n_576),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5132),
.Y(n_5160)
);

AOI211xp5_ASAP7_75t_SL g5161 ( 
.A1(n_5144),
.A2(n_571),
.B(n_577),
.C(n_578),
.Y(n_5161)
);

OAI211xp5_ASAP7_75t_L g5162 ( 
.A1(n_5116),
.A2(n_578),
.B(n_579),
.C(n_580),
.Y(n_5162)
);

A2O1A1Ixp33_ASAP7_75t_L g5163 ( 
.A1(n_5129),
.A2(n_579),
.B(n_580),
.C(n_581),
.Y(n_5163)
);

OAI211xp5_ASAP7_75t_L g5164 ( 
.A1(n_5117),
.A2(n_581),
.B(n_582),
.C(n_583),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5138),
.B(n_583),
.Y(n_5165)
);

O2A1O1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_5124),
.A2(n_585),
.B(n_586),
.C(n_587),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_5148),
.B(n_5120),
.Y(n_5167)
);

OAI211xp5_ASAP7_75t_SL g5168 ( 
.A1(n_5160),
.A2(n_5123),
.B(n_5141),
.C(n_5131),
.Y(n_5168)
);

NOR3x1_ASAP7_75t_L g5169 ( 
.A(n_5164),
.B(n_5165),
.C(n_5162),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_SL g5170 ( 
.A(n_5154),
.B(n_5140),
.Y(n_5170)
);

NAND3xp33_ASAP7_75t_L g5171 ( 
.A(n_5150),
.B(n_5161),
.C(n_5163),
.Y(n_5171)
);

O2A1O1Ixp33_ASAP7_75t_L g5172 ( 
.A1(n_5166),
.A2(n_5119),
.B(n_5122),
.C(n_588),
.Y(n_5172)
);

AOI221xp5_ASAP7_75t_L g5173 ( 
.A1(n_5152),
.A2(n_585),
.B1(n_586),
.B2(n_588),
.C(n_589),
.Y(n_5173)
);

NOR3xp33_ASAP7_75t_L g5174 ( 
.A(n_5156),
.B(n_5151),
.C(n_5158),
.Y(n_5174)
);

NOR4xp75_ASAP7_75t_L g5175 ( 
.A(n_5153),
.B(n_589),
.C(n_590),
.D(n_591),
.Y(n_5175)
);

NOR3xp33_ASAP7_75t_SL g5176 ( 
.A(n_5157),
.B(n_591),
.C(n_592),
.Y(n_5176)
);

NOR2x1_ASAP7_75t_L g5177 ( 
.A(n_5159),
.B(n_5146),
.Y(n_5177)
);

NOR2x1_ASAP7_75t_L g5178 ( 
.A(n_5145),
.B(n_593),
.Y(n_5178)
);

NOR3x1_ASAP7_75t_L g5179 ( 
.A(n_5147),
.B(n_593),
.C(n_594),
.Y(n_5179)
);

NAND4xp25_ASAP7_75t_L g5180 ( 
.A(n_5155),
.B(n_594),
.C(n_595),
.D(n_597),
.Y(n_5180)
);

INVxp67_ASAP7_75t_SL g5181 ( 
.A(n_5149),
.Y(n_5181)
);

AOI21xp5_ASAP7_75t_L g5182 ( 
.A1(n_5158),
.A2(n_597),
.B(n_598),
.Y(n_5182)
);

NAND5xp2_ASAP7_75t_L g5183 ( 
.A(n_5172),
.B(n_599),
.C(n_600),
.D(n_601),
.E(n_602),
.Y(n_5183)
);

OAI21xp5_ASAP7_75t_SL g5184 ( 
.A1(n_5168),
.A2(n_602),
.B(n_603),
.Y(n_5184)
);

AND4x1_ASAP7_75t_L g5185 ( 
.A(n_5174),
.B(n_603),
.C(n_604),
.D(n_605),
.Y(n_5185)
);

NOR3xp33_ASAP7_75t_L g5186 ( 
.A(n_5170),
.B(n_604),
.C(n_605),
.Y(n_5186)
);

NAND4xp25_ASAP7_75t_L g5187 ( 
.A(n_5169),
.B(n_606),
.C(n_607),
.D(n_608),
.Y(n_5187)
);

OAI211xp5_ASAP7_75t_SL g5188 ( 
.A1(n_5176),
.A2(n_607),
.B(n_610),
.C(n_611),
.Y(n_5188)
);

AOI22xp5_ASAP7_75t_L g5189 ( 
.A1(n_5181),
.A2(n_5180),
.B1(n_5171),
.B2(n_5173),
.Y(n_5189)
);

NOR3x1_ASAP7_75t_L g5190 ( 
.A(n_5167),
.B(n_612),
.C(n_613),
.Y(n_5190)
);

NAND4xp25_ASAP7_75t_SL g5191 ( 
.A(n_5182),
.B(n_612),
.C(n_614),
.D(n_615),
.Y(n_5191)
);

NOR3xp33_ASAP7_75t_L g5192 ( 
.A(n_5177),
.B(n_614),
.C(n_617),
.Y(n_5192)
);

NAND4xp25_ASAP7_75t_L g5193 ( 
.A(n_5179),
.B(n_617),
.C(n_618),
.D(n_619),
.Y(n_5193)
);

NOR2xp33_ASAP7_75t_L g5194 ( 
.A(n_5178),
.B(n_618),
.Y(n_5194)
);

AOI221xp5_ASAP7_75t_L g5195 ( 
.A1(n_5175),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.C(n_622),
.Y(n_5195)
);

NOR2xp33_ASAP7_75t_L g5196 ( 
.A(n_5180),
.B(n_622),
.Y(n_5196)
);

NOR2xp67_ASAP7_75t_L g5197 ( 
.A(n_5180),
.B(n_623),
.Y(n_5197)
);

NOR4xp75_ASAP7_75t_L g5198 ( 
.A(n_5170),
.B(n_623),
.C(n_624),
.D(n_625),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_5180),
.B(n_624),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5179),
.B(n_625),
.Y(n_5200)
);

NAND4xp25_ASAP7_75t_SL g5201 ( 
.A(n_5173),
.B(n_626),
.C(n_627),
.D(n_629),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_5190),
.B(n_626),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5200),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5198),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_5185),
.B(n_627),
.Y(n_5205)
);

INVxp67_ASAP7_75t_L g5206 ( 
.A(n_5183),
.Y(n_5206)
);

AOI22xp5_ASAP7_75t_L g5207 ( 
.A1(n_5184),
.A2(n_630),
.B1(n_631),
.B2(n_632),
.Y(n_5207)
);

AOI22xp5_ASAP7_75t_L g5208 ( 
.A1(n_5186),
.A2(n_630),
.B1(n_633),
.B2(n_634),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_5197),
.B(n_633),
.Y(n_5209)
);

OAI22xp5_ASAP7_75t_L g5210 ( 
.A1(n_5189),
.A2(n_5199),
.B1(n_5196),
.B2(n_5195),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5194),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5193),
.Y(n_5212)
);

NOR2x1_ASAP7_75t_L g5213 ( 
.A(n_5187),
.B(n_635),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5188),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_5191),
.Y(n_5215)
);

OAI211xp5_ASAP7_75t_SL g5216 ( 
.A1(n_5192),
.A2(n_636),
.B(n_637),
.C(n_638),
.Y(n_5216)
);

AND2x4_ASAP7_75t_L g5217 ( 
.A(n_5201),
.B(n_636),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5200),
.Y(n_5218)
);

INVx2_ASAP7_75t_L g5219 ( 
.A(n_5190),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_5207),
.B(n_638),
.Y(n_5220)
);

NAND4xp25_ASAP7_75t_L g5221 ( 
.A(n_5213),
.B(n_639),
.C(n_640),
.D(n_641),
.Y(n_5221)
);

NOR2x1_ASAP7_75t_L g5222 ( 
.A(n_5219),
.B(n_639),
.Y(n_5222)
);

INVx1_ASAP7_75t_SL g5223 ( 
.A(n_5202),
.Y(n_5223)
);

NAND4xp25_ASAP7_75t_L g5224 ( 
.A(n_5205),
.B(n_641),
.C(n_642),
.D(n_643),
.Y(n_5224)
);

NAND3xp33_ASAP7_75t_SL g5225 ( 
.A(n_5209),
.B(n_642),
.C(n_643),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5217),
.Y(n_5226)
);

OR2x2_ASAP7_75t_L g5227 ( 
.A(n_5204),
.B(n_644),
.Y(n_5227)
);

NAND3xp33_ASAP7_75t_SL g5228 ( 
.A(n_5208),
.B(n_645),
.C(n_646),
.Y(n_5228)
);

NAND3xp33_ASAP7_75t_SL g5229 ( 
.A(n_5215),
.B(n_645),
.C(n_647),
.Y(n_5229)
);

NAND4xp75_ASAP7_75t_L g5230 ( 
.A(n_5212),
.B(n_648),
.C(n_649),
.D(n_650),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5216),
.Y(n_5231)
);

NAND4xp25_ASAP7_75t_L g5232 ( 
.A(n_5227),
.B(n_5214),
.C(n_5206),
.D(n_5210),
.Y(n_5232)
);

NAND2x1_ASAP7_75t_L g5233 ( 
.A(n_5222),
.B(n_5211),
.Y(n_5233)
);

AND2x4_ASAP7_75t_L g5234 ( 
.A(n_5226),
.B(n_5218),
.Y(n_5234)
);

NOR3xp33_ASAP7_75t_L g5235 ( 
.A(n_5223),
.B(n_5203),
.C(n_5225),
.Y(n_5235)
);

AND2x4_ASAP7_75t_L g5236 ( 
.A(n_5231),
.B(n_650),
.Y(n_5236)
);

NOR2xp67_ASAP7_75t_L g5237 ( 
.A(n_5221),
.B(n_5229),
.Y(n_5237)
);

XNOR2x1_ASAP7_75t_L g5238 ( 
.A(n_5230),
.B(n_651),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5236),
.Y(n_5239)
);

NOR3xp33_ASAP7_75t_SL g5240 ( 
.A(n_5232),
.B(n_5228),
.C(n_5220),
.Y(n_5240)
);

NOR2xp67_ASAP7_75t_L g5241 ( 
.A(n_5237),
.B(n_5224),
.Y(n_5241)
);

AND2x4_ASAP7_75t_L g5242 ( 
.A(n_5235),
.B(n_651),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5242),
.Y(n_5243)
);

HB1xp67_ASAP7_75t_L g5244 ( 
.A(n_5241),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5244),
.Y(n_5245)
);

HB1xp67_ASAP7_75t_L g5246 ( 
.A(n_5245),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_5246),
.B(n_5238),
.Y(n_5247)
);

OAI211xp5_ASAP7_75t_L g5248 ( 
.A1(n_5247),
.A2(n_5233),
.B(n_5240),
.C(n_5239),
.Y(n_5248)
);

AOI221xp5_ASAP7_75t_L g5249 ( 
.A1(n_5248),
.A2(n_5234),
.B1(n_5243),
.B2(n_655),
.C(n_656),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5249),
.Y(n_5250)
);

OA22x2_ASAP7_75t_L g5251 ( 
.A1(n_5250),
.A2(n_653),
.B1(n_654),
.B2(n_656),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5251),
.Y(n_5252)
);

NAND2x1_ASAP7_75t_L g5253 ( 
.A(n_5252),
.B(n_653),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5253),
.Y(n_5254)
);

NAND2xp33_ASAP7_75t_L g5255 ( 
.A(n_5254),
.B(n_657),
.Y(n_5255)
);

OR2x6_ASAP7_75t_L g5256 ( 
.A(n_5254),
.B(n_658),
.Y(n_5256)
);

OAI221xp5_ASAP7_75t_R g5257 ( 
.A1(n_5255),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.C(n_661),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_5257),
.A2(n_5256),
.B1(n_660),
.B2(n_661),
.Y(n_5258)
);

AOI211xp5_ASAP7_75t_L g5259 ( 
.A1(n_5258),
.A2(n_659),
.B(n_662),
.C(n_663),
.Y(n_5259)
);


endmodule