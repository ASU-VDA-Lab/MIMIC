module fake_jpeg_20880_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_38),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_20),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_55),
.B1(n_36),
.B2(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_20),
.B1(n_15),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_25),
.B1(n_17),
.B2(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_18),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_38),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_76),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_78),
.C(n_74),
.Y(n_101)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_74),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_79),
.B1(n_55),
.B2(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_37),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_57),
.C(n_47),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_47),
.B1(n_54),
.B2(n_42),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_84),
.B1(n_98),
.B2(n_60),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_54),
.B1(n_43),
.B2(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_95),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_46),
.B1(n_43),
.B2(n_40),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_61),
.B1(n_77),
.B2(n_62),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_60),
.C(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_108),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_66),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_127),
.B(n_106),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_103),
.B1(n_86),
.B2(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_65),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_79),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_43),
.B1(n_67),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_126),
.B1(n_39),
.B2(n_44),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_76),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_89),
.B1(n_84),
.B2(n_96),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_89),
.B1(n_98),
.B2(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_134),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_113),
.B(n_121),
.C(n_110),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_103),
.B(n_104),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_148),
.B(n_25),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_19),
.B(n_27),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_112),
.B(n_118),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_122),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_114),
.B(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_168),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_99),
.C(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.C(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_99),
.C(n_34),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_148),
.B1(n_22),
.B2(n_23),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_26),
.C(n_30),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_25),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_134),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_179),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_143),
.B1(n_149),
.B2(n_150),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_177),
.B1(n_187),
.B2(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_152),
.B1(n_144),
.B2(n_130),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_133),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_183),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

AOI321xp33_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_145),
.A3(n_141),
.B1(n_147),
.B2(n_132),
.C(n_28),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_16),
.B(n_1),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_132),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_22),
.C(n_16),
.Y(n_198)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_154),
.B1(n_171),
.B2(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_36),
.B1(n_30),
.B2(n_23),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_170),
.B1(n_163),
.B2(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_194),
.B1(n_197),
.B2(n_0),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_174),
.B(n_179),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_0),
.B(n_2),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_166),
.B1(n_165),
.B2(n_169),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_185),
.C(n_173),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_207),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_13),
.C(n_12),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_190),
.C(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_209),
.B1(n_193),
.B2(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_12),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_206),
.A2(n_189),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_203),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_0),
.B(n_3),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_3),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_221),
.B(n_222),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_201),
.B(n_5),
.C(n_7),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_216),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_7),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_213),
.B(n_5),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_4),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.C(n_7),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_231),
.B(n_9),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_9),
.C(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_10),
.Y(n_233)
);


endmodule