module real_aes_6313_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g264 ( .A(n_0), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_1), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_2), .A2(n_43), .B1(n_153), .B2(n_157), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_3), .A2(n_30), .B1(n_219), .B2(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_4), .B(n_244), .Y(n_253) );
INVx1_ASAP7_75t_L g200 ( .A(n_5), .Y(n_200) );
AND2x6_ASAP7_75t_L g237 ( .A(n_5), .B(n_198), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_5), .B(n_518), .Y(n_517) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_6), .A2(n_25), .B1(n_92), .B2(n_97), .Y(n_101) );
INVx1_ASAP7_75t_L g215 ( .A(n_7), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_8), .A2(n_76), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_8), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_8), .B(n_223), .Y(n_292) );
INVx1_ASAP7_75t_L g257 ( .A(n_9), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_10), .B(n_211), .Y(n_328) );
AO32x2_ASAP7_75t_L g270 ( .A1(n_11), .A2(n_210), .A3(n_236), .B1(n_244), .B2(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_12), .B(n_219), .Y(n_296) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_13), .A2(n_27), .B1(n_92), .B2(n_93), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_14), .B(n_211), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_15), .A2(n_40), .B1(n_219), .B2(n_273), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g312 ( .A1(n_16), .A2(n_61), .B1(n_219), .B2(n_223), .Y(n_312) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_16), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_17), .B(n_219), .Y(n_285) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_18), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_19), .B(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_20), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_21), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_22), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_23), .B(n_239), .Y(n_287) );
INVx2_ASAP7_75t_L g221 ( .A(n_24), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_26), .B(n_219), .Y(n_218) );
OAI221xp5_ASAP7_75t_L g191 ( .A1(n_27), .A2(n_46), .B1(n_56), .B2(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_27), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_28), .B(n_239), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_29), .A2(n_81), .B1(n_171), .B2(n_172), .Y(n_80) );
INVxp67_ASAP7_75t_L g171 ( .A(n_29), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_31), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_32), .A2(n_58), .B1(n_135), .B2(n_138), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_33), .B(n_219), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_34), .A2(n_57), .B1(n_123), .B2(n_130), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_35), .A2(n_69), .B1(n_273), .B2(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_36), .B(n_219), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_37), .B(n_219), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_38), .A2(n_81), .B1(n_172), .B2(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_38), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_39), .B(n_231), .Y(n_251) );
AOI222xp33_ASAP7_75t_L g161 ( .A1(n_41), .A2(n_47), .B1(n_60), .B2(n_162), .C1(n_163), .C2(n_167), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_42), .A2(n_48), .B1(n_219), .B2(n_223), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_44), .B(n_219), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_45), .B(n_219), .Y(n_291) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_46), .A2(n_65), .B1(n_92), .B2(n_93), .Y(n_91) );
INVxp67_ASAP7_75t_L g195 ( .A(n_46), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_49), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_50), .B(n_219), .Y(n_265) );
INVx1_ASAP7_75t_L g214 ( .A(n_51), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_52), .Y(n_192) );
AO32x2_ASAP7_75t_L g308 ( .A1(n_53), .A2(n_236), .A3(n_244), .B1(n_309), .B2(n_313), .Y(n_308) );
INVx1_ASAP7_75t_L g229 ( .A(n_54), .Y(n_229) );
INVx1_ASAP7_75t_L g282 ( .A(n_55), .Y(n_282) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_56), .A2(n_73), .B1(n_92), .B2(n_97), .Y(n_96) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_59), .B(n_223), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_62), .A2(n_74), .B1(n_177), .B2(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g178 ( .A(n_62), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_63), .B(n_273), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_64), .B(n_223), .Y(n_286) );
INVx2_ASAP7_75t_L g212 ( .A(n_66), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_67), .B(n_223), .Y(n_248) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_68), .A2(n_181), .B1(n_182), .B2(n_185), .Y(n_180) );
CKINVDCx14_ASAP7_75t_R g185 ( .A(n_68), .Y(n_185) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_69), .A2(n_81), .B1(n_172), .B2(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_69), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_70), .A2(n_77), .B1(n_223), .B2(n_224), .Y(n_325) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_71), .A2(n_174), .B1(n_175), .B2(n_187), .Y(n_173) );
INVx1_ASAP7_75t_L g187 ( .A(n_71), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g177 ( .A(n_74), .Y(n_177) );
INVx1_ASAP7_75t_L g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
INVx1_ASAP7_75t_L g184 ( .A(n_76), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_76), .B(n_223), .Y(n_222) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_188), .B1(n_201), .B2(n_506), .C(n_512), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_173), .Y(n_79) );
INVx2_ASAP7_75t_SL g172 ( .A(n_81), .Y(n_172) );
AND4x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_121), .C(n_141), .D(n_161), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_110), .Y(n_82) );
OAI22xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_85), .B1(n_102), .B2(n_103), .Y(n_83) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx6_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_98), .Y(n_88) );
AND2x2_ASAP7_75t_L g115 ( .A(n_89), .B(n_108), .Y(n_115) );
AND2x6_ASAP7_75t_L g127 ( .A(n_89), .B(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_L g162 ( .A(n_89), .B(n_160), .Y(n_162) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g120 ( .A(n_90), .B(n_96), .Y(n_120) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g106 ( .A(n_91), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_91), .B(n_96), .Y(n_133) );
AND2x2_ASAP7_75t_L g156 ( .A(n_91), .B(n_101), .Y(n_156) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g97 ( .A(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g107 ( .A(n_96), .Y(n_107) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
AND2x2_ASAP7_75t_L g137 ( .A(n_98), .B(n_106), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_98), .B(n_120), .Y(n_150) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_100), .Y(n_98) );
INVx2_ASAP7_75t_L g109 ( .A(n_99), .Y(n_109) );
OR2x2_ASAP7_75t_L g129 ( .A(n_99), .B(n_100), .Y(n_129) );
INVx1_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
AND2x2_ASAP7_75t_L g160 ( .A(n_99), .B(n_101), .Y(n_160) );
AND2x2_ASAP7_75t_L g108 ( .A(n_100), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
AND2x4_ASAP7_75t_L g119 ( .A(n_108), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g131 ( .A(n_108), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g165 ( .A(n_109), .B(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B1(n_116), .B2(n_117), .Y(n_110) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_134), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx11_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g144 ( .A(n_129), .B(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x6_ASAP7_75t_L g139 ( .A(n_133), .B(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx8_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx6_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI221xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_146), .B1(n_147), .B2(n_151), .C(n_152), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x4_ASAP7_75t_L g164 ( .A(n_156), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g169 ( .A(n_156), .B(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_166), .Y(n_170) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B1(n_180), .B2(n_186), .Y(n_175) );
INVx1_ASAP7_75t_L g186 ( .A(n_176), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
AND3x1_ASAP7_75t_SL g190 ( .A(n_191), .B(n_196), .C(n_199), .Y(n_190) );
INVxp67_ASAP7_75t_L g518 ( .A(n_191), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_SL g519 ( .A(n_196), .Y(n_519) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_196), .A2(n_511), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g529 ( .A(n_196), .Y(n_529) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_197), .B(n_200), .Y(n_521) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_SL g528 ( .A(n_199), .B(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR3x1_ASAP7_75t_L g203 ( .A(n_204), .B(n_434), .C(n_483), .Y(n_203) );
NAND5xp2_ASAP7_75t_L g204 ( .A(n_205), .B(n_349), .C(n_377), .D(n_407), .E(n_421), .Y(n_204) );
AOI221xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_267), .B1(n_299), .B2(n_304), .C(n_315), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_240), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_207), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g329 ( .A(n_208), .Y(n_329) );
AND2x2_ASAP7_75t_L g337 ( .A(n_208), .B(n_243), .Y(n_337) );
AND2x2_ASAP7_75t_L g360 ( .A(n_208), .B(n_242), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_208), .B(n_254), .Y(n_375) );
OR2x2_ASAP7_75t_L g384 ( .A(n_208), .B(n_322), .Y(n_384) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_208), .Y(n_387) );
AND2x2_ASAP7_75t_L g495 ( .A(n_208), .B(n_322), .Y(n_495) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_216), .B(n_238), .Y(n_208) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_209), .A2(n_255), .B(n_266), .Y(n_254) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_212), .B(n_213), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_228), .B(n_236), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_222), .B(n_225), .Y(n_217) );
INVx3_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
BUFx3_ASAP7_75t_L g311 ( .A(n_220), .Y(n_311) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g224 ( .A(n_221), .Y(n_224) );
INVx1_ASAP7_75t_L g232 ( .A(n_221), .Y(n_232) );
INVx2_ASAP7_75t_L g258 ( .A(n_223), .Y(n_258) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_225), .A2(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_SL g280 ( .A1(n_225), .A2(n_281), .B(n_282), .C(n_283), .Y(n_280) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g309 ( .A1(n_226), .A2(n_235), .B1(n_310), .B2(n_312), .Y(n_309) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
INVx1_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
AND2x2_ASAP7_75t_L g511 ( .A(n_227), .B(n_232), .Y(n_511) );
O2A1O1Ixp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_233), .C(n_234), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_230), .A2(n_252), .B(n_264), .C(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_234), .A2(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_235), .A2(n_252), .B1(n_272), .B2(n_274), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_235), .A2(n_252), .B1(n_325), .B2(n_326), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_236), .B(n_323), .C(n_324), .Y(n_348) );
BUFx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_237), .A2(n_246), .B(n_249), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_237), .A2(n_256), .B(n_263), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_237), .A2(n_280), .B(n_284), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_237), .A2(n_290), .B(n_295), .Y(n_289) );
AND2x4_ASAP7_75t_L g510 ( .A(n_237), .B(n_511), .Y(n_510) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_239), .A2(n_279), .B(n_287), .Y(n_278) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_239), .A2(n_289), .B(n_298), .Y(n_288) );
INVx2_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_240), .B(n_387), .Y(n_443) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OAI311xp33_ASAP7_75t_L g385 ( .A1(n_241), .A2(n_386), .A3(n_387), .B1(n_388), .C1(n_403), .Y(n_385) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_254), .Y(n_241) );
AND2x2_ASAP7_75t_L g346 ( .A(n_242), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g353 ( .A(n_242), .Y(n_353) );
AND2x2_ASAP7_75t_L g474 ( .A(n_242), .B(n_303), .Y(n_474) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_243), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g330 ( .A(n_243), .B(n_254), .Y(n_330) );
AND2x2_ASAP7_75t_L g382 ( .A(n_243), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g396 ( .A(n_243), .B(n_329), .Y(n_396) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_253), .Y(n_243) );
INVx4_ASAP7_75t_L g323 ( .A(n_244), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_252), .Y(n_249) );
INVx2_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
AND2x2_ASAP7_75t_L g345 ( .A(n_254), .B(n_329), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_259), .C(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_285), .B(n_286), .Y(n_284) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_275), .Y(n_267) );
OR2x2_ASAP7_75t_L g440 ( .A(n_268), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_268), .B(n_446), .Y(n_457) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_269), .B(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g314 ( .A(n_270), .Y(n_314) );
AND2x2_ASAP7_75t_L g381 ( .A(n_270), .B(n_308), .Y(n_381) );
AND2x2_ASAP7_75t_L g392 ( .A(n_270), .B(n_288), .Y(n_392) );
AND2x2_ASAP7_75t_L g401 ( .A(n_270), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_275), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_275), .B(n_342), .Y(n_386) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g373 ( .A(n_276), .B(n_332), .Y(n_373) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_288), .Y(n_276) );
INVx2_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
AND2x2_ASAP7_75t_L g400 ( .A(n_277), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
OR2x2_ASAP7_75t_L g417 ( .A(n_278), .B(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_278), .Y(n_480) );
AND2x2_ASAP7_75t_L g319 ( .A(n_288), .B(n_314), .Y(n_319) );
INVx1_ASAP7_75t_L g340 ( .A(n_288), .Y(n_340) );
AND2x2_ASAP7_75t_L g361 ( .A(n_288), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g402 ( .A(n_288), .Y(n_402) );
INVx1_ASAP7_75t_L g418 ( .A(n_288), .Y(n_418) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_288), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_301), .B(n_406), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_301), .A2(n_391), .B1(n_440), .B2(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI211xp5_ASAP7_75t_SL g483 ( .A1(n_302), .A2(n_484), .B(n_486), .C(n_504), .Y(n_483) );
INVx2_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
AND2x2_ASAP7_75t_L g394 ( .A(n_303), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g405 ( .A(n_303), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_304), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AND2x2_ASAP7_75t_L g378 ( .A(n_305), .B(n_342), .Y(n_378) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g410 ( .A(n_306), .B(n_401), .Y(n_410) );
AND2x2_ASAP7_75t_L g429 ( .A(n_306), .B(n_343), .Y(n_429) );
AND2x4_ASAP7_75t_L g365 ( .A(n_307), .B(n_339), .Y(n_365) );
AND2x2_ASAP7_75t_L g503 ( .A(n_307), .B(n_479), .Y(n_503) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_314), .Y(n_307) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx1_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
INVx1_ASAP7_75t_L g442 ( .A(n_308), .Y(n_442) );
OR2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_318), .Y(n_333) );
AND2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_343), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_314), .B(n_363), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B1(n_331), .B2(n_334), .C(n_338), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_317), .A2(n_339), .B(n_341), .C(n_344), .Y(n_338) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_318), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_318), .B(n_340), .Y(n_446) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_318), .Y(n_453) );
AND2x2_ASAP7_75t_L g371 ( .A(n_319), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g408 ( .A(n_319), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_330), .Y(n_320) );
INVx2_ASAP7_75t_L g399 ( .A(n_321), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_321), .A2(n_332), .B1(n_449), .B2(n_451), .C1(n_452), .C2(n_454), .Y(n_448) );
AND2x2_ASAP7_75t_L g505 ( .A(n_321), .B(n_474), .Y(n_505) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_329), .Y(n_321) );
INVx1_ASAP7_75t_L g395 ( .A(n_322), .Y(n_395) );
AO21x1_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g347 ( .A(n_328), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g433 ( .A(n_330), .B(n_367), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_331), .A2(n_445), .B(n_447), .Y(n_444) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_339), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_332), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx3_ASAP7_75t_L g398 ( .A(n_336), .Y(n_398) );
OR2x2_ASAP7_75t_L g450 ( .A(n_336), .B(n_372), .Y(n_450) );
AND2x2_ASAP7_75t_L g366 ( .A(n_337), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_337), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_337), .B(n_398), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_337), .B(n_394), .Y(n_420) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_406), .Y(n_424) );
INVxp67_ASAP7_75t_L g356 ( .A(n_339), .Y(n_356) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_341), .A2(n_414), .B1(n_419), .B2(n_420), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_341), .B(n_446), .Y(n_476) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g462 ( .A(n_342), .B(n_453), .Y(n_462) );
AND2x2_ASAP7_75t_L g491 ( .A(n_342), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g496 ( .A(n_342), .B(n_446), .Y(n_496) );
INVx1_ASAP7_75t_L g409 ( .A(n_343), .Y(n_409) );
BUFx2_ASAP7_75t_L g415 ( .A(n_343), .Y(n_415) );
INVx1_ASAP7_75t_L g500 ( .A(n_344), .Y(n_500) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_345), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
NOR2x1_ASAP7_75t_L g352 ( .A(n_347), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_347), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
INVx3_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
OR2x2_ASAP7_75t_L g472 ( .A(n_347), .B(n_473), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B(n_357), .C(n_369), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_350), .A2(n_487), .B1(n_494), .B2(n_496), .C(n_497), .Y(n_486) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_358), .B(n_364), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_360), .B(n_398), .Y(n_412) );
AND2x2_ASAP7_75t_L g454 ( .A(n_360), .B(n_394), .Y(n_454) );
INVx1_ASAP7_75t_SL g467 ( .A(n_361), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_361), .B(n_415), .Y(n_470) );
INVx1_ASAP7_75t_L g488 ( .A(n_362), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_366), .A2(n_456), .B1(n_458), .B2(n_462), .C(n_463), .Y(n_455) );
AND2x2_ASAP7_75t_L g482 ( .A(n_367), .B(n_474), .Y(n_482) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g466 ( .A(n_368), .Y(n_466) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_373), .B(n_374), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g437 ( .A(n_372), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
INVx1_ASAP7_75t_L g451 ( .A(n_374), .Y(n_451) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_382), .C(n_385), .Y(n_377) );
OAI31xp33_ASAP7_75t_L g504 ( .A1(n_378), .A2(n_416), .A3(n_503), .B(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g478 ( .A(n_381), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g499 ( .A(n_381), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_383), .B(n_398), .Y(n_426) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g501 ( .A(n_384), .B(n_398), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B1(n_397), .B2(n_400), .Y(n_388) );
NAND2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_392), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g428 ( .A(n_392), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_392), .B(n_415), .Y(n_431) );
AND2x2_ASAP7_75t_L g485 ( .A(n_392), .B(n_480), .Y(n_485) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
OAI32xp33_ASAP7_75t_L g463 ( .A1(n_398), .A2(n_432), .A3(n_464), .B1(n_466), .B2(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_401), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_411), .C(n_413), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_409), .B(n_446), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_410), .A2(n_422), .B1(n_423), .B2(n_424), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_420), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_430), .B2(n_432), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND4xp25_ASAP7_75t_SL g487 ( .A(n_430), .B(n_488), .C(n_489), .D(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
NAND4xp25_ASAP7_75t_SL g434 ( .A(n_435), .B(n_448), .C(n_455), .D(n_468), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_443), .C(n_444), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g465 ( .A(n_441), .Y(n_465) );
INVx2_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
OR2x2_ASAP7_75t_L g498 ( .A(n_453), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_475), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g494 ( .A(n_474), .B(n_495), .Y(n_494) );
AOI21xp33_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B(n_481), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_497) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI322xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_515), .A3(n_519), .B1(n_520), .B2(n_522), .C1(n_524), .C2(n_526), .Y(n_512) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
endmodule