module fake_aes_6088_n_22 (n_1, n_2, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
NAND2xp5_ASAP7_75t_SL g6 ( .A(n_2), .B(n_3), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVxp67_ASAP7_75t_SL g8 ( .A(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g9 ( .A(n_3), .B(n_2), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_0), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_13), .B(n_10), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_11), .B(n_7), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_11), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
OAI21xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_12), .B(n_15), .Y(n_18) );
OAI22xp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_7), .B1(n_9), .B2(n_3), .Y(n_19) );
OAI21xp5_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_1), .B(n_2), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AOI222xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_4), .B1(n_5), .B2(n_19), .C1(n_20), .C2(n_18), .Y(n_22) );
endmodule