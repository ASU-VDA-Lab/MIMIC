module fake_jpeg_4297_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_10),
.B(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_44),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_53),
.B1(n_69),
.B2(n_21),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_63),
.B1(n_43),
.B2(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_32),
.C(n_23),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_17),
.C(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_44),
.B1(n_19),
.B2(n_18),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_76),
.B1(n_82),
.B2(n_63),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_42),
.B1(n_37),
.B2(n_19),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_44),
.B1(n_19),
.B2(n_32),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_41),
.C(n_40),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_93),
.C(n_19),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_56),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_41),
.C(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_60),
.A3(n_46),
.B1(n_40),
.B2(n_41),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_87),
.B(n_74),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_106),
.Y(n_120)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_107),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_108),
.B1(n_115),
.B2(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_58),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_49),
.B1(n_47),
.B2(n_62),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_49),
.B1(n_62),
.B2(n_48),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_48),
.B(n_47),
.C(n_41),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_35),
.B1(n_18),
.B2(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_78),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_72),
.B1(n_85),
.B2(n_78),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_143),
.B(n_115),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_124),
.B(n_141),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_131),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_145),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_74),
.B(n_89),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_90),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_77),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_137),
.B(n_91),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_117),
.C(n_101),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_158),
.C(n_123),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_101),
.C(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_164),
.B1(n_136),
.B2(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_115),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_168),
.B(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_102),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_114),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_166),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_133),
.B1(n_165),
.B2(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_176),
.B1(n_160),
.B2(n_164),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_136),
.B1(n_108),
.B2(n_144),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_192),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_184),
.C(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_126),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_126),
.C(n_122),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_86),
.C(n_129),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_143),
.C(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_188),
.C(n_193),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_143),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_81),
.B(n_137),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_195),
.B(n_153),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_89),
.C(n_113),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_121),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_195),
.B(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_153),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_146),
.C(n_149),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_219),
.C(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_121),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_168),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_150),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_151),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_170),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_168),
.C(n_165),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_191),
.B1(n_173),
.B2(n_190),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_235),
.B1(n_25),
.B2(n_22),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_0),
.B(n_1),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_173),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_237),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_219),
.A2(n_194),
.B1(n_183),
.B2(n_172),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_239),
.B1(n_228),
.B2(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_198),
.C(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_215),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_171),
.B1(n_154),
.B2(n_150),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_156),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_171),
.B1(n_154),
.B2(n_88),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_249),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_218),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_246),
.B(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_248),
.C(n_225),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_203),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_223),
.B(n_230),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_198),
.C(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_205),
.B1(n_201),
.B2(n_25),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_252),
.B1(n_16),
.B2(n_22),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_10),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_22),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_224),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_258),
.C(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_261),
.B(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_223),
.C(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_248),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_234),
.C(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

OAI322xp33_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_65),
.A3(n_52),
.B1(n_16),
.B2(n_9),
.C1(n_4),
.C2(n_5),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_7),
.B(n_15),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_240),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_5),
.C(n_14),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_265),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_4),
.C2(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_273),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_287),
.B(n_274),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_9),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_270),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_12),
.B(n_1),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_290),
.B(n_280),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_276),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_292),
.B(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_274),
.Y(n_293)
);

NOR3x1_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_0),
.C(n_2),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_287),
.B(n_282),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_297),
.A2(n_298),
.B(n_294),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_300),
.A3(n_296),
.B1(n_3),
.B2(n_2),
.C1(n_65),
.C2(n_52),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_3),
.C(n_294),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_3),
.Y(n_303)
);


endmodule