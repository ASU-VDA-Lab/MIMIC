module fake_jpeg_21902_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_24),
.B1(n_17),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_60),
.B1(n_17),
.B2(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_57),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_24),
.B1(n_17),
.B2(n_27),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_24),
.B1(n_17),
.B2(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_64),
.B1(n_89),
.B2(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_80),
.B1(n_16),
.B2(n_31),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_29),
.B1(n_19),
.B2(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_33),
.B(n_28),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_49),
.CI(n_56),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_107),
.B1(n_79),
.B2(n_19),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_58),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_54),
.B1(n_64),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_112),
.B1(n_23),
.B2(n_26),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_62),
.A3(n_63),
.B1(n_36),
.B2(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_92),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_86),
.C(n_73),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_98),
.CI(n_112),
.CON(n_140),
.SN(n_140)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_73),
.B(n_79),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_134),
.B(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_132),
.B1(n_113),
.B2(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_94),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_128),
.B1(n_129),
.B2(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_44),
.B1(n_41),
.B2(n_31),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_44),
.B1(n_31),
.B2(n_23),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_105),
.B1(n_85),
.B2(n_77),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_30),
.B1(n_16),
.B2(n_32),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_30),
.B(n_20),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_104),
.B(n_115),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_84),
.B(n_18),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_33),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_42),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_155),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_163),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_113),
.B(n_42),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_95),
.B1(n_111),
.B2(n_90),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_161),
.B1(n_128),
.B2(n_129),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_117),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_33),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_97),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_97),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_130),
.C(n_126),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_173),
.C(n_185),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_184),
.Y(n_201)
);

OAI22x1_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_133),
.B1(n_137),
.B2(n_132),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_183),
.B1(n_161),
.B2(n_145),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_153),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_186),
.B(n_153),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_81),
.B1(n_97),
.B2(n_0),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_28),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_28),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_157),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_191),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_146),
.C(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_199),
.C(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_196),
.B(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_205),
.B1(n_169),
.B2(n_167),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_143),
.C(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_155),
.B1(n_140),
.B2(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_149),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_164),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_183),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_175),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_177),
.B1(n_175),
.B2(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_186),
.C(n_181),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_15),
.B(n_4),
.Y(n_239)
);

OAI22x1_ASAP7_75t_SL g218 ( 
.A1(n_208),
.A2(n_172),
.B1(n_140),
.B2(n_168),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_225),
.B1(n_8),
.B2(n_1),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.C(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_150),
.C(n_28),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_150),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_200),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_226),
.B(n_192),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_207),
.B1(n_209),
.B2(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_237),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_205),
.B1(n_197),
.B2(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_233),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_228),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_198),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_238),
.B1(n_217),
.B2(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_28),
.C(n_0),
.Y(n_237)
);

OA21x2_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_1),
.B(n_3),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_239),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_219),
.B1(n_221),
.B2(n_213),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_248),
.B1(n_230),
.B2(n_236),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_250),
.B(n_6),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_5),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_227),
.C(n_229),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_255),
.B(n_241),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_237),
.B(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_259),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_266),
.C(n_251),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_249),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_6),
.B(n_7),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_11),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_8),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_266),
.C(n_12),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_8),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_11),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_274),
.C(n_11),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_268),
.B(n_12),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.C(n_13),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_13),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_14),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_14),
.Y(n_280)
);


endmodule