module fake_jpeg_31532_n_393 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_21),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_14),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_55),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_67),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_60),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_64),
.Y(n_125)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_81),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_13),
.CON(n_64),
.SN(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_30),
.B1(n_45),
.B2(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_1),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_37),
.Y(n_95)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_35),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_71),
.B1(n_78),
.B2(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_86),
.A2(n_48),
.B1(n_55),
.B2(n_9),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_88),
.B(n_6),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_35),
.B1(n_24),
.B2(n_29),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_100),
.B1(n_107),
.B2(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_61),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_35),
.B1(n_33),
.B2(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_98),
.A2(n_105),
.B1(n_126),
.B2(n_127),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_124),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_35),
.B1(n_24),
.B2(n_29),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_33),
.B1(n_30),
.B2(n_40),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_108),
.B1(n_114),
.B2(n_119),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_33),
.B1(n_45),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_30),
.B1(n_39),
.B2(n_31),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_46),
.B1(n_31),
.B2(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_48),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_46),
.B1(n_39),
.B2(n_42),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_134),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_46),
.B1(n_34),
.B2(n_32),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_27),
.B1(n_22),
.B2(n_4),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_136),
.B1(n_60),
.B2(n_58),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_70),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_48),
.B1(n_62),
.B2(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_55),
.B(n_2),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_53),
.B1(n_72),
.B2(n_66),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_144),
.B1(n_149),
.B2(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_49),
.B1(n_60),
.B2(n_58),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_146),
.A2(n_121),
.B1(n_117),
.B2(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_62),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_92),
.B(n_61),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_160),
.Y(n_188)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_170),
.B(n_87),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_161),
.B1(n_178),
.B2(n_113),
.Y(n_199)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_94),
.B(n_6),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_161)
);

NAND4xp25_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_8),
.C(n_12),
.D(n_13),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_166),
.Y(n_187)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_13),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_169),
.Y(n_194)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_88),
.B(n_125),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_R g171 ( 
.A(n_125),
.B(n_90),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_176),
.B(n_115),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_133),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_135),
.C(n_95),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_106),
.C(n_101),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_115),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_113),
.B1(n_123),
.B2(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_132),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_124),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_196),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_120),
.C(n_101),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_106),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_142),
.B(n_169),
.C(n_159),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_106),
.Y(n_196)
);

CKINVDCx11_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_145),
.B(n_87),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_202),
.B1(n_154),
.B2(n_165),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_214),
.B1(n_151),
.B2(n_162),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_151),
.B1(n_139),
.B2(n_137),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_181),
.B1(n_199),
.B2(n_182),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_120),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_213),
.B(n_156),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_96),
.C(n_116),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_96),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_217),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_159),
.A2(n_116),
.B(n_117),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_172),
.B(n_129),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_218),
.A2(n_225),
.B(n_243),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_169),
.B(n_138),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_220),
.B(n_239),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_147),
.B(n_140),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_226),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_234),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_183),
.A2(n_137),
.B1(n_152),
.B2(n_144),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_240),
.B1(n_246),
.B2(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_235),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_161),
.B1(n_170),
.B2(n_175),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_180),
.A2(n_157),
.B1(n_129),
.B2(n_174),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_181),
.A2(n_123),
.B1(n_166),
.B2(n_158),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_242),
.B1(n_191),
.B2(n_200),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_184),
.A2(n_123),
.B1(n_141),
.B2(n_143),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_158),
.B(n_168),
.C(n_164),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_249),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_192),
.A2(n_209),
.B1(n_200),
.B2(n_184),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_210),
.B(n_215),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_211),
.B(n_196),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_188),
.B(n_192),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_248),
.C(n_228),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_253),
.C(n_261),
.Y(n_284)
);

OAI22x1_ASAP7_75t_L g252 ( 
.A1(n_219),
.A2(n_217),
.B1(n_186),
.B2(n_205),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_231),
.B1(n_237),
.B2(n_221),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_228),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_258),
.B1(n_275),
.B2(n_276),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_186),
.B1(n_194),
.B2(n_212),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_193),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_240),
.B1(n_244),
.B2(n_227),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_194),
.C(n_188),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_269),
.C(n_273),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_271),
.B(n_239),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_216),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_216),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_246),
.A2(n_216),
.B1(n_209),
.B2(n_208),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_225),
.A2(n_216),
.B1(n_209),
.B2(n_208),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_292),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_291),
.B1(n_293),
.B2(n_296),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_224),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_221),
.B(n_241),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_289),
.B(n_295),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_286),
.A2(n_298),
.B1(n_299),
.B2(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_223),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_236),
.B1(n_242),
.B2(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_237),
.B1(n_222),
.B2(n_243),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_237),
.C(n_220),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_261),
.C(n_250),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_251),
.A2(n_243),
.B(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_222),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_267),
.B1(n_252),
.B2(n_257),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_243),
.B1(n_234),
.B2(n_233),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_300),
.B(n_314),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_307),
.B1(n_277),
.B2(n_291),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_254),
.B(n_243),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_279),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_258),
.B1(n_256),
.B2(n_276),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_264),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_316),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_254),
.C(n_273),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_299),
.C(n_298),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_256),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_262),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_294),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_274),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_282),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_243),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_330),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_336),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_309),
.B1(n_322),
.B2(n_332),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_287),
.C(n_281),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_326),
.C(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_285),
.C(n_288),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_285),
.B(n_297),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_328),
.B(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_280),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_295),
.C(n_277),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_334),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_303),
.A2(n_289),
.B(n_295),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_293),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_296),
.C(n_292),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_312),
.C(n_320),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_310),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_314),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_339),
.B(n_343),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_321),
.A2(n_305),
.B1(n_312),
.B2(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_346),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_325),
.B(n_335),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_319),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_344),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_311),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_324),
.C(n_327),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_349),
.B(n_350),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_326),
.B(n_329),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_337),
.C(n_327),
.Y(n_357)
);

INVx11_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_353),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_270),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_357),
.A2(n_352),
.B1(n_348),
.B2(n_345),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_351),
.A2(n_310),
.B1(n_306),
.B2(n_301),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_259),
.B1(n_270),
.B2(n_266),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_361),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_340),
.B(n_324),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_363),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_340),
.B(n_302),
.C(n_259),
.Y(n_363)
);

OAI321xp33_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_279),
.A3(n_306),
.B1(n_346),
.B2(n_271),
.C(n_349),
.Y(n_364)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_279),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_367),
.B(n_370),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_358),
.A2(n_279),
.B(n_344),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_372),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_355),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_363),
.Y(n_378)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_374),
.A2(n_203),
.B1(n_249),
.B2(n_376),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_355),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_375),
.A2(n_266),
.B1(n_235),
.B2(n_238),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_359),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_360),
.C(n_356),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_380),
.B(n_368),
.C(n_357),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_377),
.A2(n_369),
.B(n_370),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_384),
.C(n_385),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_381),
.C(n_375),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_388),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_391),
.C(n_379),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_387),
.A2(n_379),
.B(n_203),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_203),
.Y(n_393)
);


endmodule