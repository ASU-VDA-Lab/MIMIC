module fake_jpeg_470_n_13 (n_0, n_2, n_1, n_13);

input n_0;
input n_2;
input n_1;

output n_13;

wire n_11;
wire n_3;
wire n_10;
wire n_12;
wire n_4;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_L g3 ( 
.A(n_2),
.B(n_1),
.Y(n_3)
);

INVx4_ASAP7_75t_L g4 ( 
.A(n_1),
.Y(n_4)
);

INVx4_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

HB1xp67_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_0),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_7),
.A2(n_8),
.B(n_3),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_3),
.A2(n_0),
.B(n_1),
.Y(n_8)
);

AO221x1_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.C(n_10),
.Y(n_11)
);

AOI31xp67_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_4),
.A3(n_5),
.B(n_9),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_12),
.B(n_5),
.Y(n_13)
);


endmodule