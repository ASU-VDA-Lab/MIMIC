module fake_jpeg_22362_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_25),
.B1(n_13),
.B2(n_20),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_28),
.B1(n_29),
.B2(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_25),
.B1(n_20),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_13),
.B1(n_16),
.B2(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_12),
.B1(n_35),
.B2(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_60),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_51),
.B(n_37),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_34),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_62),
.B1(n_39),
.B2(n_37),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_2),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_3),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_60),
.C(n_50),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_41),
.B(n_47),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_48),
.B(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_51),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_51),
.B(n_58),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_62),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_82),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_48),
.C(n_53),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_65),
.C(n_64),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_78),
.C(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_82),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_71),
.C(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_70),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_94),
.B1(n_72),
.B2(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_88),
.B1(n_85),
.B2(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_72),
.B1(n_90),
.B2(n_73),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_103),
.B(n_10),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

AOI21x1_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_66),
.B(n_7),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_8),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_11),
.B(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule