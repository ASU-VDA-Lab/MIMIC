module real_jpeg_15531_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_434),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_1),
.B(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_2),
.A2(n_54),
.B1(n_130),
.B2(n_151),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_2),
.A2(n_54),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_2),
.A2(n_54),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_3),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_3),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_123),
.B1(n_125),
.B2(n_129),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_6),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_84),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_84),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_92)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_103),
.A3(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_11),
.A2(n_159),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_11),
.B(n_134),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_11),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_11),
.B(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g173 ( 
.A(n_12),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_12),
.Y(n_175)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_212),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_210),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_190),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_SL g211 ( 
.A(n_18),
.B(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.C(n_153),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_19),
.A2(n_135),
.B1(n_136),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_19),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_55),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_20),
.A2(n_192),
.B1(n_193),
.B2(n_207),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_20),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_20),
.B(n_393),
.Y(n_397)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_30),
.B1(n_42),
.B2(n_50),
.Y(n_20)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_21),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_21),
.A2(n_30),
.B1(n_42),
.B2(n_50),
.Y(n_195)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_26),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_26),
.B(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_30),
.B(n_42),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_37),
.B(n_42),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_31),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_39),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g354 ( 
.A(n_41),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_42),
.Y(n_323)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_90),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_56),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_56),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_80),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_139),
.B(n_157),
.Y(n_156)
);

AOI21x1_ASAP7_75t_SL g334 ( 
.A1(n_58),
.A2(n_335),
.B(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_69),
.Y(n_68)
);

AO22x2_ASAP7_75t_L g238 ( 
.A1(n_59),
.A2(n_68),
.B1(n_158),
.B2(n_239),
.Y(n_238)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_59),
.A2(n_68),
.B1(n_158),
.B2(n_239),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_59)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_62),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_63),
.Y(n_369)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_65),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_71),
.Y(n_244)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_138),
.B1(n_147),
.B2(n_148),
.Y(n_137)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_90),
.B(n_207),
.C(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B1(n_122),
.B2(n_134),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_92),
.A2(n_101),
.B1(n_113),
.B2(n_150),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_92),
.A2(n_101),
.B1(n_113),
.B2(n_150),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_92),
.A2(n_101),
.B(n_113),
.Y(n_393)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_97),
.Y(n_350)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_98),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_98),
.B(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_122),
.B1(n_134),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2x1p5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OA22x2_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_118),
.Y(n_271)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_123),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_124),
.A2(n_145),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_125),
.A2(n_342),
.B1(n_351),
.B2(n_355),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_136),
.A2(n_137),
.B(n_149),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_148),
.B(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_149),
.A2(n_319),
.B1(n_320),
.B2(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_149),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_149),
.B(n_297),
.C(n_322),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_149),
.B(n_195),
.C(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_149),
.A2(n_194),
.B1(n_195),
.B2(n_324),
.Y(n_409)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_153),
.B(n_431),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_168),
.B(n_186),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_155),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_156),
.A2(n_167),
.B1(n_168),
.B2(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_156),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_158),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B(n_164),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_164),
.A2(n_180),
.A3(n_268),
.B1(n_272),
.B2(n_276),
.Y(n_267)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_166),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_167),
.A2(n_168),
.B1(n_186),
.B2(n_187),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_169),
.A2(n_251),
.B1(n_364),
.B2(n_370),
.Y(n_363)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_175),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_177),
.B(n_230),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_182),
.Y(n_296)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_208),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_194),
.A2(n_195),
.B1(n_237),
.B2(n_245),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_195),
.B(n_237),
.C(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_207),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_207),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_207),
.B(n_245),
.C(n_334),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_427),
.B(n_433),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

AO221x1_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_357),
.B1(n_359),
.B2(n_420),
.C(n_426),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_328),
.B(n_356),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_312),
.B(n_327),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_264),
.B(n_311),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_247),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_219),
.B(n_247),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_220),
.B(n_238),
.C(n_245),
.Y(n_326)
);

XOR2x2_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_221),
.B(n_228),
.Y(n_315)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_251),
.B1(n_252),
.B2(n_259),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_245),
.B2(n_246),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_237),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_237),
.A2(n_245),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_238),
.A2(n_246),
.B1(n_267),
.B2(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_238),
.B(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_238),
.A2(n_246),
.B1(n_387),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_263),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_248),
.A2(n_249),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_315),
.C(n_317),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_248),
.A2(n_249),
.B1(n_363),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_249),
.B(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_302),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_250),
.A2(n_283),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_298),
.B(n_300),
.Y(n_297)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_258),
.Y(n_367)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_286),
.B(n_310),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_282),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_266),
.B(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_283),
.B(n_341),
.Y(n_401)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_305),
.B(n_309),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_301),
.B(n_304),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_297),
.A2(n_306),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_300),
.A2(n_364),
.B(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_326),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_317),
.B1(n_318),
.B2(n_325),
.Y(n_313)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_330),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_337),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_338),
.C(n_339),
.Y(n_406)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_404),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_394),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_379),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_360),
.B(n_379),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_375),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_361),
.B(n_376),
.C(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_382),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.C(n_385),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_383),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_391),
.C(n_392),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_402),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_402),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_400),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_398),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_416),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_407),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_412),
.C(n_414),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_414),
.B2(n_415),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_416),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_419),
.Y(n_421)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B(n_424),
.C(n_425),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_430),
.Y(n_433)
);


endmodule