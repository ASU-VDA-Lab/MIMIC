module fake_jpeg_24789_n_322 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_8),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_50),
.Y(n_69)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_60),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_38),
.B1(n_30),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_27),
.B1(n_24),
.B2(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_24),
.B1(n_36),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_20),
.B1(n_36),
.B2(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_47),
.B1(n_45),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_78),
.B(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_39),
.B(n_37),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_69),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_41),
.A2(n_29),
.B1(n_31),
.B2(n_2),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_86),
.B1(n_11),
.B2(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_29),
.B1(n_1),
.B2(n_3),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_92),
.A2(n_72),
.B1(n_57),
.B2(n_6),
.Y(n_153)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_100),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_98),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_102),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_11),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_119),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_109),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_76),
.B1(n_88),
.B2(n_87),
.Y(n_138)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_73),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_69),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_69),
.B1(n_64),
.B2(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_149),
.B1(n_97),
.B2(n_92),
.Y(n_166)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_68),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_153),
.B1(n_92),
.B2(n_109),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_81),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_63),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_55),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_4),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_70),
.B1(n_57),
.B2(n_62),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_104),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_111),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_72),
.A3(n_55),
.B1(n_7),
.B2(n_8),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_104),
.B(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_173),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_111),
.B(n_115),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_160),
.A2(n_172),
.B(n_179),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_165),
.B(n_129),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_166),
.B1(n_170),
.B2(n_174),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_106),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_113),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_92),
.B1(n_101),
.B2(n_97),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_121),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_96),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_93),
.B1(n_113),
.B2(n_91),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_133),
.A2(n_91),
.B1(n_94),
.B2(n_117),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_189),
.B1(n_138),
.B2(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_150),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_184),
.A2(n_150),
.B1(n_127),
.B2(n_145),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_137),
.B(n_141),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_157),
.B(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_98),
.Y(n_187)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_94),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_125),
.B(n_142),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_189),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_130),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_198),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_202),
.B(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_155),
.C(n_152),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_201),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_156),
.B1(n_152),
.B2(n_142),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_219),
.B1(n_179),
.B2(n_190),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_213),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_152),
.B(n_129),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_214),
.B(n_220),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_127),
.B1(n_136),
.B2(n_135),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_168),
.B(n_178),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_157),
.Y(n_213)
);

NOR2x1p5_ASAP7_75t_SL g214 ( 
.A(n_172),
.B(n_5),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_136),
.B1(n_135),
.B2(n_13),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_165),
.B(n_11),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_234),
.B(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_186),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_203),
.B1(n_164),
.B2(n_170),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_181),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_160),
.C(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_236),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_171),
.B(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_180),
.B(n_172),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_195),
.A2(n_169),
.B(n_159),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_204),
.B1(n_215),
.B2(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_244),
.Y(n_255)
);

NAND2x1p5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_173),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_159),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_243),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_193),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_253),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_215),
.B1(n_175),
.B2(n_187),
.Y(n_276)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_252),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_227),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_259),
.B1(n_228),
.B2(n_234),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_238),
.B(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_205),
.B1(n_198),
.B2(n_204),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_209),
.C(n_169),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_243),
.C(n_240),
.Y(n_271)
);

AOI221xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_230),
.B1(n_221),
.B2(n_176),
.C(n_174),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_275),
.Y(n_285)
);

OAI31xp33_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_236),
.A3(n_222),
.B(n_229),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_231),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_248),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_250),
.B1(n_258),
.B2(n_254),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_229),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_246),
.B1(n_262),
.B2(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.C(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_208),
.C(n_240),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_279),
.B1(n_256),
.B2(n_245),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_182),
.C(n_173),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_183),
.B1(n_135),
.B2(n_136),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_191),
.C(n_13),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_259),
.Y(n_286)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_269),
.B1(n_278),
.B2(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_291),
.B1(n_292),
.B2(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_255),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_277),
.B1(n_251),
.B2(n_265),
.Y(n_291)
);

FAx1_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_12),
.CI(n_13),
.CON(n_293),
.SN(n_293)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_267),
.B(n_266),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_293),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_286),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_271),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_287),
.B1(n_283),
.B2(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_285),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_313),
.B1(n_304),
.B2(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_297),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_300),
.B1(n_281),
.B2(n_285),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_306),
.B(n_307),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_14),
.A3(n_15),
.B1(n_17),
.B2(n_282),
.C1(n_293),
.C2(n_317),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_310),
.B(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_14),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_14),
.Y(n_322)
);


endmodule