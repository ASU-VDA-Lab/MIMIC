module real_aes_8547_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g575 ( .A1(n_0), .A2(n_175), .B(n_576), .C(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_1), .B(n_521), .Y(n_580) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_2), .B(n_114), .C(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g128 ( .A(n_2), .Y(n_128) );
INVx1_ASAP7_75t_L g209 ( .A(n_3), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_4), .B(n_167), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_5), .A2(n_490), .B(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_6), .A2(n_152), .B(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_36), .B1(n_161), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_8), .B(n_152), .Y(n_178) );
AND2x6_ASAP7_75t_L g176 ( .A(n_9), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_10), .A2(n_176), .B(n_480), .C(n_482), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_11), .A2(n_461), .B1(n_753), .B2(n_754), .C1(n_763), .C2(n_767), .Y(n_460) );
INVx1_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_12), .B(n_37), .Y(n_129) );
INVx1_ASAP7_75t_L g157 ( .A(n_13), .Y(n_157) );
INVx1_ASAP7_75t_L g202 ( .A(n_14), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_15), .B(n_165), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_16), .B(n_167), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_17), .B(n_153), .Y(n_214) );
AO32x2_ASAP7_75t_L g236 ( .A1(n_18), .A2(n_152), .A3(n_182), .B1(n_193), .B2(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_19), .B(n_161), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_20), .B(n_153), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_21), .A2(n_56), .B1(n_161), .B2(n_239), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g261 ( .A1(n_22), .A2(n_84), .B1(n_161), .B2(n_165), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_23), .B(n_161), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_24), .A2(n_193), .B(n_480), .C(n_541), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_25), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_25), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_26), .A2(n_193), .B(n_480), .C(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_27), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_28), .B(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_29), .A2(n_490), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_30), .B(n_195), .Y(n_233) );
INVx2_ASAP7_75t_L g163 ( .A(n_31), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_32), .A2(n_492), .B(n_500), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_33), .B(n_161), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_34), .B(n_195), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_35), .B(n_247), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_37), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_38), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_39), .B(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_40), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_41), .A2(n_80), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_41), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_42), .B(n_167), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_43), .B(n_490), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g141 ( .A1(n_44), .A2(n_81), .B1(n_142), .B2(n_143), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_44), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_45), .A2(n_492), .B(n_494), .C(n_500), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_46), .A2(n_758), .B1(n_761), .B2(n_762), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_46), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_47), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g577 ( .A(n_48), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_49), .A2(n_93), .B1(n_239), .B2(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g495 ( .A(n_50), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_51), .B(n_161), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_52), .B(n_161), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_53), .A2(n_132), .B1(n_133), .B2(n_136), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_53), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_54), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_55), .B(n_173), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g218 ( .A1(n_57), .A2(n_61), .B1(n_161), .B2(n_165), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_58), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_59), .B(n_161), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_60), .B(n_161), .Y(n_244) );
INVx1_ASAP7_75t_L g177 ( .A(n_62), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_63), .B(n_490), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_64), .B(n_521), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_65), .A2(n_173), .B(n_205), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_66), .B(n_161), .Y(n_210) );
INVx1_ASAP7_75t_L g156 ( .A(n_67), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_69), .B(n_167), .Y(n_531) );
AO32x2_ASAP7_75t_L g257 ( .A1(n_70), .A2(n_152), .A3(n_193), .B1(n_258), .B2(n_262), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_71), .B(n_168), .Y(n_483) );
INVx1_ASAP7_75t_L g188 ( .A(n_72), .Y(n_188) );
INVx1_ASAP7_75t_L g228 ( .A(n_73), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_74), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_75), .B(n_497), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_76), .A2(n_480), .B(n_500), .C(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_77), .B(n_165), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_78), .Y(n_516) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_80), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_81), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_81), .A2(n_143), .B1(n_144), .B2(n_454), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_82), .A2(n_89), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_82), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_83), .B(n_496), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_85), .B(n_239), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_86), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_87), .B(n_165), .Y(n_232) );
INVx2_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_89), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_90), .B(n_192), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_91), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
OR2x2_ASAP7_75t_L g125 ( .A(n_92), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g465 ( .A(n_92), .B(n_127), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_94), .A2(n_104), .B1(n_165), .B2(n_166), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_95), .B(n_490), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_96), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_97), .A2(n_106), .B1(n_118), .B2(n_772), .Y(n_105) );
INVxp67_ASAP7_75t_L g519 ( .A(n_98), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_99), .B(n_165), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_100), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g476 ( .A(n_101), .Y(n_476) );
INVx1_ASAP7_75t_L g554 ( .A(n_102), .Y(n_554) );
AND2x2_ASAP7_75t_L g502 ( .A(n_103), .B(n_195), .Y(n_502) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g772 ( .A(n_108), .Y(n_772) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g752 ( .A(n_114), .B(n_127), .Y(n_752) );
NOR2x2_ASAP7_75t_L g769 ( .A(n_114), .B(n_126), .Y(n_769) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_459), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g771 ( .A(n_121), .Y(n_771) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_130), .B(n_455), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g458 ( .A(n_125), .Y(n_458) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
XOR2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_135), .B(n_219), .Y(n_558) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B1(n_144), .B2(n_454), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g454 ( .A(n_144), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_378), .Y(n_144) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_336), .Y(n_145) );
NOR4xp25_ASAP7_75t_L g146 ( .A(n_147), .B(n_276), .C(n_312), .D(n_326), .Y(n_146) );
OAI221xp5_ASAP7_75t_SL g147 ( .A1(n_148), .A2(n_220), .B1(n_252), .B2(n_263), .C(n_267), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_148), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_196), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_179), .Y(n_150) );
AND2x2_ASAP7_75t_L g273 ( .A(n_151), .B(n_180), .Y(n_273) );
INVx3_ASAP7_75t_L g281 ( .A(n_151), .Y(n_281) );
AND2x2_ASAP7_75t_L g335 ( .A(n_151), .B(n_199), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_151), .B(n_198), .Y(n_371) );
AND2x2_ASAP7_75t_L g429 ( .A(n_151), .B(n_291), .Y(n_429) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_158), .B(n_178), .Y(n_151) );
INVx4_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_152), .A2(n_507), .B(n_508), .Y(n_506) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_152), .Y(n_513) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_154), .B(n_155), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_170), .B(n_176), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_164), .B(n_167), .Y(n_159) );
INVx3_ASAP7_75t_L g227 ( .A(n_161), .Y(n_227) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_161), .Y(n_556) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
BUFx3_ASAP7_75t_L g260 ( .A(n_162), .Y(n_260) );
AND2x6_ASAP7_75t_L g480 ( .A(n_162), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
INVx2_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g175 ( .A(n_167), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_185), .B(n_186), .Y(n_184) );
O2A1O1Ixp5_ASAP7_75t_SL g226 ( .A1(n_167), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_167), .B(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g258 ( .A1(n_168), .A2(n_192), .B1(n_259), .B2(n_261), .Y(n_258) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
INVx1_ASAP7_75t_L g247 ( .A(n_169), .Y(n_247) );
AND2x2_ASAP7_75t_L g478 ( .A(n_169), .B(n_174), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_169), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_175), .Y(n_170) );
INVx2_ASAP7_75t_L g189 ( .A(n_173), .Y(n_189) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_175), .A2(n_189), .B(n_209), .C(n_210), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_175), .A2(n_192), .B1(n_217), .B2(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_175), .A2(n_192), .B1(n_238), .B2(n_240), .Y(n_237) );
BUFx3_ASAP7_75t_L g193 ( .A(n_176), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_176), .A2(n_201), .B(n_208), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_176), .A2(n_226), .B(n_230), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_176), .A2(n_243), .B(n_248), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_176), .B(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g490 ( .A(n_176), .B(n_478), .Y(n_490) );
INVx4_ASAP7_75t_SL g501 ( .A(n_176), .Y(n_501) );
AND2x2_ASAP7_75t_L g264 ( .A(n_179), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g278 ( .A(n_179), .B(n_199), .Y(n_278) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_180), .B(n_199), .Y(n_293) );
AND2x2_ASAP7_75t_L g305 ( .A(n_180), .B(n_281), .Y(n_305) );
OR2x2_ASAP7_75t_L g307 ( .A(n_180), .B(n_265), .Y(n_307) );
AND2x2_ASAP7_75t_L g342 ( .A(n_180), .B(n_265), .Y(n_342) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_180), .Y(n_387) );
INVx1_ASAP7_75t_L g395 ( .A(n_180), .Y(n_395) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B(n_194), .Y(n_180) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_181), .A2(n_200), .B(n_211), .Y(n_199) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_182), .B(n_486), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_193), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .C(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_189), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_191), .A2(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx4_ASAP7_75t_L g578 ( .A(n_192), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_193), .B(n_216), .C(n_219), .Y(n_215) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_195), .A2(n_225), .B(n_233), .Y(n_224) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_195), .A2(n_242), .B(n_251), .Y(n_241) );
INVx2_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_195), .A2(n_489), .B(n_491), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_195), .A2(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g547 ( .A(n_195), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_196), .A2(n_313), .B1(n_317), .B2(n_321), .C(n_322), .Y(n_312) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g272 ( .A(n_197), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
INVx2_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
AND2x2_ASAP7_75t_L g324 ( .A(n_198), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g343 ( .A(n_198), .B(n_281), .Y(n_343) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g406 ( .A(n_199), .B(n_281), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .C(n_205), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_203), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_203), .A2(n_510), .B(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_205), .A2(n_554), .B(n_555), .C(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_206), .A2(n_231), .B(n_232), .Y(n_230) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g497 ( .A(n_207), .Y(n_497) );
AND2x2_ASAP7_75t_L g328 ( .A(n_212), .B(n_273), .Y(n_328) );
OAI322xp33_ASAP7_75t_L g396 ( .A1(n_212), .A2(n_352), .A3(n_397), .B1(n_399), .B2(n_402), .C1(n_404), .C2(n_408), .Y(n_396) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_213), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
AND2x2_ASAP7_75t_L g401 ( .A(n_213), .B(n_281), .Y(n_401) );
AND2x2_ASAP7_75t_L g433 ( .A(n_213), .B(n_305), .Y(n_433) );
OR2x2_ASAP7_75t_L g436 ( .A(n_213), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
AO21x1_ASAP7_75t_L g265 ( .A1(n_216), .A2(n_219), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_219), .A2(n_475), .B(n_485), .Y(n_474) );
INVx3_ASAP7_75t_L g521 ( .A(n_219), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_219), .B(n_533), .Y(n_532) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_219), .A2(n_551), .B(n_558), .Y(n_550) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_234), .Y(n_221) );
INVx1_ASAP7_75t_L g449 ( .A(n_222), .Y(n_449) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g254 ( .A(n_223), .B(n_241), .Y(n_254) );
INVx2_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g311 ( .A(n_224), .Y(n_311) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_224), .Y(n_319) );
OR2x2_ASAP7_75t_L g443 ( .A(n_224), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g268 ( .A(n_234), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g308 ( .A(n_234), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g360 ( .A(n_234), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
AND2x2_ASAP7_75t_L g255 ( .A(n_235), .B(n_256), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g315 ( .A(n_235), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g369 ( .A(n_235), .B(n_257), .Y(n_369) );
OR2x2_ASAP7_75t_L g377 ( .A(n_235), .B(n_311), .Y(n_377) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx2_ASAP7_75t_L g286 ( .A(n_236), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_236), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g320 ( .A(n_236), .B(n_241), .Y(n_320) );
AND2x2_ASAP7_75t_L g384 ( .A(n_236), .B(n_257), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_241), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_241), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
INVx1_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g314 ( .A(n_241), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_241), .Y(n_392) );
INVx1_ASAP7_75t_L g444 ( .A(n_241), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_246), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g421 ( .A(n_253), .B(n_330), .Y(n_421) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g348 ( .A(n_255), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g447 ( .A(n_255), .B(n_382), .Y(n_447) );
INVx1_ASAP7_75t_L g269 ( .A(n_256), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_256), .B(n_289), .Y(n_295) );
BUFx2_ASAP7_75t_L g354 ( .A(n_256), .Y(n_354) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_257), .Y(n_275) );
INVx1_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_260), .Y(n_499) );
INVx2_ASAP7_75t_L g579 ( .A(n_260), .Y(n_579) );
INVx1_ASAP7_75t_L g544 ( .A(n_262), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g423 ( .A(n_263), .B(n_270), .Y(n_423) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI32xp33_ASAP7_75t_L g267 ( .A1(n_264), .A2(n_268), .A3(n_270), .B1(n_272), .B2(n_274), .Y(n_267) );
AND2x2_ASAP7_75t_L g407 ( .A(n_264), .B(n_280), .Y(n_407) );
AND2x2_ASAP7_75t_L g445 ( .A(n_264), .B(n_343), .Y(n_445) );
INVx1_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_269), .B(n_331), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_270), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_270), .B(n_273), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_270), .B(n_342), .Y(n_424) );
OR2x2_ASAP7_75t_L g438 ( .A(n_270), .B(n_307), .Y(n_438) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g365 ( .A(n_271), .B(n_273), .Y(n_365) );
OR2x2_ASAP7_75t_L g374 ( .A(n_271), .B(n_361), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_273), .B(n_324), .Y(n_346) );
INVx2_ASAP7_75t_L g361 ( .A(n_275), .Y(n_361) );
OR2x2_ASAP7_75t_L g376 ( .A(n_275), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g391 ( .A(n_275), .B(n_392), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_275), .A2(n_368), .B(n_449), .C(n_450), .Y(n_448) );
OAI321xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_282), .A3(n_287), .B1(n_290), .B2(n_294), .C(n_298), .Y(n_276) );
INVx1_ASAP7_75t_L g389 ( .A(n_277), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g400 ( .A(n_278), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g352 ( .A(n_280), .Y(n_352) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_281), .B(n_395), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_282), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
AND2x2_ASAP7_75t_L g357 ( .A(n_284), .B(n_331), .Y(n_357) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_285), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_287), .A2(n_328), .B(n_373), .C(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g339 ( .A(n_289), .B(n_296), .Y(n_339) );
BUFx2_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
INVx1_ASAP7_75t_L g364 ( .A(n_289), .Y(n_364) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g370 ( .A(n_292), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g453 ( .A(n_292), .Y(n_453) );
INVx1_ASAP7_75t_L g446 ( .A(n_293), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g299 ( .A(n_295), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g403 ( .A(n_295), .B(n_320), .Y(n_403) );
INVx1_ASAP7_75t_L g332 ( .A(n_296), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_303), .B1(n_306), .B2(n_308), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_300), .B(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g368 ( .A(n_301), .B(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_302), .B(n_311), .Y(n_331) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g323 ( .A(n_305), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g333 ( .A(n_307), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_310), .A2(n_428), .B1(n_430), .B2(n_431), .C(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g316 ( .A(n_311), .Y(n_316) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_311), .Y(n_382) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_314), .B(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_315), .A2(n_320), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_318), .B(n_328), .Y(n_425) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g394 ( .A(n_319), .Y(n_394) );
AND2x2_ASAP7_75t_L g353 ( .A(n_320), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g442 ( .A(n_320), .Y(n_442) );
INVx1_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
INVx1_ASAP7_75t_L g413 ( .A(n_324), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_332), .B2(n_333), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_330), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_331), .B(n_369), .Y(n_435) );
OR2x2_ASAP7_75t_L g408 ( .A(n_332), .B(n_361), .Y(n_408) );
INVx1_ASAP7_75t_L g347 ( .A(n_333), .Y(n_347) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_335), .B(n_386), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_355), .C(n_366), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_344), .C(n_350), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_339), .A2(n_410), .B1(n_414), .B2(n_417), .C(n_419), .Y(n_409) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g351 ( .A(n_342), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g405 ( .A(n_342), .B(n_406), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g390 ( .A1(n_343), .A2(n_391), .B(n_393), .C(n_395), .Y(n_390) );
INVx2_ASAP7_75t_L g437 ( .A(n_343), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_347), .B(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_369), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_359), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_365), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_360), .B(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_365), .B(n_452), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B(n_372), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g393 ( .A(n_369), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND4x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_409), .C(n_426), .D(n_448), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_396), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_385), .B(n_388), .C(n_390), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_384), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_395), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
INVx2_ASAP7_75t_SL g418 ( .A(n_406), .Y(n_418) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g431 ( .A(n_416), .Y(n_431) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g426 ( .A(n_427), .B(n_434), .Y(n_426) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .B1(n_438), .B2(n_439), .C(n_440), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_455), .B(n_460), .C(n_770), .Y(n_459) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_463), .B1(n_466), .B2(n_750), .Y(n_461) );
INVx1_ASAP7_75t_L g764 ( .A(n_462), .Y(n_764) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g765 ( .A(n_464), .Y(n_765) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_467), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
OR3x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_648), .C(n_713), .Y(n_467) );
NAND4xp25_ASAP7_75t_SL g468 ( .A(n_469), .B(n_589), .C(n_615), .D(n_638), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_522), .B1(n_559), .B2(n_566), .C(n_581), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_471), .A2(n_582), .B1(n_606), .B2(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_503), .Y(n_471) );
INVx1_ASAP7_75t_SL g642 ( .A(n_472), .Y(n_642) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_487), .Y(n_472) );
OR2x2_ASAP7_75t_L g564 ( .A(n_473), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g584 ( .A(n_473), .B(n_504), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_473), .B(n_512), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_473), .B(n_487), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_473), .B(n_562), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_473), .B(n_613), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_473), .B(n_503), .Y(n_735) );
AOI211xp5_ASAP7_75t_SL g746 ( .A1(n_473), .A2(n_652), .B(n_747), .C(n_748), .Y(n_746) );
INVx5_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_474), .B(n_504), .Y(n_618) );
AND2x2_ASAP7_75t_L g621 ( .A(n_474), .B(n_505), .Y(n_621) );
OR2x2_ASAP7_75t_L g666 ( .A(n_474), .B(n_504), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_474), .B(n_512), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_479), .Y(n_475) );
INVx5_ASAP7_75t_L g493 ( .A(n_480), .Y(n_493) );
INVx5_ASAP7_75t_SL g565 ( .A(n_487), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_487), .B(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_487), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_487), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g701 ( .A(n_487), .B(n_512), .Y(n_701) );
OR2x2_ASAP7_75t_L g707 ( .A(n_487), .B(n_597), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_487), .B(n_657), .Y(n_716) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_502), .Y(n_487) );
BUFx2_ASAP7_75t_L g539 ( .A(n_490), .Y(n_539) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_493), .A2(n_501), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g573 ( .A1(n_493), .A2(n_501), .B(n_574), .C(n_575), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_498), .C(n_499), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_496), .A2(n_499), .B(n_530), .C(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
AND2x2_ASAP7_75t_L g598 ( .A(n_504), .B(n_565), .Y(n_598) );
INVx1_ASAP7_75t_SL g611 ( .A(n_504), .Y(n_611) );
OR2x2_ASAP7_75t_L g646 ( .A(n_504), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g652 ( .A(n_504), .B(n_512), .Y(n_652) );
AND2x2_ASAP7_75t_L g710 ( .A(n_504), .B(n_562), .Y(n_710) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_505), .B(n_565), .Y(n_637) );
INVx3_ASAP7_75t_L g562 ( .A(n_512), .Y(n_562) );
OR2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_565), .Y(n_603) );
AND2x2_ASAP7_75t_L g613 ( .A(n_512), .B(n_611), .Y(n_613) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_512), .Y(n_661) );
AND2x2_ASAP7_75t_L g670 ( .A(n_512), .B(n_584), .Y(n_670) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_520), .Y(n_512) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_521), .A2(n_572), .B(n_580), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_522), .A2(n_687), .B1(n_689), .B2(n_691), .C(n_694), .Y(n_686) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .Y(n_523) );
AND2x2_ASAP7_75t_L g660 ( .A(n_524), .B(n_641), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_524), .B(n_719), .Y(n_723) );
OR2x2_ASAP7_75t_L g744 ( .A(n_524), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_524), .B(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx5_ASAP7_75t_L g591 ( .A(n_525), .Y(n_591) );
AND2x2_ASAP7_75t_L g668 ( .A(n_525), .B(n_536), .Y(n_668) );
AND2x2_ASAP7_75t_L g729 ( .A(n_525), .B(n_608), .Y(n_729) );
AND2x2_ASAP7_75t_L g742 ( .A(n_525), .B(n_562), .Y(n_742) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_532), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_548), .Y(n_534) );
AND2x4_ASAP7_75t_L g569 ( .A(n_535), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_535), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g594 ( .A(n_535), .Y(n_594) );
AND2x2_ASAP7_75t_L g663 ( .A(n_535), .B(n_641), .Y(n_663) );
AND2x2_ASAP7_75t_L g673 ( .A(n_535), .B(n_591), .Y(n_673) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_535), .Y(n_681) );
AND2x2_ASAP7_75t_L g693 ( .A(n_535), .B(n_571), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_535), .B(n_625), .Y(n_697) );
AND2x2_ASAP7_75t_L g734 ( .A(n_535), .B(n_729), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_535), .B(n_608), .Y(n_745) );
OR2x2_ASAP7_75t_L g747 ( .A(n_535), .B(n_683), .Y(n_747) );
INVx5_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g633 ( .A(n_536), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g643 ( .A(n_536), .B(n_588), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_536), .B(n_571), .Y(n_655) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_536), .Y(n_685) );
AND2x4_ASAP7_75t_L g719 ( .A(n_536), .B(n_570), .Y(n_719) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
AOI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_540), .B(n_544), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
BUFx2_ASAP7_75t_L g568 ( .A(n_548), .Y(n_568) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g608 ( .A(n_549), .Y(n_608) );
AND2x2_ASAP7_75t_L g641 ( .A(n_549), .B(n_571), .Y(n_641) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g588 ( .A(n_550), .B(n_571), .Y(n_588) );
BUFx2_ASAP7_75t_L g634 ( .A(n_550), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_557), .Y(n_551) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_561), .B(n_642), .Y(n_721) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_562), .B(n_584), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_562), .B(n_565), .Y(n_623) );
AND2x2_ASAP7_75t_L g678 ( .A(n_562), .B(n_614), .Y(n_678) );
AOI221xp5_ASAP7_75t_SL g615 ( .A1(n_563), .A2(n_616), .B1(n_624), .B2(n_626), .C(n_630), .Y(n_615) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g610 ( .A(n_564), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g651 ( .A(n_564), .B(n_652), .Y(n_651) );
OAI321xp33_ASAP7_75t_L g658 ( .A1(n_564), .A2(n_617), .A3(n_659), .B1(n_661), .B2(n_662), .C(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_565), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_568), .B(n_719), .Y(n_737) );
AND2x2_ASAP7_75t_L g624 ( .A(n_569), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_569), .B(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_570), .Y(n_600) );
AND2x2_ASAP7_75t_L g607 ( .A(n_570), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_570), .B(n_682), .Y(n_712) );
INVx1_ASAP7_75t_L g749 ( .A(n_570), .Y(n_749) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_586), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_583), .A2(n_693), .B(n_742), .C(n_743), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_584), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_584), .B(n_622), .Y(n_688) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g631 ( .A(n_588), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_588), .B(n_591), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_588), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_588), .B(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B1(n_604), .B2(n_609), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g605 ( .A(n_591), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g628 ( .A(n_591), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g640 ( .A(n_591), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_591), .B(n_634), .Y(n_676) );
OR2x2_ASAP7_75t_L g683 ( .A(n_591), .B(n_608), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_591), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g733 ( .A(n_591), .B(n_719), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_599), .B2(n_601), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g639 ( .A(n_594), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_597), .A2(n_612), .B1(n_680), .B2(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g727 ( .A(n_598), .Y(n_727) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_602), .A2(n_639), .B1(n_642), .B2(n_643), .C(n_644), .Y(n_638) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g617 ( .A(n_603), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_607), .B(n_673), .Y(n_705) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_608), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_608), .Y(n_629) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
AND2x2_ASAP7_75t_L g656 ( .A(n_614), .B(n_657), .Y(n_656) );
NAND2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g700 ( .A(n_621), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_624), .A2(n_650), .B1(n_653), .B2(n_656), .C(n_658), .Y(n_649) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_628), .B(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B(n_635), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_635), .Y(n_732) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OR2x2_ASAP7_75t_L g674 ( .A(n_637), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g695 ( .A(n_640), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_640), .B(n_700), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_643), .B(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_667), .C(n_686), .D(n_699), .Y(n_648) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g657 ( .A(n_652), .Y(n_657) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g690 ( .A(n_661), .B(n_666), .Y(n_690) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_671), .C(n_679), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g738 ( .A1(n_669), .A2(n_711), .B(n_739), .C(n_746), .Y(n_738) );
INVx1_ASAP7_75t_SL g698 ( .A(n_670), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g702 ( .A(n_676), .Y(n_702) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_682), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_682), .B(n_693), .Y(n_726) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g703 ( .A(n_693), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .Y(n_694) );
INVxp33_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .A3(n_703), .B1(n_704), .B2(n_706), .C1(n_708), .C2(n_711), .Y(n_699) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND3xp33_ASAP7_75t_SL g713 ( .A(n_714), .B(n_731), .C(n_738), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_720), .B2(n_722), .C(n_724), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g730 ( .A(n_719), .Y(n_730) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_735), .C(n_736), .Y(n_731) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g766 ( .A(n_751), .Y(n_766) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g761 ( .A(n_758), .Y(n_761) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
endmodule