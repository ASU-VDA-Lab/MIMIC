module fake_jpeg_21687_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_40),
.B1(n_31),
.B2(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_27),
.B1(n_40),
.B2(n_31),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_69),
.Y(n_85)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_74),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_61),
.B1(n_77),
.B2(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_51),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_34),
.C(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_34),
.B(n_25),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_92),
.B(n_55),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_53),
.B1(n_41),
.B2(n_32),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_77),
.B1(n_65),
.B2(n_72),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_93),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_34),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_69),
.B1(n_57),
.B2(n_58),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_98),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_25),
.B(n_22),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_25),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_17),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_104),
.B1(n_108),
.B2(n_118),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_65),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_55),
.B1(n_74),
.B2(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_16),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_71),
.B(n_70),
.C(n_28),
.Y(n_113)
);

OAI22x1_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_82),
.B1(n_101),
.B2(n_87),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_22),
.B1(n_18),
.B2(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_14),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_80),
.C(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.C(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_86),
.C(n_88),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_92),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_105),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_93),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_85),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_131),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_87),
.C(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_93),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_81),
.B(n_117),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_113),
.B1(n_105),
.B2(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_154),
.C(n_122),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_148),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_113),
.B1(n_118),
.B2(n_103),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_28),
.B1(n_21),
.B2(n_4),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_113),
.B1(n_109),
.B2(n_85),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_157),
.B(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g156 ( 
.A(n_136),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_132),
.B1(n_125),
.B2(n_136),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_164),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_125),
.B1(n_123),
.B2(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_157),
.Y(n_173)
);

AOI321xp33_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_126),
.A3(n_137),
.B1(n_129),
.B2(n_124),
.C(n_117),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_150),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_21),
.B1(n_13),
.B2(n_11),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_21),
.C(n_13),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_154),
.C(n_148),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_2),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_165),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_159),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_147),
.C(n_3),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_176),
.B1(n_178),
.B2(n_170),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_164),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_163),
.B(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_180),
.B1(n_183),
.B2(n_6),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_4),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_192),
.B(n_194),
.Y(n_195)
);

AOI21x1_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_5),
.B(n_6),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_189),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_196),
.B(n_6),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.C(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_8),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_9),
.Y(n_201)
);


endmodule