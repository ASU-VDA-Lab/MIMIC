module fake_netlist_6_3455_n_407 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_66, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_65, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_407);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_66;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_65;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_407;

wire n_91;
wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_68;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_125;
wire n_384;
wire n_297;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_78;
wire n_84;
wire n_392;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_67;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_71;
wire n_74;
wire n_229;
wire n_305;
wire n_72;
wire n_173;
wire n_250;
wire n_372;
wire n_111;
wire n_314;
wire n_378;
wire n_377;
wire n_183;
wire n_79;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_73;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_397;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_70;
wire n_234;
wire n_381;
wire n_82;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_80;
wire n_196;
wire n_402;
wire n_352;
wire n_107;
wire n_89;
wire n_374;
wire n_366;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_69;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_83;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_90;
wire n_347;
wire n_328;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_75;
wire n_401;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_81;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVxp33_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_4),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_6),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_8),
.Y(n_93)
);

INVxp33_ASAP7_75t_SL g94 ( 
.A(n_27),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

INVxp33_ASAP7_75t_SL g96 ( 
.A(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_22),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_55),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_52),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_14),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_23),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_34),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_3),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_54),
.Y(n_110)
);

INVxp33_ASAP7_75t_SL g111 ( 
.A(n_56),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_53),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_40),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_30),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_41),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_13),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_62),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_R g138 ( 
.A(n_96),
.B(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_95),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_1),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_2),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_R g159 ( 
.A(n_119),
.B(n_2),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_113),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_R g179 ( 
.A(n_122),
.B(n_5),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_117),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_71),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_85),
.Y(n_186)
);

NAND2x1p5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_89),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_96),
.B1(n_94),
.B2(n_111),
.Y(n_189)
);

NAND2x1p5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_121),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_182),
.B1(n_137),
.B2(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_97),
.Y(n_195)
);

AO22x2_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_118),
.B1(n_112),
.B2(n_104),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_92),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

OAI221xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_116),
.B1(n_125),
.B2(n_75),
.C(n_126),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2x1p5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_111),
.Y(n_203)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_160),
.B(n_124),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_150),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_101),
.Y(n_209)
);

NAND2x1p5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_94),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_68),
.Y(n_211)
);

OR2x2_ASAP7_75t_SL g212 ( 
.A(n_163),
.B(n_124),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_5),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_26),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_25),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_140),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_148),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g225 ( 
.A1(n_153),
.A2(n_10),
.B1(n_12),
.B2(n_16),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_R g230 ( 
.A(n_134),
.B(n_17),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_157),
.B(n_31),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_159),
.B(n_35),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_171),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_185),
.B1(n_183),
.B2(n_151),
.Y(n_237)
);

OR2x6_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_217),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_164),
.B(n_138),
.C(n_159),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_165),
.Y(n_241)
);

NOR2x1_ASAP7_75t_R g242 ( 
.A(n_205),
.B(n_133),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_162),
.B(n_175),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_138),
.B(n_179),
.C(n_129),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_173),
.B1(n_170),
.B2(n_132),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_156),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_156),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_141),
.B1(n_45),
.B2(n_63),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_43),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_141),
.B(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_190),
.B(n_195),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_212),
.B1(n_210),
.B2(n_203),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_197),
.B(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_203),
.B(n_210),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_190),
.B(n_195),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_198),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_193),
.A2(n_194),
.B(n_197),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_193),
.A2(n_194),
.B(n_207),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_216),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_234),
.B(n_231),
.C(n_224),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_196),
.A2(n_188),
.B(n_214),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_214),
.B(n_230),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_214),
.B(n_230),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_196),
.A2(n_188),
.B(n_192),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_196),
.A2(n_219),
.B(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_208),
.B(n_213),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_215),
.B(n_213),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_208),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_208),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_215),
.Y(n_285)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_225),
.B(n_278),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_275),
.B1(n_257),
.B2(n_261),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_254),
.B1(n_277),
.B2(n_238),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_254),
.A2(n_238),
.B1(n_251),
.B2(n_282),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_241),
.B(n_250),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_281),
.B(n_263),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_262),
.A2(n_260),
.B(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_268),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

AO32x2_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_237),
.A3(n_238),
.B1(n_276),
.B2(n_248),
.Y(n_298)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_243),
.A2(n_266),
.B(n_265),
.Y(n_299)
);

OR2x6_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_239),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_237),
.B1(n_247),
.B2(n_245),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_253),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_267),
.A2(n_264),
.B(n_253),
.C(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

OAI222xp33_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_189),
.B1(n_238),
.B2(n_249),
.C1(n_222),
.C2(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

AOI221xp5_ASAP7_75t_L g310 ( 
.A1(n_237),
.A2(n_189),
.B1(n_245),
.B2(n_254),
.C(n_96),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_270),
.A2(n_278),
.B(n_256),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_278),
.B(n_256),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_273),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_274),
.A2(n_189),
.B(n_278),
.C(n_270),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_270),
.A2(n_278),
.B(n_279),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_270),
.A2(n_278),
.B(n_256),
.Y(n_323)
);

OAI211xp5_ASAP7_75t_L g324 ( 
.A1(n_244),
.A2(n_189),
.B(n_168),
.C(n_200),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_274),
.A2(n_273),
.B1(n_189),
.B2(n_278),
.Y(n_325)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_310),
.B(n_302),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_287),
.A2(n_325),
.B1(n_318),
.B2(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_320),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_319),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_288),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_304),
.B1(n_321),
.B2(n_297),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_285),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_297),
.B1(n_286),
.B2(n_299),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_291),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_R g340 ( 
.A(n_303),
.B(n_319),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_288),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_292),
.C(n_308),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_289),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_323),
.B(n_295),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_314),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_SL g348 ( 
.A(n_306),
.B(n_293),
.C(n_309),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_322),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_R g351 ( 
.A(n_305),
.B(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

AO21x2_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_348),
.B(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_329),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_305),
.B(n_307),
.Y(n_356)
);

OAI221xp5_ASAP7_75t_L g357 ( 
.A1(n_342),
.A2(n_298),
.B1(n_301),
.B2(n_316),
.C(n_314),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_312),
.B(n_294),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_305),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

AOI222xp33_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_294),
.B1(n_298),
.B2(n_301),
.C1(n_316),
.C2(n_337),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_298),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_333),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_333),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_330),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_339),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_339),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_361),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_357),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_356),
.B1(n_343),
.B2(n_344),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_350),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_373),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_353),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_374),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_365),
.Y(n_385)
);

OAI321xp33_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_370),
.A3(n_364),
.B1(n_368),
.B2(n_371),
.C(n_372),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_365),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_340),
.B1(n_370),
.B2(n_351),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_385),
.B(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_384),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_384),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

AO22x2_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_389),
.B1(n_379),
.B2(n_383),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_395),
.A2(n_358),
.B(n_334),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_389),
.B(n_376),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_391),
.C(n_396),
.Y(n_400)
);

NAND2x1_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_393),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_400),
.Y(n_402)
);

AOI31xp33_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_399),
.A3(n_331),
.B(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_403),
.Y(n_404)
);

OAI322xp33_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_398),
.A3(n_402),
.B1(n_354),
.B2(n_341),
.C1(n_298),
.C2(n_381),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_341),
.B1(n_381),
.B2(n_368),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_350),
.B(n_349),
.Y(n_407)
);


endmodule