module fake_jpeg_71_n_155 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_155);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_49),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_19),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_26),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_28),
.B1(n_30),
.B2(n_18),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_73),
.B1(n_23),
.B2(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_14),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_26),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_80),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_69),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_39),
.B(n_50),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_91),
.C(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_77),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_10),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_48),
.B1(n_42),
.B2(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_20),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_20),
.B1(n_34),
.B2(n_8),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_20),
.B1(n_7),
.B2(n_9),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_72),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_77),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_60),
.B(n_71),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_60),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_112),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_57),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_69),
.A3(n_67),
.B1(n_70),
.B2(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_5),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_91),
.C(n_82),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_79),
.C(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_106),
.B1(n_99),
.B2(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_130),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_122),
.B1(n_101),
.B2(n_124),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_133),
.B1(n_123),
.B2(n_126),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_119),
.B(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_99),
.B1(n_111),
.B2(n_104),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_117),
.Y(n_141)
);

OAI321xp33_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_140),
.A3(n_134),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_139),
.C(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND4xp25_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_131),
.C(n_133),
.D(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_144),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_142),
.B1(n_137),
.B2(n_116),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_149),
.A3(n_142),
.B1(n_86),
.B2(n_138),
.C1(n_80),
.C2(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_70),
.A3(n_61),
.B1(n_67),
.B2(n_80),
.C1(n_7),
.C2(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_152),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_61),
.Y(n_155)
);


endmodule