module fake_jpeg_12242_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_25),
.C(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_31),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_33),
.B1(n_37),
.B2(n_34),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_48),
.B1(n_53),
.B2(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_36),
.B1(n_37),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_36),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_22),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_64),
.B(n_2),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_1),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_1),
.B(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_74),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_3),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_68),
.B1(n_65),
.B2(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_79),
.B1(n_67),
.B2(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_59),
.B1(n_53),
.B2(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_66),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_82),
.B(n_76),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_77),
.B(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_73),
.B1(n_78),
.B2(n_75),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_4),
.B(n_5),
.Y(n_86)
);

AOI211xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_87)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_14),
.Y(n_88)
);


endmodule