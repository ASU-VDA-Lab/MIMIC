module real_jpeg_21209_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_0),
.A2(n_25),
.B1(n_27),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_0),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_162),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_162),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_162),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_2),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_135),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_135),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_135),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_24),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_14),
.B(n_49),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_166),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_4),
.A2(n_80),
.B1(n_153),
.B2(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_4),
.B(n_197),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_4),
.B(n_27),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_4),
.A2(n_27),
.B(n_248),
.Y(n_252)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_6),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_168),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_168),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_168),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_7),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_9),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_31),
.B1(n_48),
.B2(n_49),
.Y(n_174)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_94),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.C(n_76),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_20),
.B(n_67),
.CI(n_76),
.CON(n_139),
.SN(n_139)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_21),
.A2(n_22),
.B1(n_96),
.B2(n_109),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_22),
.B(n_39),
.C(n_55),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_23),
.A2(n_28),
.B1(n_90),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_23),
.A2(n_90),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_23),
.A2(n_90),
.B1(n_134),
.B2(n_179),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_24),
.B(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_24),
.A2(n_35),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_25),
.A2(n_36),
.B1(n_165),
.B2(n_172),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g247 ( 
.A1(n_25),
.A2(n_42),
.A3(n_59),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_26),
.B(n_27),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g165 ( 
.A(n_30),
.B(n_166),
.CON(n_165),
.SN(n_165)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_40),
.B1(n_101),
.B2(n_107),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_41),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_41),
.A2(n_47),
.B1(n_86),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_41),
.A2(n_51),
.B(n_87),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_41),
.A2(n_47),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_41),
.A2(n_47),
.B1(n_219),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_41),
.A2(n_47),
.B1(n_239),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_41),
.A2(n_71),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_43),
.A2(n_50),
.B(n_166),
.C(n_215),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g249 ( 
.A(n_43),
.B(n_58),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_47),
.A2(n_73),
.B(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_47),
.B(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_48),
.B(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_65),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_56),
.A2(n_103),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_56),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_56),
.A2(n_65),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_57),
.A2(n_61),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_57),
.A2(n_61),
.B1(n_196),
.B2(n_252),
.Y(n_251)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_69),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_66),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_68),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_89),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_78),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_80),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_80),
.A2(n_150),
.B1(n_153),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_80),
.A2(n_82),
.B1(n_208),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_80),
.A2(n_128),
.B(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_81),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_81),
.A2(n_84),
.B(n_152),
.Y(n_246)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_108),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_317),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_139),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_115),
.B(n_139),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_116),
.B(n_120),
.Y(n_315)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_121),
.A2(n_122),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.C(n_137),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_123),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_124),
.B(n_130),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_153),
.B(n_174),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_139),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_311),
.B(n_316),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_299),
.B(n_310),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_199),
.B(n_278),
.C(n_298),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_184),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_144),
.B(n_184),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_169),
.B2(n_183),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_147),
.B(n_156),
.C(n_183),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_155),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_148),
.B(n_155),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_153),
.B(n_166),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_164),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_170),
.B(n_176),
.C(n_181),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_194),
.B(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_277),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_272),
.B(n_276),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_260),
.B(n_271),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_242),
.B(n_259),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_231),
.B(n_241),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_220),
.B(n_230),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_212),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_216),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_229),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_250),
.B1(n_257),
.B2(n_258),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_245),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_269),
.C(n_270),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_296),
.B2(n_297),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.C(n_297),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_295),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_293),
.C(n_295),
.Y(n_309)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_307),
.C(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);


endmodule