module fake_ariane_284_n_2002 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2002);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2002;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_363;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_43),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_107),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_116),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_72),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_76),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_126),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_11),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_93),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_3),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_29),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_86),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_51),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_44),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_53),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_68),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_47),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_121),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_189),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_141),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_74),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_138),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_39),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_11),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_105),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_52),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_160),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_96),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_155),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_34),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_169),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_112),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_25),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_101),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_127),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_5),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_44),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_87),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_163),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_148),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_187),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_90),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_89),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_99),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_109),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_120),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_113),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_136),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_94),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_142),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_173),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_55),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_184),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_4),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_150),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_192),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_165),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_135),
.Y(n_303)
);

BUFx8_ASAP7_75t_SL g304 ( 
.A(n_65),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_122),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_54),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_42),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_77),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_168),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_62),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_191),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_63),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_54),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_114),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_98),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_202),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_115),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_159),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_119),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_123),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_15),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_58),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_111),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_143),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_59),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_130),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_58),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_18),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_70),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_80),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_166),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_88),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_91),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_144),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_34),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_199),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_8),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_108),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_26),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_13),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_81),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_16),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_158),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_25),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_12),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_41),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_172),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_46),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_60),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_179),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_134),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_82),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_117),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_9),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_53),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_92),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_131),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_20),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_17),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_190),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_27),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_13),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_33),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_125),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_151),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_66),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_49),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_14),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_193),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_200),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_64),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_183),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_20),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_162),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_49),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_30),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_69),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_79),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_52),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_157),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_197),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_28),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_37),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_38),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_167),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_174),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_194),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_42),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_97),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_32),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_73),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_128),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_171),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_43),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_15),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_145),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_27),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_29),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_154),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_2),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_304),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_318),
.B(n_0),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_302),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_236),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_243),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_302),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_254),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_318),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_326),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_240),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_268),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_326),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_206),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_337),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_319),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_384),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_206),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_214),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_236),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_385),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_214),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_334),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_227),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_227),
.B(n_0),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_242),
.B(n_2),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_228),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_228),
.B(n_3),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_335),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_387),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_236),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_397),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_232),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_232),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_290),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_236),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_290),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_248),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_239),
.Y(n_456)
);

BUFx6f_ASAP7_75t_SL g457 ( 
.A(n_274),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_239),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_207),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_211),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_216),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_249),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_307),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_249),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_252),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_252),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_270),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_217),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_231),
.B(n_235),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_236),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_314),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_259),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_270),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_231),
.B(n_5),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_235),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_255),
.B(n_6),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_285),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_285),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_299),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_238),
.B(n_10),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_299),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_346),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_306),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_306),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_219),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_220),
.Y(n_486)
);

INVx4_ASAP7_75t_R g487 ( 
.A(n_274),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_331),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_221),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_222),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_331),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_226),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_238),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_230),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_332),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_234),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_259),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_247),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_257),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_266),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_272),
.Y(n_501)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_295),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_340),
.B(n_14),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_273),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_280),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_241),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_241),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_332),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_339),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_339),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_281),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_259),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_R g513 ( 
.A(n_208),
.B(n_67),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_292),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_293),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_490),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_469),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_423),
.B(n_338),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_476),
.B(n_259),
.Y(n_525)
);

BUFx8_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_470),
.B(n_348),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_423),
.B(n_259),
.Y(n_528)
);

BUFx8_ASAP7_75t_L g529 ( 
.A(n_457),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_492),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_497),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_432),
.B(n_233),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_472),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_512),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_494),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_503),
.B(n_323),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_264),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_412),
.B(n_229),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_437),
.B(n_440),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_475),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_475),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_493),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_457),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_506),
.B(n_233),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_261),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_462),
.B(n_429),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_434),
.B(n_261),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_413),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_477),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_416),
.B(n_264),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_425),
.B(n_269),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_478),
.B(n_323),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_479),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_481),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_483),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_427),
.B(n_265),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_430),
.B(n_265),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_419),
.Y(n_583)
);

CKINVDCx8_ASAP7_75t_R g584 ( 
.A(n_411),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_491),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_509),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_422),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_502),
.B(n_323),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_442),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_438),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_441),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_473),
.B(n_269),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_450),
.B(n_480),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_439),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_535),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_551),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_522),
.B(n_459),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_551),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_518),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_551),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_424),
.C(n_422),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

INVxp33_ASAP7_75t_L g610 ( 
.A(n_544),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_535),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_542),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_551),
.B(n_283),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_548),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_501),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_424),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_551),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_594),
.B(n_426),
.Y(n_620)
);

CKINVDCx6p67_ASAP7_75t_R g621 ( 
.A(n_540),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_561),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_540),
.B(n_459),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_594),
.B(n_426),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_535),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_594),
.B(n_460),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_460),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_548),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_593),
.B(n_461),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_552),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_549),
.B(n_282),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_461),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_540),
.B(n_485),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_548),
.A2(n_591),
.B1(n_573),
.B2(n_546),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_552),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_549),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_596),
.B(n_486),
.C(n_485),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_552),
.Y(n_644)
);

BUFx6f_ASAP7_75t_SL g645 ( 
.A(n_548),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_549),
.B(n_486),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_557),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_536),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_584),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_552),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

INVx4_ASAP7_75t_SL g653 ( 
.A(n_524),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_556),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_526),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_542),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_556),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_556),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_591),
.A2(n_496),
.B1(n_498),
.B2(n_489),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_557),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_560),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_560),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_596),
.B(n_520),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_523),
.B(n_489),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_560),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_541),
.Y(n_671)
);

CKINVDCx6p67_ASAP7_75t_R g672 ( 
.A(n_540),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_523),
.B(n_496),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_516),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_516),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_516),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_534),
.B(n_498),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_541),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_524),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_500),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_540),
.B(n_500),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_550),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_533),
.B(n_504),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_571),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_521),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_530),
.B(n_504),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_521),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_550),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_540),
.B(n_511),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_553),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_530),
.B(n_511),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_546),
.B(n_454),
.C(n_452),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_526),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_521),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_528),
.B(n_282),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_526),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_562),
.B(n_350),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_530),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_540),
.B(n_499),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_562),
.B(n_455),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_518),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_562),
.A2(n_350),
.B1(n_360),
.B2(n_351),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_521),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_554),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_526),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_573),
.A2(n_353),
.B1(n_364),
.B2(n_349),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_540),
.B(n_505),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_521),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_565),
.B(n_351),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_538),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_531),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_538),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_539),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_540),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_530),
.A2(n_532),
.B1(n_537),
.B2(n_565),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_532),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_555),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_532),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_528),
.B(n_288),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_532),
.B(n_215),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_597),
.B(n_514),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_531),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_399),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_537),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_517),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_537),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_565),
.A2(n_365),
.B1(n_395),
.B2(n_370),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_517),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_517),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_567),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_571),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_517),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_527),
.B(n_402),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_571),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_527),
.B(n_288),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_517),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_584),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_571),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_517),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_547),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_526),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_283),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_565),
.B(n_443),
.Y(n_746)
);

AND2x2_ASAP7_75t_SL g747 ( 
.A(n_555),
.B(n_229),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_517),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_534),
.B(n_360),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_654),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_626),
.B(n_567),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_743),
.B(n_586),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_618),
.B(n_583),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_615),
.B(n_555),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_642),
.A2(n_586),
.B(n_563),
.C(n_569),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_736),
.B(n_586),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_650),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_622),
.B(n_586),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_654),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_622),
.B(n_586),
.Y(n_761)
);

INVx8_ASAP7_75t_L g762 ( 
.A(n_740),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_620),
.B(n_583),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_701),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_655),
.B(n_589),
.Y(n_765)
);

BUFx4_ASAP7_75t_L g766 ( 
.A(n_740),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_658),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_658),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_628),
.B(n_589),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_604),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_606),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_571),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_645),
.A2(n_568),
.B1(n_578),
.B2(n_566),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_671),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_628),
.B(n_443),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_600),
.B(n_529),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_612),
.A2(n_545),
.B(n_525),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_600),
.B(n_529),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_604),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_671),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_723),
.A2(n_547),
.B(n_564),
.C(n_563),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_529),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_740),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_665),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_660),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_668),
.B(n_529),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_660),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_697),
.B(n_531),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_662),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_652),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_645),
.A2(n_555),
.B1(n_569),
.B2(n_564),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_624),
.B(n_525),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_650),
.B(n_444),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_615),
.B(n_528),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_686),
.A2(n_545),
.B(n_566),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_696),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_SL g797 ( 
.A(n_663),
.B(n_444),
.C(n_411),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_738),
.B(n_598),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_678),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_662),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_691),
.A2(n_568),
.B(n_566),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_655),
.B(n_570),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_645),
.A2(n_568),
.B1(n_578),
.B2(n_566),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_646),
.B(n_570),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_635),
.B(n_665),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_599),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_599),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_610),
.A2(n_647),
.B1(n_697),
.B2(n_673),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_682),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_602),
.Y(n_812)
);

NOR2x1p5_ASAP7_75t_L g813 ( 
.A(n_608),
.B(n_576),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_634),
.B(n_577),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_603),
.B(n_577),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_615),
.B(n_543),
.Y(n_816)
);

NOR3xp33_ASAP7_75t_L g817 ( 
.A(n_643),
.B(n_543),
.C(n_393),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_697),
.A2(n_580),
.B1(n_590),
.B2(n_543),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_747),
.B(n_528),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_602),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_693),
.B(n_415),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_733),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_713),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_688),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_724),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_688),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_747),
.B(n_528),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_698),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_634),
.B(n_524),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_611),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_634),
.B(n_580),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_634),
.B(n_590),
.Y(n_832)
);

AO221x1_ASAP7_75t_L g833 ( 
.A1(n_708),
.A2(n_323),
.B1(n_365),
.B2(n_366),
.C(n_367),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_669),
.A2(n_578),
.B(n_581),
.C(n_568),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_747),
.B(n_528),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_634),
.B(n_534),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_656),
.A2(n_657),
.B(n_661),
.C(n_659),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_634),
.B(n_558),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_680),
.B(n_592),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_683),
.A2(n_581),
.B(n_585),
.C(n_578),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_611),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_690),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_690),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_702),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_677),
.B(n_558),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_677),
.B(n_558),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_652),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_616),
.B(n_592),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_746),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_702),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_656),
.B(n_581),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_733),
.B(n_595),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_733),
.B(n_595),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_693),
.B(n_581),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_692),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_722),
.B(n_559),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_652),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_559),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_697),
.A2(n_588),
.B1(n_587),
.B2(n_585),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_707),
.B(n_559),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_707),
.B(n_585),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_749),
.B(n_367),
.C(n_366),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_700),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_711),
.B(n_592),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_711),
.B(n_705),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_629),
.B(n_585),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_711),
.B(n_592),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_625),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_625),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_706),
.B(n_575),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_639),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_706),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_639),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_641),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_698),
.B(n_575),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_749),
.B(n_375),
.C(n_370),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_417),
.Y(n_878)
);

AND2x6_ASAP7_75t_SL g879 ( 
.A(n_664),
.B(n_375),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_698),
.B(n_575),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_718),
.B(n_575),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_718),
.B(n_575),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_718),
.B(n_575),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_720),
.B(n_587),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_699),
.B(n_572),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_720),
.B(n_587),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_727),
.B(n_587),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_727),
.B(n_588),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_695),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_641),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_696),
.B(n_574),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_657),
.A2(n_588),
.B(n_579),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_709),
.B(n_572),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_659),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_648),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_661),
.B(n_579),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_744),
.B(n_574),
.Y(n_897)
);

O2A1O1Ixp5_ASAP7_75t_L g898 ( 
.A1(n_729),
.A2(n_588),
.B(n_582),
.C(n_258),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_695),
.A2(n_574),
.B1(n_582),
.B2(n_395),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_744),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_729),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_664),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_685),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_666),
.A2(n_404),
.B(n_405),
.C(n_305),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_623),
.B(n_294),
.Y(n_905)
);

INVx8_ASAP7_75t_L g906 ( 
.A(n_695),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_695),
.A2(n_404),
.B1(n_405),
.B2(n_316),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_717),
.B(n_305),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_648),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_666),
.B(n_316),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_652),
.B(n_317),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_667),
.B(n_317),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_621),
.B(n_421),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_667),
.B(n_320),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_649),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_670),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_652),
.B(n_320),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_649),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_823),
.B(n_703),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_866),
.A2(n_681),
.B1(n_689),
.B2(n_637),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_837),
.A2(n_605),
.B(n_601),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_774),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_757),
.A2(n_605),
.B(n_601),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_753),
.A2(n_614),
.B(n_607),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_851),
.A2(n_803),
.B(n_792),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_851),
.A2(n_614),
.B(n_607),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_849),
.B(n_428),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_825),
.B(n_436),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_752),
.B(n_695),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_752),
.B(n_695),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_754),
.B(n_763),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_754),
.B(n_695),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_763),
.B(n_719),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_896),
.A2(n_619),
.B(n_617),
.Y(n_934)
);

AND2x6_ASAP7_75t_L g935 ( 
.A(n_796),
.B(n_670),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_848),
.B(n_721),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_848),
.B(n_721),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_765),
.B(n_719),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_793),
.B(n_446),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_815),
.B(n_721),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_896),
.A2(n_619),
.B(n_617),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_810),
.B(n_719),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_808),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_884),
.A2(n_887),
.B(n_886),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_806),
.A2(n_687),
.B(n_694),
.C(n_685),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_769),
.B(n_684),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_770),
.B(n_453),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_762),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_780),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_795),
.A2(n_630),
.B(n_627),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_815),
.B(n_721),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_786),
.B(n_684),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_857),
.B(n_721),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_796),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_779),
.B(n_463),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_782),
.B(n_684),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_888),
.A2(n_716),
.B(n_630),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_898),
.A2(n_632),
.B(n_627),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_771),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_822),
.B(n_684),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_772),
.A2(n_716),
.B(n_633),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_839),
.A2(n_716),
.B(n_633),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_790),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_777),
.A2(n_636),
.B(n_632),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_906),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_859),
.B(n_721),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_807),
.B(n_471),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_798),
.B(n_730),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_891),
.B(n_653),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_809),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_758),
.B(n_482),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_799),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_885),
.A2(n_737),
.B(n_734),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_885),
.A2(n_750),
.B(n_651),
.C(n_609),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_801),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_790),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_764),
.B(n_609),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_845),
.B(n_712),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_894),
.A2(n_636),
.B(n_644),
.C(n_640),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_784),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_839),
.A2(n_644),
.B(n_640),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_809),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_759),
.A2(n_737),
.B(n_734),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_846),
.B(n_714),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_781),
.A2(n_710),
.B(n_687),
.C(n_694),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_893),
.B(n_714),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_761),
.A2(n_741),
.B(n_651),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_775),
.B(n_715),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_790),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_802),
.A2(n_621),
.B1(n_672),
.B2(n_651),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_818),
.B(n_684),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_819),
.A2(n_750),
.B1(n_609),
.B2(n_741),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_864),
.A2(n_710),
.B(n_704),
.C(n_675),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_900),
.B(n_704),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_878),
.B(n_726),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_834),
.A2(n_731),
.B(n_728),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_811),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_899),
.B(n_726),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_840),
.A2(n_731),
.B(n_728),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_899),
.B(n_674),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_812),
.Y(n_1001)
);

NOR2xp67_ASAP7_75t_L g1002 ( 
.A(n_797),
.B(n_674),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_824),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_812),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_876),
.A2(n_735),
.B(n_732),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_826),
.B(n_676),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_842),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_880),
.A2(n_735),
.B(n_732),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_843),
.B(n_676),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_881),
.A2(n_742),
.B(n_739),
.Y(n_1010)
);

CKINVDCx10_ASAP7_75t_R g1011 ( 
.A(n_788),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_844),
.A2(n_672),
.B1(n_297),
.B2(n_298),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_850),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_819),
.A2(n_745),
.B1(n_613),
.B2(n_742),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_905),
.A2(n_748),
.B(n_739),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_882),
.A2(n_748),
.B(n_613),
.Y(n_1016)
);

AND2x2_ASAP7_75t_SL g1017 ( 
.A(n_821),
.B(n_487),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_788),
.B(n_309),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_883),
.A2(n_745),
.B(n_330),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_853),
.B(n_873),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_756),
.A2(n_330),
.B(n_329),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_892),
.A2(n_210),
.B(n_209),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_836),
.B(n_838),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_906),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_901),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_860),
.B(n_311),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_856),
.B(n_313),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_814),
.A2(n_336),
.B(n_329),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_831),
.A2(n_352),
.B(n_336),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_832),
.A2(n_355),
.B(n_352),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_863),
.B(n_322),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_820),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_877),
.B(n_324),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_891),
.B(n_325),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_762),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_871),
.A2(n_358),
.B(n_355),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_852),
.B(n_854),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_902),
.A2(n_362),
.B(n_358),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_897),
.B(n_341),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_368),
.B(n_362),
.Y(n_1040)
);

CKINVDCx10_ASAP7_75t_R g1041 ( 
.A(n_766),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_897),
.B(n_513),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_906),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_827),
.A2(n_373),
.B(n_368),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_820),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_830),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_751),
.A2(n_386),
.B(n_373),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_907),
.B(n_343),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_751),
.A2(n_396),
.B(n_386),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_762),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_827),
.A2(n_213),
.B(n_212),
.Y(n_1051)
);

AND2x6_ASAP7_75t_L g1052 ( 
.A(n_790),
.B(n_653),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_907),
.B(n_344),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_865),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_905),
.A2(n_396),
.B(n_278),
.C(n_277),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_SL g1056 ( 
.A1(n_911),
.A2(n_262),
.B(n_401),
.C(n_260),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_900),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_835),
.A2(n_256),
.B(n_409),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_835),
.A2(n_253),
.B(n_406),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_816),
.B(n_354),
.C(n_410),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_913),
.B(n_361),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_889),
.B(n_804),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_913),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_813),
.Y(n_1064)
);

BUFx4f_ASAP7_75t_L g1065 ( 
.A(n_783),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_776),
.B(n_653),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_778),
.B(n_369),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_868),
.B(n_371),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_794),
.B(n_379),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_828),
.A2(n_245),
.B(n_403),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_817),
.B(n_381),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_794),
.B(n_388),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_828),
.A2(n_237),
.B(n_218),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_760),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_904),
.A2(n_394),
.B(n_356),
.C(n_392),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_910),
.A2(n_391),
.B(n_398),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_773),
.B(n_653),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_783),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_773),
.B(n_400),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_805),
.A2(n_408),
.B1(n_407),
.B2(n_323),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_783),
.B(n_16),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_805),
.B(n_223),
.Y(n_1082)
);

AO21x2_ASAP7_75t_L g1083 ( 
.A1(n_912),
.A2(n_519),
.B(n_517),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_SL g1084 ( 
.A(n_855),
.B(n_679),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_767),
.A2(n_519),
.B(n_679),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_861),
.B(n_224),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_867),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_833),
.B(n_519),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_914),
.A2(n_791),
.B(n_917),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_908),
.B(n_225),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_903),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_768),
.B(n_244),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_847),
.B(n_679),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_768),
.B(n_21),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_879),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_847),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_785),
.A2(n_519),
.B(n_246),
.C(n_321),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_785),
.B(n_250),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_847),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_787),
.A2(n_519),
.B(n_679),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_944),
.A2(n_858),
.B(n_847),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_931),
.A2(n_858),
.B1(n_789),
.B2(n_800),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_988),
.B(n_787),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_995),
.B(n_789),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_SL g1105 ( 
.A1(n_956),
.A2(n_917),
.B(n_911),
.C(n_862),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_933),
.A2(n_858),
.B(n_829),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1027),
.B(n_1054),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_947),
.B(n_800),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_1057),
.B(n_755),
.Y(n_1109)
);

OR2x6_ASAP7_75t_SL g1110 ( 
.A(n_1081),
.B(n_251),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_922),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_948),
.B(n_858),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_955),
.B(n_271),
.C(n_263),
.Y(n_1113)
);

BUFx8_ASAP7_75t_SL g1114 ( 
.A(n_1095),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_936),
.A2(n_755),
.B(n_918),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_973),
.A2(n_918),
.B(n_915),
.C(n_909),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_927),
.A2(n_380),
.B1(n_287),
.B2(n_286),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1041),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_967),
.B(n_841),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1050),
.B(n_841),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_919),
.A2(n_915),
.B1(n_909),
.B2(n_895),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_980),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_943),
.Y(n_1123)
);

AO32x1_ASAP7_75t_L g1124 ( 
.A1(n_1088),
.A2(n_1080),
.A3(n_920),
.B1(n_1025),
.B2(n_972),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_948),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_928),
.B(n_869),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_949),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_929),
.A2(n_890),
.B1(n_875),
.B2(n_874),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_968),
.B(n_869),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_975),
.B(n_890),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_930),
.A2(n_875),
.B1(n_874),
.B2(n_872),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_959),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_1003),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1035),
.B(n_870),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_L g1135 ( 
.A(n_1042),
.B(n_872),
.C(n_870),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_971),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_932),
.A2(n_519),
.B(n_276),
.C(n_275),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_970),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_939),
.B(n_279),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_937),
.A2(n_342),
.B(n_289),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_982),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1071),
.A2(n_524),
.B1(n_679),
.B2(n_519),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1007),
.B(n_1013),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_934),
.A2(n_345),
.B(n_291),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_969),
.B(n_519),
.Y(n_1145)
);

OR2x4_ASAP7_75t_L g1146 ( 
.A(n_1037),
.B(n_23),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_969),
.B(n_679),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1064),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1018),
.B(n_284),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_940),
.B(n_296),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1094),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1055),
.A2(n_347),
.B(n_390),
.C(n_389),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1031),
.A2(n_24),
.B(n_30),
.C(n_31),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1011),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1069),
.A2(n_524),
.B1(n_383),
.B2(n_382),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1020),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1001),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_934),
.A2(n_300),
.B(n_378),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_R g1160 ( 
.A(n_1061),
.B(n_301),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1091),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1065),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_954),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1072),
.A2(n_524),
.B1(n_377),
.B2(n_374),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1065),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_986),
.B(n_32),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1063),
.B(n_35),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1004),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_SL g1169 ( 
.A(n_963),
.B(n_303),
.Y(n_1169)
);

O2A1O1Ixp5_ASAP7_75t_L g1170 ( 
.A1(n_952),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_941),
.A2(n_308),
.B(n_372),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1079),
.A2(n_310),
.B1(n_312),
.B2(n_315),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_951),
.A2(n_363),
.B(n_359),
.C(n_357),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1078),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1017),
.B(n_40),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_977),
.B(n_327),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_941),
.A2(n_925),
.B(n_1016),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_963),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1044),
.A2(n_333),
.B(n_338),
.C(n_283),
.Y(n_1180)
);

HAxp5_ASAP7_75t_L g1181 ( 
.A(n_1033),
.B(n_41),
.CON(n_1181),
.SN(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_981),
.A2(n_338),
.B(n_85),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1075),
.A2(n_1044),
.B1(n_1087),
.B2(n_1053),
.C(n_1048),
.Y(n_1183)
);

AND2x6_ASAP7_75t_L g1184 ( 
.A(n_965),
.B(n_338),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_978),
.B(n_45),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_925),
.A2(n_283),
.B(n_524),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1012),
.B(n_283),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_923),
.A2(n_962),
.B(n_924),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1057),
.B(n_100),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1034),
.B(n_46),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1026),
.A2(n_524),
.B1(n_283),
.B2(n_50),
.Y(n_1191)
);

BUFx8_ASAP7_75t_L g1192 ( 
.A(n_935),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_984),
.B(n_47),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1068),
.B(n_48),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_935),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1002),
.A2(n_283),
.B(n_524),
.C(n_51),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1074),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_950),
.A2(n_283),
.B(n_524),
.Y(n_1198)
);

AO32x1_ASAP7_75t_L g1199 ( 
.A1(n_1032),
.A2(n_48),
.A3(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_SL g1200 ( 
.A(n_946),
.B(n_57),
.C(n_59),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_935),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1039),
.B(n_60),
.C(n_61),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_965),
.B(n_61),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1067),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_SL g1205 ( 
.A(n_1076),
.B(n_71),
.C(n_75),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1006),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_923),
.A2(n_78),
.B(n_83),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_953),
.B(n_84),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_1021),
.A2(n_102),
.B(n_104),
.C(n_106),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1009),
.A2(n_110),
.B1(n_124),
.B2(n_137),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1045),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1046),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_924),
.A2(n_146),
.B(n_147),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_966),
.B(n_152),
.C(n_170),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1005),
.A2(n_177),
.B(n_182),
.Y(n_1215)
);

OAI22x1_ASAP7_75t_L g1216 ( 
.A1(n_991),
.A2(n_185),
.B1(n_186),
.B2(n_201),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_985),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1000),
.A2(n_203),
.B1(n_998),
.B2(n_992),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1023),
.A2(n_1030),
.B1(n_1022),
.B2(n_1014),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1038),
.A2(n_1040),
.B(n_993),
.C(n_1047),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1052),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_935),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1082),
.A2(n_976),
.B1(n_963),
.B2(n_989),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_942),
.B(n_1096),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1049),
.B(n_1060),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1096),
.B(n_960),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_945),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1005),
.A2(n_1010),
.B(n_1008),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1008),
.A2(n_1010),
.B(n_957),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_976),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1024),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1038),
.B(n_1040),
.Y(n_1233)
);

BUFx8_ASAP7_75t_L g1234 ( 
.A(n_976),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_994),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_989),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1024),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_989),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1036),
.B(n_1099),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1043),
.B(n_1099),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1028),
.B(n_1029),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1089),
.A2(n_999),
.B(n_996),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1021),
.A2(n_1029),
.B1(n_1028),
.B2(n_974),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1019),
.A2(n_1015),
.B(n_1016),
.C(n_926),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_994),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_996),
.A2(n_999),
.B(n_964),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1052),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1052),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1052),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1092),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1052),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1246),
.A2(n_990),
.B(n_979),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1244),
.A2(n_1097),
.A3(n_1100),
.B(n_1085),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1221),
.B(n_1019),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1224),
.A2(n_1059),
.B(n_1058),
.C(n_1051),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1122),
.B(n_1098),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1107),
.B(n_1073),
.Y(n_1258)
);

BUFx2_ASAP7_75t_R g1259 ( 
.A(n_1118),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1186),
.A2(n_921),
.B(n_926),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1111),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_SL g1262 ( 
.A(n_1221),
.B(n_938),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1158),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1229),
.A2(n_921),
.B(n_1100),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1119),
.B(n_1070),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1127),
.Y(n_1266)
);

NOR4xp25_ASAP7_75t_L g1267 ( 
.A(n_1153),
.B(n_958),
.C(n_1062),
.D(n_1066),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1178),
.A2(n_983),
.B(n_1085),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1226),
.A2(n_961),
.B(n_987),
.C(n_1084),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1158),
.Y(n_1270)
);

INVx4_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1132),
.Y(n_1272)
);

NAND2x1_ASAP7_75t_L g1273 ( 
.A(n_1222),
.B(n_1093),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1056),
.B(n_1083),
.C(n_1183),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1133),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1234),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1242),
.A2(n_1188),
.B(n_1243),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1114),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1101),
.A2(n_1219),
.B(n_1178),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1198),
.A2(n_1116),
.B(n_1182),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1241),
.A2(n_1218),
.B(n_1220),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1129),
.A2(n_1137),
.A3(n_1180),
.B(n_1102),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1146),
.A2(n_1181),
.B1(n_1149),
.B2(n_1117),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1223),
.A2(n_1228),
.B(n_1239),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1215),
.B(n_1105),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1126),
.B(n_1136),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1194),
.A2(n_1204),
.B(n_1166),
.C(n_1190),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1117),
.B(n_1250),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1174),
.A2(n_1209),
.B(n_1193),
.C(n_1185),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1161),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1176),
.B(n_1167),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1151),
.B(n_1143),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1177),
.B(n_1200),
.C(n_1202),
.Y(n_1293)
);

AOI221xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1152),
.A2(n_1196),
.B1(n_1233),
.B2(n_1217),
.C(n_1171),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1148),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1247),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1221),
.B(n_1201),
.Y(n_1297)
);

NAND2xp33_ASAP7_75t_L g1298 ( 
.A(n_1248),
.B(n_1247),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1106),
.A2(n_1222),
.B(n_1150),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1208),
.A2(n_1213),
.B(n_1207),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1156),
.B(n_1139),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1165),
.B(n_1162),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1165),
.B(n_1162),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_1214),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1236),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1206),
.B(n_1104),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1155),
.A2(n_1164),
.B1(n_1195),
.B2(n_1203),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1138),
.A2(n_1141),
.B1(n_1157),
.B2(n_1212),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_1245),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1234),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1238),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_SL g1312 ( 
.A1(n_1235),
.A2(n_1130),
.B(n_1103),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1197),
.A2(n_1124),
.A3(n_1168),
.B(n_1211),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1205),
.B(n_1164),
.C(n_1155),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1247),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1175),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1203),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1134),
.B(n_1163),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1225),
.A2(n_1135),
.B(n_1113),
.C(n_1214),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1134),
.B(n_1172),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1124),
.A2(n_1120),
.B(n_1210),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1187),
.A2(n_1210),
.B(n_1170),
.C(n_1159),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1125),
.A2(n_1251),
.B1(n_1145),
.B2(n_1144),
.Y(n_1323)
);

AO32x2_ASAP7_75t_L g1324 ( 
.A1(n_1124),
.A2(n_1199),
.A3(n_1125),
.B1(n_1110),
.B2(n_1173),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1249),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1154),
.B(n_1231),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1147),
.B(n_1145),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1191),
.A2(n_1109),
.B(n_1140),
.C(n_1227),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1109),
.A2(n_1121),
.B(n_1240),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1189),
.A2(n_1252),
.B(n_1142),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1249),
.Y(n_1331)
);

NAND2xp33_ASAP7_75t_SL g1332 ( 
.A(n_1249),
.B(n_1169),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1252),
.A2(n_1120),
.B(n_1112),
.C(n_1237),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1112),
.A2(n_1237),
.B(n_1232),
.C(n_1147),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1179),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1232),
.A2(n_1192),
.B(n_1184),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1199),
.A2(n_1154),
.B1(n_1192),
.B2(n_1145),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1179),
.B(n_1184),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1184),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1199),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1122),
.B(n_784),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1156),
.B(n_807),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1224),
.A2(n_931),
.B(n_723),
.C(n_849),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1156),
.B(n_807),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1224),
.A2(n_931),
.B(n_723),
.C(n_849),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1244),
.A2(n_973),
.A3(n_1229),
.B(n_1089),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1111),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1156),
.B(n_807),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1107),
.B(n_650),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1123),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1247),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1355)
);

AOI221x1_ASAP7_75t_L g1356 ( 
.A1(n_1216),
.A2(n_1210),
.B1(n_1246),
.B2(n_1219),
.C(n_1243),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1156),
.B(n_807),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1224),
.A2(n_931),
.B(n_723),
.C(n_849),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1111),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1132),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1156),
.B(n_807),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1224),
.A2(n_931),
.B(n_723),
.C(n_849),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1229),
.A2(n_1230),
.B(n_973),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1234),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1118),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1107),
.B(n_849),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1107),
.B(n_650),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1181),
.A2(n_931),
.B(n_603),
.C(n_522),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1111),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1122),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1111),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1158),
.Y(n_1375)
);

AOI221x1_ASAP7_75t_L g1376 ( 
.A1(n_1216),
.A2(n_1210),
.B1(n_1246),
.B2(n_1219),
.C(n_1243),
.Y(n_1376)
);

AOI221x1_ASAP7_75t_L g1377 ( 
.A1(n_1216),
.A2(n_1210),
.B1(n_1246),
.B2(n_1219),
.C(n_1243),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1242),
.A2(n_1246),
.B(n_1229),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1158),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1156),
.B(n_807),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1119),
.B(n_807),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1119),
.B(n_807),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1111),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1107),
.B(n_650),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1118),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_SL g1388 ( 
.A1(n_1174),
.A2(n_931),
.B(n_933),
.C(n_930),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1123),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1107),
.B(n_650),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1234),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1165),
.B(n_1158),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1156),
.B(n_807),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1156),
.B(n_807),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1220),
.A2(n_937),
.B(n_936),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_973),
.A3(n_1229),
.B(n_1089),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1111),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1398)
);

OAI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1226),
.A2(n_931),
.B(n_522),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1132),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1186),
.A2(n_1229),
.B(n_1101),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1119),
.B(n_807),
.Y(n_1402)
);

BUFx4_ASAP7_75t_SL g1403 ( 
.A(n_1118),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1244),
.A2(n_973),
.A3(n_1229),
.B(n_1089),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1119),
.B(n_807),
.Y(n_1405)
);

OAI21xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1233),
.A2(n_931),
.B(n_827),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1224),
.A2(n_931),
.B(n_723),
.C(n_849),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1246),
.A2(n_1101),
.B(n_1188),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1158),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1340),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1283),
.A2(n_1288),
.B1(n_1399),
.B2(n_1314),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1283),
.A2(n_1314),
.B1(n_1336),
.B2(n_1291),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1368),
.A2(n_1293),
.B1(n_1399),
.B2(n_1307),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1325),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1293),
.A2(n_1301),
.B1(n_1382),
.B2(n_1383),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1261),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1345),
.A2(n_1364),
.B1(n_1407),
.B2(n_1359),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1266),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1311),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1402),
.A2(n_1405),
.B1(n_1258),
.B2(n_1338),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1349),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1403),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1265),
.A2(n_1338),
.B1(n_1352),
.B2(n_1389),
.Y(n_1423)
);

INVx3_ASAP7_75t_SL g1424 ( 
.A(n_1387),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1347),
.A2(n_1393),
.B1(n_1357),
.B2(n_1344),
.Y(n_1425)
);

INVx5_ASAP7_75t_L g1426 ( 
.A(n_1340),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1351),
.A2(n_1390),
.B1(n_1386),
.B2(n_1370),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1360),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1286),
.A2(n_1350),
.B1(n_1346),
.B2(n_1394),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1392),
.Y(n_1430)
);

BUFx8_ASAP7_75t_L g1431 ( 
.A(n_1367),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1372),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1374),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1363),
.A2(n_1381),
.B1(n_1371),
.B2(n_1281),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1406),
.A2(n_1304),
.B1(n_1306),
.B2(n_1292),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1356),
.A2(n_1376),
.B1(n_1377),
.B2(n_1257),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1305),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1304),
.A2(n_1330),
.B1(n_1321),
.B2(n_1341),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1353),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1384),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1397),
.A2(n_1395),
.B1(n_1317),
.B2(n_1295),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1316),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1276),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1287),
.A2(n_1319),
.B(n_1305),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1272),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1313),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1308),
.A2(n_1329),
.B1(n_1330),
.B2(n_1312),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1329),
.A2(n_1332),
.B1(n_1373),
.B2(n_1395),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1341),
.A2(n_1297),
.B1(n_1327),
.B2(n_1324),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1310),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1353),
.B(n_1337),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1297),
.A2(n_1324),
.B1(n_1279),
.B2(n_1318),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1324),
.A2(n_1320),
.B1(n_1323),
.B2(n_1309),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1335),
.Y(n_1454)
);

BUFx12f_ASAP7_75t_L g1455 ( 
.A(n_1366),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1284),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1326),
.B(n_1290),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1325),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1271),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1333),
.B(n_1267),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1362),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_1277),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1400),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1391),
.A2(n_1298),
.B1(n_1392),
.B2(n_1409),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1259),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1263),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1325),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1263),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1263),
.A2(n_1379),
.B1(n_1375),
.B2(n_1270),
.Y(n_1469)
);

BUFx2_ASAP7_75t_SL g1470 ( 
.A(n_1271),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1339),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1253),
.A2(n_1294),
.B1(n_1267),
.B2(n_1331),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1270),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1270),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1375),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1375),
.A2(n_1409),
.B1(n_1379),
.B2(n_1300),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1379),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1302),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1296),
.Y(n_1479)
);

BUFx4f_ASAP7_75t_SL g1480 ( 
.A(n_1296),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1315),
.A2(n_1255),
.B1(n_1303),
.B2(n_1262),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1294),
.A2(n_1315),
.B1(n_1268),
.B2(n_1365),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1378),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1334),
.A2(n_1255),
.B1(n_1273),
.B2(n_1328),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1299),
.A2(n_1268),
.B1(n_1365),
.B2(n_1285),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1264),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

BUFx2_ASAP7_75t_R g1488 ( 
.A(n_1388),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1289),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1256),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1396),
.B(n_1404),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1269),
.Y(n_1492)
);

BUFx4_ASAP7_75t_R g1493 ( 
.A(n_1322),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1396),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1260),
.A2(n_1280),
.B1(n_1408),
.B2(n_1369),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1343),
.A2(n_1380),
.B1(n_1398),
.B2(n_1385),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1404),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1254),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1274),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1354),
.A2(n_1361),
.B1(n_1355),
.B2(n_1358),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1254),
.B(n_1282),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1282),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1401),
.Y(n_1503)
);

CKINVDCx14_ASAP7_75t_R g1504 ( 
.A(n_1278),
.Y(n_1504)
);

BUFx10_ASAP7_75t_L g1505 ( 
.A(n_1387),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1261),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1283),
.A2(n_1288),
.B1(n_723),
.B2(n_927),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1325),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1261),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1399),
.A2(n_522),
.B(n_849),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1367),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1353),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1314),
.A2(n_1146),
.B1(n_931),
.B2(n_638),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1261),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1261),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1288),
.A2(n_1110),
.B1(n_939),
.B2(n_821),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1399),
.A2(n_931),
.B1(n_1283),
.B2(n_1293),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1261),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1348),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1283),
.A2(n_1314),
.B1(n_417),
.B2(n_421),
.Y(n_1520)
);

CKINVDCx11_ASAP7_75t_R g1521 ( 
.A(n_1367),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1367),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1283),
.A2(n_1288),
.B1(n_444),
.B2(n_443),
.Y(n_1523)
);

INVx6_ASAP7_75t_L g1524 ( 
.A(n_1353),
.Y(n_1524)
);

BUFx10_ASAP7_75t_L g1525 ( 
.A(n_1387),
.Y(n_1525)
);

INVx4_ASAP7_75t_L g1526 ( 
.A(n_1311),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1283),
.A2(n_1314),
.B1(n_417),
.B2(n_421),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1275),
.B(n_1399),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1342),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1325),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1311),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1348),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1399),
.A2(n_931),
.B1(n_1283),
.B2(n_1293),
.Y(n_1533)
);

INVx6_ASAP7_75t_L g1534 ( 
.A(n_1353),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1314),
.A2(n_1146),
.B1(n_931),
.B2(n_638),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1275),
.B(n_1399),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1367),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1311),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1283),
.A2(n_1288),
.B1(n_931),
.B2(n_1399),
.Y(n_1539)
);

INVx6_ASAP7_75t_L g1540 ( 
.A(n_1353),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1278),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1446),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1478),
.Y(n_1543)
);

INVx4_ASAP7_75t_SL g1544 ( 
.A(n_1492),
.Y(n_1544)
);

AO21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1460),
.A2(n_1420),
.B(n_1491),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1437),
.B(n_1507),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1496),
.A2(n_1485),
.B(n_1495),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1442),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1416),
.B(n_1418),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1421),
.B(n_1428),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1519),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1503),
.A2(n_1456),
.B(n_1462),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1487),
.B(n_1497),
.Y(n_1554)
);

AOI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1434),
.A2(n_1460),
.B(n_1491),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1520),
.A2(n_1527),
.B1(n_1499),
.B2(n_1411),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_SL g1557 ( 
.A(n_1431),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1532),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1529),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1532),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1528),
.Y(n_1561)
);

AO21x1_ASAP7_75t_SL g1562 ( 
.A1(n_1420),
.A2(n_1411),
.B(n_1501),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1502),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1432),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1494),
.B(n_1490),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1462),
.A2(n_1497),
.B(n_1487),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1490),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1528),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1483),
.A2(n_1498),
.B(n_1476),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1440),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1478),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1461),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1506),
.B(n_1509),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1424),
.B(n_1445),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1434),
.A2(n_1417),
.B(n_1536),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1514),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1517),
.A2(n_1533),
.B(n_1539),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1536),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1515),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1518),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1433),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1463),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1479),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1483),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1449),
.B(n_1438),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1492),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1465),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1492),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1490),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1500),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1410),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1457),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1426),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1500),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1429),
.B(n_1435),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1486),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1482),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1449),
.B(n_1438),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1466),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1476),
.A2(n_1484),
.B(n_1451),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1454),
.Y(n_1601)
);

CKINVDCx6p67_ASAP7_75t_R g1602 ( 
.A(n_1424),
.Y(n_1602)
);

AO21x1_ASAP7_75t_SL g1603 ( 
.A1(n_1435),
.A2(n_1441),
.B(n_1448),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1423),
.A2(n_1447),
.B(n_1441),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1471),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1451),
.A2(n_1417),
.B(n_1481),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1482),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1453),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1453),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1472),
.Y(n_1610)
);

INVx5_ASAP7_75t_L g1611 ( 
.A(n_1426),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1472),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1436),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1468),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1436),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1520),
.A2(n_1527),
.B1(n_1539),
.B2(n_1535),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1459),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1425),
.A2(n_1517),
.B(n_1533),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1413),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1444),
.B(n_1513),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1513),
.A2(n_1535),
.B1(n_1430),
.B2(n_1450),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1452),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1489),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1414),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1464),
.A2(n_1415),
.B(n_1412),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1458),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1452),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1443),
.B(n_1455),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1488),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1477),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1510),
.A2(n_1427),
.B(n_1474),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1488),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1458),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1439),
.A2(n_1534),
.B(n_1540),
.Y(n_1634)
);

BUFx2_ASAP7_75t_SL g1635 ( 
.A(n_1467),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1467),
.B(n_1508),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1467),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1530),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1530),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1473),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1469),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1459),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1572),
.B(n_1526),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_SL g1644 ( 
.A1(n_1577),
.A2(n_1504),
.B(n_1431),
.C(n_1537),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1475),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1616),
.A2(n_1523),
.B(n_1516),
.C(n_1419),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1616),
.A2(n_1531),
.B(n_1538),
.C(n_1470),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1564),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1570),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1548),
.B(n_1505),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1618),
.A2(n_1620),
.B(n_1619),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1548),
.B(n_1525),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.B(n_1583),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1557),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1551),
.A2(n_1480),
.B1(n_1459),
.B2(n_1439),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1613),
.A2(n_1422),
.B1(n_1522),
.B2(n_1511),
.C(n_1521),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1618),
.A2(n_1575),
.B(n_1546),
.Y(n_1657)
);

BUFx4f_ASAP7_75t_L g1658 ( 
.A(n_1602),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1525),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1585),
.A2(n_1512),
.B1(n_1524),
.B2(n_1534),
.Y(n_1660)
);

NAND2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1551),
.B(n_1541),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1556),
.A2(n_1512),
.B1(n_1524),
.B2(n_1534),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1585),
.A2(n_1598),
.B1(n_1551),
.B2(n_1595),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1598),
.A2(n_1615),
.B(n_1622),
.C(n_1627),
.Y(n_1665)
);

AO32x2_ASAP7_75t_L g1666 ( 
.A1(n_1543),
.A2(n_1551),
.A3(n_1617),
.B1(n_1642),
.B2(n_1591),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1605),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1565),
.B(n_1544),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1561),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1610),
.A2(n_1612),
.B1(n_1621),
.B2(n_1615),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1573),
.B(n_1636),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1565),
.B(n_1544),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1623),
.B(n_1571),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1599),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1590),
.A2(n_1594),
.B(n_1611),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1622),
.A2(n_1627),
.B1(n_1610),
.B2(n_1612),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1625),
.A2(n_1629),
.B(n_1632),
.C(n_1606),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1576),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1599),
.B(n_1630),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1630),
.B(n_1637),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1623),
.A2(n_1608),
.B1(n_1609),
.B2(n_1594),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1597),
.A2(n_1607),
.B(n_1589),
.C(n_1567),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1623),
.A2(n_1567),
.B1(n_1589),
.B2(n_1586),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1579),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1637),
.B(n_1640),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1555),
.A2(n_1590),
.B(n_1606),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1578),
.B(n_1580),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1608),
.A2(n_1609),
.B1(n_1604),
.B2(n_1607),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1555),
.A2(n_1597),
.B(n_1625),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1559),
.B(n_1568),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1629),
.A2(n_1632),
.B(n_1600),
.C(n_1567),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1589),
.A2(n_1588),
.B(n_1586),
.C(n_1603),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1601),
.B(n_1581),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_SL g1695 ( 
.A1(n_1631),
.A2(n_1642),
.B(n_1617),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1544),
.B(n_1634),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1624),
.B(n_1626),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1588),
.A2(n_1603),
.B(n_1641),
.C(n_1562),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1571),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1569),
.A2(n_1553),
.B(n_1566),
.Y(n_1700)
);

AO32x1_ASAP7_75t_L g1701 ( 
.A1(n_1591),
.A2(n_1593),
.A3(n_1641),
.B1(n_1552),
.B2(n_1560),
.Y(n_1701)
);

AO21x1_ASAP7_75t_L g1702 ( 
.A1(n_1633),
.A2(n_1639),
.B(n_1638),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1571),
.B(n_1582),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1689),
.A2(n_1562),
.B1(n_1604),
.B2(n_1545),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1700),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1547),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1700),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1670),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1648),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1649),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1668),
.B(n_1596),
.Y(n_1711)
);

AOI222xp33_ASAP7_75t_L g1712 ( 
.A1(n_1671),
.A2(n_1544),
.B1(n_1587),
.B2(n_1582),
.C1(n_1628),
.C2(n_1563),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1695),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1691),
.B(n_1558),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1657),
.B(n_1651),
.C(n_1690),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1667),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1666),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1657),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1688),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1687),
.B(n_1547),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1694),
.B(n_1558),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1687),
.B(n_1547),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1653),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1679),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1651),
.B(n_1584),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1685),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1666),
.B(n_1547),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1696),
.B(n_1554),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1584),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1702),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1680),
.Y(n_1731)
);

NOR2xp67_ASAP7_75t_SL g1732 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1675),
.B(n_1681),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1699),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1701),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1701),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1682),
.B(n_1542),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1726),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1715),
.B(n_1674),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1545),
.B1(n_1604),
.B2(n_1682),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1706),
.B(n_1663),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1713),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1715),
.B(n_1669),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1718),
.B(n_1659),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1734),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1717),
.A2(n_1646),
.B(n_1663),
.C(n_1647),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1712),
.A2(n_1665),
.B1(n_1677),
.B2(n_1671),
.C(n_1678),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1726),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1718),
.B(n_1686),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1645),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1730),
.B(n_1631),
.C(n_1677),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1730),
.A2(n_1644),
.B(n_1655),
.C(n_1684),
.Y(n_1754)
);

AO21x2_ASAP7_75t_L g1755 ( 
.A1(n_1707),
.A2(n_1698),
.B(n_1692),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1709),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1709),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1729),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1731),
.B(n_1650),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1734),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1719),
.B(n_1697),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1725),
.B(n_1724),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1731),
.B(n_1652),
.Y(n_1763)
);

AOI33xp33_ASAP7_75t_L g1764 ( 
.A1(n_1727),
.A2(n_1656),
.A3(n_1643),
.B1(n_1683),
.B2(n_1660),
.B3(n_1639),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1724),
.Y(n_1765)
);

AOI222xp33_ASAP7_75t_L g1766 ( 
.A1(n_1720),
.A2(n_1693),
.B1(n_1661),
.B2(n_1669),
.C1(n_1673),
.C2(n_1563),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1707),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1602),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1713),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1738),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1710),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1733),
.B(n_1703),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1712),
.A2(n_1662),
.B1(n_1604),
.B2(n_1631),
.C(n_1655),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1733),
.B(n_1643),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1710),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1708),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1739),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1750),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1750),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_R g1781 ( 
.A(n_1768),
.B(n_1654),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1756),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1745),
.B(n_1735),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1745),
.B(n_1736),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1762),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1767),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1747),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1758),
.B(n_1708),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1744),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1758),
.B(n_1710),
.Y(n_1791)
);

NAND2x1_ASAP7_75t_L g1792 ( 
.A(n_1765),
.B(n_1732),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1756),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1745),
.B(n_1736),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1757),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1745),
.B(n_1737),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1744),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1757),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1767),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1745),
.B(n_1752),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1752),
.B(n_1737),
.Y(n_1801)
);

OR2x6_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1673),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1711),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1743),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1751),
.B(n_1711),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1770),
.B(n_1721),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1766),
.B(n_1728),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1769),
.B(n_1723),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1769),
.B(n_1723),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1781),
.B(n_1792),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1800),
.B(n_1746),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1800),
.B(n_1746),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1777),
.B(n_1770),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1800),
.B(n_1772),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1777),
.B(n_1770),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1790),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1779),
.Y(n_1819)
);

AO22x1_ASAP7_75t_L g1820 ( 
.A1(n_1788),
.A2(n_1720),
.B1(n_1722),
.B2(n_1754),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1803),
.B(n_1772),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1803),
.B(n_1747),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1803),
.B(n_1760),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1797),
.B(n_1765),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1780),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1779),
.B(n_1762),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1808),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1807),
.B(n_1801),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1807),
.B(n_1760),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1792),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1808),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1782),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1788),
.B(n_1771),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1740),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1807),
.B(n_1774),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1801),
.B(n_1774),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1782),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1786),
.B(n_1771),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1793),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1793),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1801),
.B(n_1759),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1786),
.B(n_1775),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1806),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1795),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1810),
.B(n_1759),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1795),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1798),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1810),
.B(n_1811),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1806),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1810),
.B(n_1763),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1804),
.B(n_1761),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1811),
.B(n_1763),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1804),
.B(n_1775),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1806),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1809),
.A2(n_1753),
.B(n_1764),
.C(n_1748),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1778),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1798),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1805),
.B(n_1761),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1834),
.B(n_1811),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1819),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1855),
.A2(n_1754),
.B(n_1748),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1825),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1805),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1851),
.B(n_1789),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1848),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1818),
.B(n_1790),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_1783),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1812),
.B(n_1790),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1821),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1843),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1848),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1818),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1820),
.B(n_1789),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1843),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1819),
.Y(n_1875)
);

INVx2_ASAP7_75t_SL g1876 ( 
.A(n_1822),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1832),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1832),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1821),
.B(n_1783),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1837),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1851),
.B(n_1776),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1837),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1820),
.B(n_1776),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1836),
.B(n_1783),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1836),
.B(n_1784),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1827),
.A2(n_1802),
.B1(n_1773),
.B2(n_1749),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1839),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1816),
.B(n_1574),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1822),
.B(n_1784),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1823),
.B(n_1784),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1835),
.B(n_1794),
.Y(n_1891)
);

INVxp67_ASAP7_75t_SL g1892 ( 
.A(n_1824),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1835),
.B(n_1794),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1816),
.B(n_1794),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1839),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1861),
.B(n_1658),
.Y(n_1896)
);

OAI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1861),
.A2(n_1802),
.B1(n_1749),
.B2(n_1741),
.C(n_1773),
.Y(n_1897)
);

OAI32xp33_ASAP7_75t_L g1898 ( 
.A1(n_1873),
.A2(n_1858),
.A3(n_1827),
.B1(n_1831),
.B2(n_1830),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1894),
.Y(n_1899)
);

AND2x2_ASAP7_75t_SL g1900 ( 
.A(n_1886),
.B(n_1658),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1865),
.B(n_1841),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1860),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1894),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1873),
.A2(n_1802),
.B1(n_1722),
.B2(n_1720),
.Y(n_1904)
);

INVxp67_ASAP7_75t_SL g1905 ( 
.A(n_1868),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1860),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1865),
.B(n_1858),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1869),
.B(n_1845),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1869),
.B(n_1845),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1867),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1866),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1862),
.B(n_1830),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1876),
.B(n_1813),
.Y(n_1913)
);

NOR2x1_ASAP7_75t_L g1914 ( 
.A(n_1862),
.B(n_1824),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1879),
.B(n_1850),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1879),
.B(n_1850),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1881),
.B(n_1831),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1875),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1883),
.B(n_1830),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1871),
.B(n_1841),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1883),
.A2(n_1802),
.B1(n_1722),
.B2(n_1755),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1876),
.B(n_1823),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1872),
.Y(n_1923)
);

A2O1A1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1897),
.A2(n_1859),
.B(n_1889),
.C(n_1890),
.Y(n_1924)
);

AOI322xp5_ASAP7_75t_L g1925 ( 
.A1(n_1900),
.A2(n_1863),
.A3(n_1867),
.B1(n_1884),
.B2(n_1885),
.C1(n_1893),
.C2(n_1891),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1907),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1907),
.B(n_1863),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1896),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1912),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1902),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1906),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1921),
.A2(n_1802),
.B1(n_1892),
.B2(n_1874),
.C(n_1870),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1919),
.A2(n_1802),
.B(n_1888),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1912),
.A2(n_1898),
.B(n_1919),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1900),
.A2(n_1870),
.B1(n_1874),
.B2(n_1755),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1923),
.B(n_1864),
.Y(n_1936)
);

AOI322xp5_ASAP7_75t_L g1937 ( 
.A1(n_1923),
.A2(n_1884),
.A3(n_1885),
.B1(n_1893),
.B2(n_1891),
.C1(n_1874),
.C2(n_1870),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1905),
.A2(n_1833),
.B(n_1875),
.Y(n_1938)
);

AOI31xp33_ASAP7_75t_L g1939 ( 
.A1(n_1911),
.A2(n_1864),
.A3(n_1881),
.B(n_1882),
.Y(n_1939)
);

XNOR2xp5_ASAP7_75t_L g1940 ( 
.A(n_1913),
.B(n_1829),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1922),
.B(n_1829),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1913),
.B(n_1914),
.Y(n_1942)
);

NOR2x1_ASAP7_75t_L g1943 ( 
.A(n_1918),
.B(n_1877),
.Y(n_1943)
);

O2A1O1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1934),
.A2(n_1917),
.B(n_1903),
.C(n_1899),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1939),
.B(n_1908),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1943),
.Y(n_1946)
);

OAI21xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1937),
.A2(n_1909),
.B(n_1908),
.Y(n_1947)
);

AOI222xp33_ASAP7_75t_L g1948 ( 
.A1(n_1926),
.A2(n_1882),
.B1(n_1887),
.B2(n_1895),
.C1(n_1880),
.C2(n_1878),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1927),
.Y(n_1949)
);

NAND2x1_ASAP7_75t_L g1950 ( 
.A(n_1929),
.B(n_1913),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1940),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1927),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1936),
.B(n_1899),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1941),
.B(n_1909),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1930),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1954),
.B(n_1915),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1953),
.B(n_1915),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1945),
.A2(n_1935),
.B1(n_1928),
.B2(n_1932),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1945),
.B(n_1925),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1955),
.Y(n_1960)
);

AOI222xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1946),
.A2(n_1931),
.B1(n_1903),
.B2(n_1910),
.C1(n_1942),
.C2(n_1938),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1949),
.A2(n_1952),
.B1(n_1951),
.B2(n_1933),
.Y(n_1962)
);

NOR2x1p5_ASAP7_75t_L g1963 ( 
.A(n_1950),
.B(n_1910),
.Y(n_1963)
);

NOR3x1_ASAP7_75t_L g1964 ( 
.A(n_1944),
.B(n_1901),
.C(n_1920),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1948),
.A2(n_1904),
.B1(n_1849),
.B2(n_1843),
.Y(n_1965)
);

NOR3xp33_ASAP7_75t_L g1966 ( 
.A(n_1947),
.B(n_1924),
.C(n_1917),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1957),
.B(n_1948),
.Y(n_1967)
);

AOI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1966),
.A2(n_1877),
.B1(n_1895),
.B2(n_1887),
.C(n_1880),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1966),
.A2(n_1916),
.B(n_1878),
.Y(n_1969)
);

OAI222xp33_ASAP7_75t_L g1970 ( 
.A1(n_1959),
.A2(n_1916),
.B1(n_1854),
.B2(n_1849),
.C1(n_1856),
.C2(n_1796),
.Y(n_1970)
);

O2A1O1Ixp5_ASAP7_75t_L g1971 ( 
.A1(n_1956),
.A2(n_1856),
.B(n_1833),
.C(n_1857),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1965),
.A2(n_1854),
.B1(n_1849),
.B2(n_1856),
.C(n_1796),
.Y(n_1972)
);

OA22x2_ASAP7_75t_L g1973 ( 
.A1(n_1969),
.A2(n_1958),
.B1(n_1960),
.B2(n_1961),
.Y(n_1973)
);

AOI211xp5_ASAP7_75t_L g1974 ( 
.A1(n_1967),
.A2(n_1964),
.B(n_1962),
.C(n_1963),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1971),
.Y(n_1975)
);

AOI211xp5_ASAP7_75t_L g1976 ( 
.A1(n_1970),
.A2(n_1796),
.B(n_1857),
.C(n_1844),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1972),
.Y(n_1977)
);

AOI211xp5_ASAP7_75t_L g1978 ( 
.A1(n_1968),
.A2(n_1840),
.B(n_1844),
.C(n_1846),
.Y(n_1978)
);

AOI211xp5_ASAP7_75t_L g1979 ( 
.A1(n_1967),
.A2(n_1840),
.B(n_1847),
.C(n_1846),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1973),
.A2(n_1817),
.B(n_1815),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1977),
.A2(n_1854),
.B1(n_1815),
.B2(n_1817),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1975),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1979),
.Y(n_1983)
);

NOR2xp67_ASAP7_75t_L g1984 ( 
.A(n_1974),
.B(n_1847),
.Y(n_1984)
);

NAND4xp75_ASAP7_75t_L g1985 ( 
.A(n_1976),
.B(n_1813),
.C(n_1814),
.D(n_1852),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1984),
.B(n_1852),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1983),
.B(n_1838),
.Y(n_1987)
);

AO22x2_ASAP7_75t_L g1988 ( 
.A1(n_1982),
.A2(n_1978),
.B1(n_1814),
.B2(n_1842),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1986),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1989),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1990),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1990),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_SL g1993 ( 
.A1(n_1991),
.A2(n_1987),
.B1(n_1980),
.B2(n_1988),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1992),
.A2(n_1985),
.B1(n_1981),
.B2(n_1826),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1993),
.B(n_1838),
.Y(n_1995)
);

OA22x2_ASAP7_75t_L g1996 ( 
.A1(n_1994),
.A2(n_1842),
.B1(n_1826),
.B2(n_1778),
.Y(n_1996)
);

OR2x6_ASAP7_75t_L g1997 ( 
.A(n_1995),
.B(n_1635),
.Y(n_1997)
);

OAI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1996),
.A2(n_1778),
.B1(n_1785),
.B2(n_1787),
.C(n_1799),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1853),
.B(n_1791),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1999),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1998),
.B1(n_1785),
.B2(n_1799),
.Y(n_2001)
);

AOI211xp5_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_1853),
.B(n_1785),
.C(n_1787),
.Y(n_2002)
);


endmodule