module fake_jpeg_18568_n_285 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_57),
.B1(n_59),
.B2(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_43),
.B1(n_34),
.B2(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_34),
.B1(n_17),
.B2(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_48),
.B1(n_57),
.B2(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_106)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_65),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_44),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_68),
.A2(n_69),
.B1(n_0),
.B2(n_2),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_40),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_79),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_36),
.B1(n_52),
.B2(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_91),
.B1(n_32),
.B2(n_25),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_92),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_21),
.B1(n_35),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_80),
.B1(n_88),
.B2(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_40),
.B(n_39),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_39),
.B1(n_40),
.B2(n_32),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_25),
.B(n_1),
.C(n_2),
.Y(n_110)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_33),
.B1(n_19),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_30),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_31),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_50),
.B(n_32),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_24),
.A3(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_103),
.B(n_87),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_110),
.B1(n_68),
.B2(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_120),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_73),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_10),
.C(n_15),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_85),
.C(n_83),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_96),
.B1(n_65),
.B2(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_141),
.B1(n_142),
.B2(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_135),
.B1(n_99),
.B2(n_110),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_64),
.B1(n_102),
.B2(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_144),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_107),
.B1(n_120),
.B2(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_85),
.B1(n_68),
.B2(n_75),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_69),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_122),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_98),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_146),
.C(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_66),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_66),
.B(n_70),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_76),
.C(n_4),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_150),
.C(n_112),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_10),
.C(n_4),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_11),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_11),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_99),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_106),
.B1(n_124),
.B2(n_122),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_155),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_126),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_171),
.B(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_149),
.B1(n_150),
.B2(n_113),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_166),
.B1(n_176),
.B2(n_142),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_178),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_103),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_106),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_110),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_131),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_113),
.B1(n_111),
.B2(n_100),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_143),
.CI(n_128),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_186),
.A2(n_203),
.B1(n_161),
.B2(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_143),
.C(n_128),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_200),
.C(n_206),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_152),
.B(n_133),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_173),
.B(n_171),
.C(n_181),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_152),
.B(n_135),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_207),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_145),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_139),
.B1(n_151),
.B2(n_154),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_205),
.B1(n_156),
.B2(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_111),
.B1(n_100),
.B2(n_114),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_114),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_12),
.C(n_5),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_212),
.B1(n_197),
.B2(n_169),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_207),
.B(n_191),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_213),
.B1(n_225),
.B2(n_226),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_182),
.B1(n_165),
.B2(n_167),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_182),
.B1(n_164),
.B2(n_177),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_177),
.C(n_162),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_200),
.C(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_116),
.C(n_7),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_205),
.B1(n_204),
.B2(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_198),
.B1(n_192),
.B2(n_199),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_184),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_210),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_185),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_191),
.B1(n_184),
.B2(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_210),
.C(n_217),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_215),
.C(n_221),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_210),
.C(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_242),
.C(n_231),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

OAI211xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_243),
.B(n_235),
.C(n_239),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_227),
.B(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_264),
.C(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_233),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_251),
.B1(n_252),
.B2(n_256),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_264),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_249),
.B(n_237),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_251),
.C(n_230),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_275),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_276),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_245),
.B(n_248),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_236),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_266),
.B(n_267),
.C(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_259),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_281),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_13),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_8),
.B(n_9),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_9),
.B(n_12),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_14),
.Y(n_285)
);


endmodule