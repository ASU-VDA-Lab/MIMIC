module fake_jpeg_1455_n_463 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_463);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_463;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_52),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_1),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_65),
.A2(n_23),
.B(n_6),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_17),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_78),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_37),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_81),
.B(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_3),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_75),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_39),
.B1(n_30),
.B2(n_24),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_86),
.A2(n_87),
.B1(n_99),
.B2(n_108),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_30),
.B1(n_20),
.B2(n_24),
.Y(n_87)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_45),
.B1(n_34),
.B2(n_25),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_23),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_45),
.B1(n_17),
.B2(n_33),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_97),
.A2(n_107),
.B1(n_125),
.B2(n_126),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_30),
.B1(n_24),
.B2(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_32),
.B1(n_41),
.B2(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_24),
.B1(n_41),
.B2(n_40),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_118),
.A2(n_119),
.B1(n_129),
.B2(n_36),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_156)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_31),
.CON(n_123),
.SN(n_123)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_144),
.B(n_107),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_46),
.A2(n_42),
.B1(n_36),
.B2(n_14),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_51),
.A2(n_76),
.B1(n_66),
.B2(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_48),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_4),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_31),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_62),
.B(n_74),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_42),
.B1(n_36),
.B2(n_31),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_31),
.B1(n_23),
.B2(n_42),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_31),
.B1(n_23),
.B2(n_42),
.Y(n_135)
);

INVx5_ASAP7_75t_SL g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g183 ( 
.A(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_14),
.Y(n_148)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

OR2x4_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_42),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_171),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_14),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_153),
.B(n_169),
.Y(n_247)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_188),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_93),
.B(n_13),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_105),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_177),
.Y(n_211)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_112),
.B(n_15),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_180),
.Y(n_215)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_116),
.B(n_11),
.Y(n_180)
);

BUFx24_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_16),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_184),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_4),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_139),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_6),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_193),
.Y(n_239)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_196),
.Y(n_236)
);

NAND2x1p5_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_170),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_113),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_195),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_138),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_110),
.B1(n_102),
.B2(n_89),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_8),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_200),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_208),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_157),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_123),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_229),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_94),
.B(n_120),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_210),
.B(n_183),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_163),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_139),
.B1(n_113),
.B2(n_121),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_217),
.A2(n_205),
.B1(n_248),
.B2(n_243),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_136),
.B1(n_133),
.B2(n_89),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_151),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_150),
.B(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_221),
.B(n_225),
.Y(n_290)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_90),
.B1(n_92),
.B2(n_96),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_171),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_245),
.B1(n_183),
.B2(n_145),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_154),
.B(n_91),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_146),
.B(n_138),
.C(n_102),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_243),
.C(n_191),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_156),
.A2(n_90),
.B(n_103),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_155),
.B(n_198),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_36),
.C(n_110),
.Y(n_243)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_36),
.B1(n_35),
.B2(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_213),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_274),
.C(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_255),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_197),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_257),
.A2(n_266),
.B(n_234),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_259),
.A2(n_270),
.B1(n_276),
.B2(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_269),
.B(n_237),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_158),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_196),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_263),
.B(n_273),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_165),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_271),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_216),
.A2(n_158),
.B1(n_157),
.B2(n_147),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_216),
.A2(n_164),
.B1(n_152),
.B2(n_166),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_172),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_179),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_176),
.B1(n_174),
.B2(n_168),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_216),
.A2(n_214),
.B1(n_230),
.B2(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_279),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_211),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_235),
.B(n_215),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_280),
.B(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_172),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_167),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_247),
.B(n_159),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_221),
.A2(n_160),
.B1(n_167),
.B2(n_151),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_28),
.B1(n_9),
.B2(n_10),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_210),
.A2(n_28),
.B1(n_9),
.B2(n_10),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_8),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_236),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_208),
.B(n_9),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_222),
.C(n_244),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_284),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_295),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_297),
.A2(n_307),
.B(n_318),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_260),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_308),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_209),
.B(n_229),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_310),
.B(n_322),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_261),
.A2(n_204),
.B(n_242),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_220),
.B(n_204),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_251),
.B(n_204),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_326),
.C(n_269),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_220),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_313),
.B(n_317),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_233),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_327),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_276),
.B(n_248),
.CI(n_238),
.CON(n_317),
.SN(n_317)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_277),
.A2(n_237),
.B(n_238),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_319),
.A2(n_320),
.B(n_324),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_233),
.B(n_207),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_264),
.A2(n_207),
.B(n_212),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_228),
.B1(n_223),
.B2(n_246),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_259),
.B1(n_275),
.B2(n_264),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_277),
.A2(n_212),
.B(n_246),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_228),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_325),
.B(n_330),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_219),
.C(n_223),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_219),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_10),
.C(n_28),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_274),
.B1(n_288),
.B2(n_254),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_332),
.A2(n_335),
.B1(n_343),
.B2(n_344),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_287),
.B(n_268),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_318),
.B(n_297),
.Y(n_386)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_341),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_255),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_349),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_294),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_296),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_347),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_252),
.B1(n_271),
.B2(n_273),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_299),
.A2(n_305),
.B1(n_327),
.B2(n_303),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_316),
.A2(n_289),
.B1(n_292),
.B2(n_291),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_348),
.A2(n_351),
.B1(n_304),
.B2(n_302),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_299),
.A2(n_270),
.B1(n_250),
.B2(n_256),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_350),
.A2(n_345),
.B1(n_338),
.B2(n_344),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_323),
.A2(n_285),
.B1(n_258),
.B2(n_267),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_356),
.C(n_308),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_272),
.C(n_278),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_296),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_357),
.B(n_360),
.Y(n_366)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_293),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_307),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_300),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_377),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_368),
.A2(n_369),
.B1(n_388),
.B2(n_353),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_331),
.B1(n_302),
.B2(n_312),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_345),
.B(n_331),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_370),
.B(n_379),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_361),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_384),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_383),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_304),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_378),
.A2(n_353),
.B1(n_348),
.B2(n_351),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_333),
.A2(n_318),
.B(n_321),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_312),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_385),
.C(n_328),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_326),
.Y(n_385)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_386),
.A2(n_352),
.B(n_253),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_334),
.B(n_314),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_387),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_314),
.B1(n_317),
.B2(n_320),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_317),
.C(n_329),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_349),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_346),
.B(n_355),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_392),
.A2(n_396),
.B(n_398),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_332),
.B1(n_346),
.B2(n_350),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_393),
.A2(n_378),
.B1(n_376),
.B2(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_384),
.B(n_355),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_397),
.A2(n_380),
.B1(n_389),
.B2(n_382),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_339),
.B(n_347),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_402),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_408),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_377),
.B(n_358),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_336),
.B(n_333),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_405),
.B(n_407),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_365),
.A2(n_322),
.B(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_409),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_328),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_413),
.A2(n_397),
.B1(n_404),
.B2(n_392),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_383),
.C(n_372),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_419),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_405),
.B1(n_409),
.B2(n_410),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_408),
.C(n_390),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_367),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_421),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_372),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_381),
.C(n_375),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_394),
.C(n_393),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_366),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_407),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_295),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_406),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_404),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_431),
.A2(n_435),
.B1(n_440),
.B2(n_414),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_437),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_395),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_434),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_438),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_380),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_425),
.A2(n_253),
.B(n_329),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_411),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_411),
.B(n_422),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_413),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_445),
.B1(n_446),
.B2(n_449),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_420),
.C(n_419),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_427),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_448),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_418),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_447),
.A2(n_434),
.B1(n_415),
.B2(n_424),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_452),
.A2(n_453),
.B(n_455),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_417),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_437),
.Y(n_455)
);

AOI322xp5_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_455),
.A3(n_454),
.B1(n_441),
.B2(n_444),
.C1(n_451),
.C2(n_436),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_456),
.B(n_417),
.Y(n_459)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_450),
.A2(n_441),
.B(n_416),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_458),
.B(n_457),
.C(n_430),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_460),
.C(n_430),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_421),
.B(n_286),
.Y(n_463)
);


endmodule