module fake_jpeg_12677_n_663 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_663);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_663;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_9),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_62),
.B(n_110),
.Y(n_216)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_66),
.Y(n_223)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_68),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_75),
.A2(n_88),
.B1(n_45),
.B2(n_23),
.Y(n_188)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_78),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_83),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_18),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_89),
.Y(n_225)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_91),
.B(n_43),
.Y(n_145)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_42),
.B(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_118),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_20),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_58),
.Y(n_142)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_32),
.Y(n_130)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_40),
.Y(n_131)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

AND2x4_ASAP7_75t_SL g132 ( 
.A(n_62),
.B(n_45),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_132),
.B(n_15),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_50),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_140),
.B(n_143),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_142),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_47),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_145),
.B(n_158),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_56),
.B1(n_25),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_147),
.A2(n_160),
.B1(n_183),
.B2(n_195),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_SL g153 ( 
.A(n_67),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_153),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_50),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_61),
.A2(n_25),
.B1(n_44),
.B2(n_33),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_56),
.B1(n_25),
.B2(n_27),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_161),
.A2(n_177),
.B1(n_201),
.B2(n_32),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_54),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_166),
.B(n_167),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_43),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_65),
.A2(n_20),
.B1(n_27),
.B2(n_44),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_54),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_179),
.B(n_200),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_115),
.B(n_52),
.C(n_47),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_88),
.C(n_110),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_68),
.A2(n_81),
.B1(n_78),
.B2(n_66),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_188),
.A2(n_209),
.B1(n_219),
.B2(n_109),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_86),
.A2(n_53),
.B1(n_52),
.B2(n_44),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_198),
.B(n_35),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_64),
.B(n_53),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_69),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_77),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_204),
.B(n_221),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_77),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_222),
.B1(n_108),
.B2(n_120),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_99),
.A2(n_33),
.B1(n_28),
.B2(n_23),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_76),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_103),
.A2(n_28),
.B1(n_41),
.B2(n_13),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_104),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_93),
.B(n_35),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_106),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_227),
.Y(n_319)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_229),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_230),
.B(n_246),
.Y(n_348)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_234),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_235),
.Y(n_339)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_147),
.A2(n_72),
.B1(n_79),
.B2(n_117),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_237),
.A2(n_284),
.B1(n_292),
.B2(n_307),
.Y(n_311)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_238),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_239),
.B(n_264),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_148),
.B(n_0),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_240),
.B(n_248),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_243),
.Y(n_345)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_212),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_132),
.B(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_250),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_162),
.C(n_155),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_251),
.B(n_298),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_254),
.A2(n_164),
.B1(n_175),
.B2(n_157),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_212),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_256),
.B(n_263),
.Y(n_351)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_137),
.Y(n_258)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_259),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_260),
.A2(n_299),
.B(n_305),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_261),
.B(n_271),
.Y(n_346)
);

INVx4_ASAP7_75t_SL g263 ( 
.A(n_153),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_208),
.A2(n_123),
.B1(n_118),
.B2(n_93),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_267),
.A2(n_290),
.B1(n_294),
.B2(n_303),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_216),
.A2(n_118),
.B(n_109),
.C(n_35),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_268),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_248),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_139),
.B(n_1),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_150),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_274),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_165),
.B(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_276),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_138),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_201),
.A2(n_89),
.B1(n_96),
.B2(n_116),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_280),
.A2(n_285),
.B1(n_289),
.B2(n_297),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_281),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_357)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_282),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_163),
.B(n_32),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_283),
.B(n_295),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_160),
.A2(n_32),
.B1(n_39),
.B2(n_41),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_161),
.A2(n_41),
.B1(n_39),
.B2(n_12),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_172),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_296),
.Y(n_329)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_149),
.Y(n_287)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_177),
.Y(n_288)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_41),
.B1(n_39),
.B2(n_12),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_190),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_183),
.A2(n_39),
.B1(n_41),
.B2(n_3),
.Y(n_292)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_169),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_199),
.B(n_10),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_222),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_224),
.A2(n_39),
.B1(n_10),
.B2(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_151),
.B(n_18),
.C(n_16),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_186),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_304),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_171),
.B(n_15),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_301),
.B(n_2),
.Y(n_355)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_175),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_192),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_144),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_146),
.B(n_1),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_157),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_238),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_205),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_180),
.B1(n_211),
.B2(n_154),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_308),
.A2(n_333),
.B1(n_337),
.B2(n_340),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_214),
.B1(n_191),
.B2(n_189),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_284),
.A2(n_189),
.B1(n_197),
.B2(n_213),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_318),
.A2(n_323),
.B1(n_354),
.B2(n_256),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_241),
.A2(n_144),
.B1(n_213),
.B2(n_164),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_324),
.B(n_233),
.Y(n_406)
);

NAND2x1_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_159),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_328),
.A2(n_359),
.B(n_355),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_260),
.A2(n_180),
.B1(n_211),
.B2(n_154),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_281),
.A2(n_192),
.B1(n_193),
.B2(n_133),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_338),
.B(n_5),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_230),
.A2(n_193),
.B1(n_133),
.B2(n_152),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_228),
.A2(n_225),
.B1(n_152),
.B2(n_207),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_353),
.B1(n_357),
.B2(n_229),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_358),
.B1(n_252),
.B2(n_234),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_237),
.A2(n_225),
.B1(n_159),
.B2(n_170),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_294),
.A2(n_202),
.B1(n_206),
.B2(n_185),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_239),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_293),
.A2(n_3),
.B(n_4),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_261),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_276),
.Y(n_371)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_366),
.A2(n_299),
.B(n_305),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_369),
.B(n_396),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_371),
.B(n_380),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_251),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_378),
.C(n_381),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_373),
.A2(n_379),
.B1(n_387),
.B2(n_389),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_240),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_377),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_338),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_291),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_367),
.A2(n_271),
.B1(n_257),
.B2(n_247),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_255),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_250),
.C(n_299),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_384),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_385),
.A2(n_386),
.B1(n_402),
.B2(n_411),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_367),
.A2(n_350),
.B1(n_337),
.B2(n_308),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_311),
.A2(n_266),
.B1(n_298),
.B2(n_265),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_335),
.B(n_262),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_390),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_273),
.B1(n_290),
.B2(n_253),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_249),
.C(n_245),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_302),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_392),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_326),
.Y(n_392)
);

BUFx24_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_325),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_398),
.Y(n_438)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_332),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_329),
.A2(n_272),
.B(n_258),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_399),
.A2(n_405),
.B(n_412),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_270),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_400),
.B(n_416),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_344),
.B(n_328),
.C(n_340),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_351),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_333),
.A2(n_232),
.B1(n_244),
.B2(n_231),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_325),
.B(n_287),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_408),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_329),
.A2(n_282),
.B(n_246),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_406),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_407),
.A2(n_415),
.B(n_358),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_306),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_320),
.B(n_304),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_413),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_353),
.A2(n_242),
.B1(n_303),
.B2(n_235),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_328),
.A2(n_269),
.B(n_236),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_320),
.B(n_5),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_349),
.A2(n_6),
.B1(n_263),
.B2(n_314),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_414),
.A2(n_347),
.B1(n_343),
.B2(n_332),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_314),
.A2(n_352),
.B1(n_324),
.B2(n_347),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_322),
.B(n_359),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_408),
.A2(n_312),
.B1(n_322),
.B2(n_364),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_420),
.A2(n_427),
.B1(n_431),
.B2(n_406),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_401),
.A2(n_407),
.B(n_416),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_426),
.A2(n_430),
.B(n_440),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_324),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_429),
.B(n_445),
.C(n_396),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_412),
.A2(n_324),
.B(n_343),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_376),
.A2(n_415),
.B1(n_386),
.B2(n_414),
.Y(n_431)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_382),
.Y(n_436)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_436),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_370),
.A2(n_317),
.B(n_351),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_387),
.A2(n_309),
.B1(n_360),
.B2(n_321),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_442),
.A2(n_451),
.B1(n_453),
.B2(n_455),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_351),
.B(n_342),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_444),
.A2(n_406),
.B(n_410),
.Y(n_463)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_446),
.Y(n_482)
);

FAx1_ASAP7_75t_SL g449 ( 
.A(n_374),
.B(n_317),
.CI(n_341),
.CON(n_449),
.SN(n_449)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_378),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_389),
.A2(n_360),
.B1(n_321),
.B2(n_356),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_373),
.A2(n_356),
.B1(n_341),
.B2(n_336),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_376),
.A2(n_310),
.B1(n_330),
.B2(n_365),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_371),
.B(n_310),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_383),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_432),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_471),
.C(n_481),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_458),
.A2(n_479),
.B(n_472),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_425),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_459),
.B(n_464),
.Y(n_494)
);

O2A1O1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_394),
.B(n_370),
.C(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_385),
.B1(n_391),
.B2(n_398),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_489),
.B1(n_492),
.B2(n_444),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_466),
.A2(n_470),
.B1(n_472),
.B2(n_488),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_467),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_424),
.B(n_392),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_468),
.B(n_474),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_372),
.B1(n_378),
.B2(n_379),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_372),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_420),
.A2(n_377),
.B1(n_390),
.B2(n_403),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_424),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_413),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_476),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_400),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_447),
.A2(n_384),
.B1(n_381),
.B2(n_405),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_438),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_480),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_369),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_456),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_483),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_455),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_487),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_437),
.B(n_380),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_490),
.C(n_437),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_402),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_486),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_427),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_425),
.A2(n_404),
.B1(n_393),
.B2(n_409),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_428),
.A2(n_443),
.B1(n_452),
.B2(n_448),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_423),
.A2(n_411),
.B1(n_375),
.B2(n_342),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_491),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_423),
.A2(n_342),
.B1(n_317),
.B2(n_362),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_493),
.B(n_421),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_426),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_504),
.Y(n_533)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_498),
.A2(n_499),
.B1(n_515),
.B2(n_520),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_465),
.A2(n_419),
.B1(n_448),
.B2(n_430),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_519),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_474),
.B(n_454),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_526),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_429),
.Y(n_504)
);

AOI22x1_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_462),
.B1(n_486),
.B2(n_487),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_507),
.A2(n_486),
.B1(n_458),
.B2(n_491),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_452),
.C(n_454),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_511),
.C(n_522),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_439),
.C(n_419),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_484),
.A2(n_449),
.B1(n_450),
.B2(n_439),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_450),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_517),
.B(n_473),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_461),
.A2(n_449),
.B1(n_418),
.B2(n_441),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_461),
.A2(n_436),
.B1(n_422),
.B2(n_442),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_521),
.A2(n_528),
.B1(n_425),
.B2(n_330),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_440),
.C(n_422),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_460),
.B(n_417),
.C(n_446),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_482),
.C(n_478),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_468),
.B(n_345),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_475),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_464),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_469),
.A2(n_453),
.B(n_393),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_527),
.B(n_393),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_462),
.A2(n_480),
.B1(n_466),
.B2(n_483),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_467),
.B(n_451),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_529),
.B(n_493),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_476),
.Y(n_530)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

AOI31xp33_ASAP7_75t_L g575 ( 
.A1(n_531),
.A2(n_516),
.A3(n_513),
.B(n_514),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_534),
.A2(n_558),
.B1(n_503),
.B2(n_518),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_523),
.A2(n_460),
.B1(n_463),
.B2(n_473),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_535),
.A2(n_506),
.B1(n_521),
.B2(n_507),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_509),
.A2(n_479),
.B(n_458),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_536),
.B(n_549),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_545),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_539),
.B(n_541),
.C(n_557),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_500),
.B(n_482),
.C(n_478),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_494),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_547),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_435),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_546),
.B(n_555),
.Y(n_569)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_494),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_496),
.B(n_492),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_498),
.Y(n_563)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_501),
.B(n_435),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_551),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_508),
.B(n_362),
.Y(n_551)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_552),
.B(n_540),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_507),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_553),
.B(n_528),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_554),
.A2(n_503),
.B(n_515),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_319),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_459),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_556),
.B(n_559),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_500),
.B(n_363),
.C(n_365),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_504),
.B(n_363),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_313),
.C(n_345),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_560),
.B(n_522),
.C(n_509),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_563),
.B(n_581),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_564),
.A2(n_576),
.B1(n_535),
.B2(n_558),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_567),
.B(n_574),
.Y(n_603)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_568),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_541),
.B(n_499),
.C(n_519),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_570),
.B(n_572),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_529),
.C(n_520),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_575),
.B(n_542),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_537),
.A2(n_506),
.B1(n_512),
.B2(n_513),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_557),
.B(n_532),
.C(n_539),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_580),
.C(n_559),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_537),
.B1(n_552),
.B2(n_545),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_532),
.B(n_556),
.C(n_560),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_533),
.B(n_516),
.Y(n_581)
);

FAx1_ASAP7_75t_SL g582 ( 
.A(n_530),
.B(n_527),
.CI(n_393),
.CON(n_582),
.SN(n_582)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_538),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_316),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_584),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_533),
.B(n_334),
.Y(n_584)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_585),
.Y(n_587)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_586),
.Y(n_613)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_588),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_589),
.A2(n_572),
.B1(n_563),
.B2(n_582),
.Y(n_609)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_585),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_590),
.B(n_595),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g591 ( 
.A1(n_566),
.A2(n_536),
.B(n_544),
.Y(n_591)
);

CKINVDCx14_ASAP7_75t_R g612 ( 
.A(n_591),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_573),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_592),
.B(n_319),
.Y(n_622)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_576),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_564),
.A2(n_562),
.B1(n_570),
.B2(n_567),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_596),
.A2(n_578),
.B1(n_580),
.B2(n_581),
.Y(n_614)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_600),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_548),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_605),
.C(n_561),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_577),
.B(n_313),
.Y(n_619)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_574),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_582),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_544),
.C(n_313),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_619),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g631 ( 
.A(n_609),
.B(n_593),
.Y(n_631)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_610),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_614),
.A2(n_589),
.B1(n_602),
.B2(n_603),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_598),
.B(n_571),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_615),
.B(n_618),
.Y(n_636)
);

BUFx24_ASAP7_75t_SL g616 ( 
.A(n_603),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_616),
.B(n_622),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_595),
.A2(n_565),
.B1(n_584),
.B2(n_583),
.Y(n_617)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_617),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_577),
.C(n_565),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_316),
.C(n_327),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_620),
.B(n_597),
.C(n_593),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_604),
.A2(n_319),
.B(n_334),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_621),
.A2(n_587),
.B(n_590),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_630),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_607),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_625),
.B(n_629),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_606),
.B(n_587),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_627),
.A2(n_619),
.B(n_617),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_618),
.B(n_596),
.C(n_599),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_631),
.B(n_609),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_588),
.C(n_601),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_632),
.B(n_634),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_594),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_606),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_637),
.B(n_624),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_641),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_611),
.C(n_620),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_642),
.B(n_644),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_636),
.A2(n_613),
.B(n_621),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_643),
.A2(n_645),
.B(n_646),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_611),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_597),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_638),
.B(n_624),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_647),
.A2(n_649),
.B(n_640),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_SL g656 ( 
.A1(n_648),
.A2(n_631),
.B(n_623),
.C(n_628),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_642),
.B(n_639),
.C(n_632),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_646),
.A2(n_631),
.B(n_630),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_653),
.A2(n_339),
.B(n_327),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_654),
.B(n_656),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_SL g655 ( 
.A1(n_652),
.A2(n_641),
.B(n_633),
.C(n_627),
.Y(n_655)
);

AOI321xp33_ASAP7_75t_L g658 ( 
.A1(n_655),
.A2(n_657),
.A3(n_651),
.B1(n_650),
.B2(n_649),
.C(n_647),
.Y(n_658)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_658),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_660),
.A2(n_659),
.B(n_339),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_661),
.B(n_339),
.Y(n_662)
);

MAJx2_ASAP7_75t_L g663 ( 
.A(n_662),
.B(n_339),
.C(n_393),
.Y(n_663)
);


endmodule