module fake_jpeg_23339_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_32),
.B1(n_46),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_25),
.B1(n_36),
.B2(n_28),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_38),
.B1(n_20),
.B2(n_19),
.Y(n_112)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_86),
.B1(n_34),
.B2(n_35),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_84),
.B(n_14),
.Y(n_116)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_114),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_18),
.C(n_29),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_34),
.C(n_27),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_95),
.Y(n_148)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_103),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_1),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_106),
.B(n_34),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_1),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_65),
.B(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_58),
.B1(n_56),
.B2(n_26),
.Y(n_140)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_18),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_120),
.Y(n_143)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_57),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_77),
.B(n_14),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_132),
.C(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_88),
.B1(n_109),
.B2(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_136),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_81),
.C(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_100),
.Y(n_162)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_139),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_91),
.A3(n_106),
.B1(n_101),
.B2(n_57),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_90),
.Y(n_172)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_159),
.B1(n_142),
.B2(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_25),
.B1(n_26),
.B2(n_21),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_151),
.B1(n_156),
.B2(n_96),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_25),
.B1(n_26),
.B2(n_21),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_18),
.C(n_27),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_149),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_89),
.A2(n_27),
.B(n_18),
.C(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_27),
.B(n_25),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_99),
.A2(n_109),
.B1(n_120),
.B2(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_27),
.C(n_34),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_104),
.C(n_119),
.Y(n_176)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_7),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_27),
.B1(n_19),
.B2(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_94),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_96),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_193),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_88),
.B1(n_122),
.B2(n_107),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_155),
.B(n_139),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_136),
.B1(n_11),
.B2(n_12),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_169),
.B(n_13),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_3),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_174),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_156),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_179),
.C(n_156),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_128),
.B(n_4),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_186),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_119),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_187),
.B1(n_10),
.B2(n_12),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_184),
.B1(n_150),
.B2(n_155),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_141),
.B1(n_158),
.B2(n_126),
.Y(n_184)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_203),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_217),
.B(n_171),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_125),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_137),
.B1(n_156),
.B2(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_148),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_209),
.C(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_210),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_219),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_223),
.B1(n_162),
.B2(n_163),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_15),
.B(n_16),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_16),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_173),
.A2(n_16),
.B1(n_160),
.B2(n_166),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_173),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_246),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_160),
.CI(n_179),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_203),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_229),
.A2(n_239),
.B(n_245),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_208),
.C(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_197),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_180),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_183),
.B(n_178),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_214),
.B(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_223),
.B1(n_200),
.B2(n_198),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_256),
.B1(n_237),
.B2(n_241),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_267),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_198),
.B1(n_211),
.B2(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_264),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_239),
.B(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_195),
.B1(n_210),
.B2(n_204),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_201),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_230),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_270),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_243),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_235),
.C(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_268),
.C(n_249),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_285),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_276),
.B(n_284),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_228),
.C(n_226),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_224),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_274),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_291),
.C(n_244),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_268),
.B1(n_262),
.B2(n_266),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_257),
.C(n_258),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_252),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_296),
.A2(n_279),
.B1(n_250),
.B2(n_269),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_240),
.B1(n_237),
.B2(n_231),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_216),
.B1(n_248),
.B2(n_246),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_277),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_282),
.B(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_299),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_309),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_301),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_293),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_270),
.C(n_283),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_259),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_295),
.B(n_287),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_297),
.B(n_294),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_289),
.B1(n_292),
.B2(n_307),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_302),
.B(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_320),
.B(n_312),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_310),
.B(n_314),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_325),
.B(n_225),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_316),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_207),
.B(n_238),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_220),
.A3(n_205),
.B1(n_215),
.B2(n_238),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_205),
.Y(n_332)
);


endmodule