module fake_netlist_6_3965_n_2244 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2244);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2244;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_2016;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_119),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_49),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_77),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_28),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_181),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_102),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_197),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_45),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_85),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_65),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_210),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_138),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_207),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_101),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_97),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_8),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_143),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_221),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_146),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_110),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_129),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_18),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_89),
.Y(n_287)
);

BUFx2_ASAP7_75t_R g288 ( 
.A(n_171),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_172),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_64),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_161),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_117),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_193),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_20),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_191),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_92),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_70),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_217),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_95),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_3),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_223),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_23),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_3),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_168),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_31),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_195),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_38),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_12),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_25),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_136),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_72),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_150),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_80),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_127),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_78),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_114),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_201),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_113),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_196),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_46),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_204),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_15),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_214),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_25),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_81),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_225),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_8),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_55),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_125),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_5),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_52),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_224),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_230),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_44),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_75),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_22),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_158),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_54),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_108),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_60),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_51),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_36),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_20),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_87),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_44),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_141),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_105),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_2),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_57),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_84),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_120),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_91),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_104),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_65),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_202),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_206),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_198),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_14),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_94),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_43),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_26),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_215),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_107),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_72),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_151),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_100),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_66),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_43),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_63),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_86),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_220),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_79),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_6),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_45),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_68),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_48),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_76),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_213),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_1),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_64),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_36),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_124),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_14),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_48),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_132),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_226),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_139),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_31),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_216),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_178),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_157),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_47),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_24),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_155),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_148),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_26),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_111),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_200),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_9),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_229),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_67),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_176),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_70),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_30),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_106),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_55),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_49),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_59),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_211),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_109),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_165),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_177),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_58),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_18),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_192),
.Y(n_424)
);

BUFx10_ASAP7_75t_L g425 ( 
.A(n_186),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_68),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_1),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_19),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_53),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_128),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_35),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_6),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_164),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_144),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_147),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_42),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_11),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_17),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_153),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_40),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_69),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_73),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_39),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_21),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_4),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_22),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_67),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_122),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_156),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_189),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_140),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_123),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_154),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_52),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_135),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_187),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_32),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_235),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_336),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_R g461 ( 
.A(n_267),
.B(n_4),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_276),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_300),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_336),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_265),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_336),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_7),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_281),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_336),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_284),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_336),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_336),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_336),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_278),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_285),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_336),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_234),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_280),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_286),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_329),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_234),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_329),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_329),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_291),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_329),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_329),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_298),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_282),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_302),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_287),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_256),
.B(n_7),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_321),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_310),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_315),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_257),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g505 ( 
.A(n_411),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_335),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_316),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_317),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_363),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_319),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_409),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_331),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_414),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_232),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_380),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_418),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_333),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_243),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_251),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_363),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_380),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_337),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_232),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_339),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_363),
.Y(n_526)
);

INVxp33_ASAP7_75t_SL g527 ( 
.A(n_236),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_387),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_256),
.B(n_10),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_345),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_400),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_239),
.B(n_245),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_275),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_254),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_351),
.B(n_11),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_236),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_352),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_363),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_233),
.B(n_246),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_279),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_387),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_354),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_428),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_305),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_351),
.B(n_12),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_357),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_292),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_307),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_240),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_308),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_399),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_313),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_394),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_327),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_340),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_399),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_347),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_240),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_349),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_350),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_373),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_378),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_382),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_358),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_265),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_383),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_392),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_283),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_405),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_415),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_370),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_233),
.B(n_13),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_446),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_289),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_423),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_458),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_516),
.B(n_246),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_466),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_519),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_484),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_484),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_486),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_533),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_541),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_487),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_534),
.B(n_343),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_572),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_579),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_462),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_489),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_476),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_510),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_446),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_521),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_526),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_524),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_538),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_470),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_542),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_470),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_482),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_466),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_505),
.B(n_472),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_472),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_540),
.A2(n_465),
.B(n_460),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_548),
.B(n_531),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_478),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_543),
.B(n_294),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_478),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_466),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_544),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_546),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_467),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_555),
.B(n_305),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_560),
.B(n_294),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_473),
.B(n_238),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_474),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_483),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_475),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_483),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_520),
.B(n_288),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_488),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_481),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_479),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_488),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_491),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_481),
.B(n_305),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_569),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_R g648 ( 
.A(n_491),
.B(n_290),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_569),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_493),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_577),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_569),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_501),
.B(n_238),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_551),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_501),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_493),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_557),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_497),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_497),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_552),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_500),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_492),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_494),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_557),
.Y(n_666)
);

CKINVDCx8_ASAP7_75t_R g667 ( 
.A(n_507),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_581),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_265),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_507),
.Y(n_670)
);

CKINVDCx16_ASAP7_75t_R g671 ( 
.A(n_496),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_508),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_556),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_558),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_588),
.A2(n_502),
.B1(n_461),
.B2(n_469),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_634),
.B(n_273),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_646),
.B(n_508),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_632),
.B(n_511),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_632),
.B(n_511),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_634),
.B(n_604),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_646),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_562),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_642),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_648),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_599),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_622),
.B(n_468),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_635),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_635),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_638),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_618),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_273),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_638),
.B(n_513),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_618),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_643),
.B(n_513),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_634),
.B(n_274),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_640),
.B(n_274),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_643),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_595),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_527),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_631),
.B(n_518),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_631),
.B(n_518),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_669),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_633),
.B(n_523),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_642),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_614),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_611),
.B(n_463),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_587),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_630),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_669),
.B(n_523),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_591),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_592),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_669),
.B(n_265),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_657),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_657),
.B(n_527),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_630),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_634),
.B(n_297),
.Y(n_720)
);

CKINVDCx16_ASAP7_75t_R g721 ( 
.A(n_671),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_669),
.A2(n_529),
.B1(n_535),
.B2(n_495),
.Y(n_722)
);

INVx4_ASAP7_75t_SL g723 ( 
.A(n_669),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_477),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_623),
.B(n_464),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_674),
.B(n_536),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_639),
.B(n_504),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_621),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_654),
.B(n_297),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_656),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_662),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_621),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_654),
.B(n_485),
.Y(n_733)
);

BUFx4f_ASAP7_75t_L g734 ( 
.A(n_654),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_654),
.B(n_334),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_675),
.B(n_334),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_674),
.B(n_536),
.Y(n_737)
);

AND2x6_ASAP7_75t_L g738 ( 
.A(n_659),
.B(n_455),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_675),
.B(n_455),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_667),
.A2(n_459),
.B1(n_553),
.B2(n_530),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_672),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_619),
.B(n_525),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_674),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_616),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_618),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_672),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_603),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_666),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_669),
.A2(n_549),
.B1(n_459),
.B2(n_441),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_674),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_620),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_669),
.B(n_525),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_603),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_605),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_674),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_675),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_675),
.B(n_553),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_596),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_675),
.B(n_530),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_668),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_584),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_625),
.A2(n_537),
.B1(n_550),
.B2(n_545),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_595),
.Y(n_765)
);

BUFx6f_ASAP7_75t_SL g766 ( 
.A(n_651),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_668),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_668),
.A2(n_447),
.B1(n_440),
.B2(n_416),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_613),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_668),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_584),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_671),
.B(n_265),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_659),
.B(n_394),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_607),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_607),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_608),
.B(n_537),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_653),
.B(n_545),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_637),
.B(n_485),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_651),
.A2(n_532),
.B1(n_432),
.B2(n_559),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_653),
.B(n_550),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_598),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_655),
.B(n_584),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_652),
.B(n_532),
.Y(n_783)
);

NOR2x1p5_ASAP7_75t_L g784 ( 
.A(n_641),
.B(n_522),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_613),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_666),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_666),
.Y(n_787)
);

BUFx4f_ASAP7_75t_L g788 ( 
.A(n_586),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_615),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_615),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_655),
.B(n_568),
.Y(n_791)
);

OR2x2_ASAP7_75t_SL g792 ( 
.A(n_667),
.B(n_480),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_644),
.B(n_568),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_SL g794 ( 
.A(n_645),
.B(n_369),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_584),
.Y(n_795)
);

AND2x6_ASAP7_75t_L g796 ( 
.A(n_647),
.B(n_237),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_650),
.B(n_575),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_666),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_658),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_660),
.B(n_575),
.C(n_522),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_586),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_608),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_589),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_609),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_589),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_609),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_609),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_582),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_612),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_612),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_661),
.B(n_244),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_663),
.B(n_250),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_609),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_590),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_601),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_590),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_610),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_670),
.B(n_498),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_617),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_610),
.B(n_269),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_610),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_593),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_673),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_627),
.B(n_499),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_628),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_593),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_610),
.B(n_379),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_626),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_628),
.B(n_503),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_690),
.B(n_594),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_691),
.B(n_594),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_702),
.B(n_706),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_597),
.Y(n_834)
);

O2A1O1Ixp5_ASAP7_75t_L g835 ( 
.A1(n_681),
.A2(n_649),
.B(n_647),
.C(n_600),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_702),
.A2(n_509),
.B(n_311),
.C(n_431),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_734),
.B(n_394),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_749),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_734),
.B(n_394),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_700),
.B(n_597),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_725),
.Y(n_841)
);

AND2x4_ASAP7_75t_SL g842 ( 
.A(n_686),
.B(n_664),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_749),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_786),
.Y(n_844)
);

BUFx6f_ASAP7_75t_SL g845 ( 
.A(n_686),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_733),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_694),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_778),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_600),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_768),
.A2(n_270),
.B1(n_397),
.B2(n_376),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_722),
.B(n_602),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_678),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_786),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_683),
.B(n_395),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_776),
.B(n_388),
.C(n_377),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

AND2x6_ASAP7_75t_SL g857 ( 
.A(n_727),
.B(n_561),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_731),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_722),
.B(n_761),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_740),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_768),
.A2(n_443),
.B1(n_261),
.B2(n_271),
.C(n_444),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_742),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_763),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_761),
.B(n_602),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_703),
.B(n_506),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_679),
.B(n_348),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_705),
.B(n_394),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_705),
.B(n_750),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_774),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_726),
.B(n_606),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_704),
.A2(n_514),
.B1(n_517),
.B2(n_512),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_818),
.B(n_563),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_705),
.B(n_394),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_677),
.A2(n_720),
.B(n_698),
.C(n_729),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_798),
.Y(n_877)
);

OAI221xp5_ASAP7_75t_L g878 ( 
.A1(n_750),
.A2(n_567),
.B1(n_564),
.B2(n_565),
.C(n_566),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_717),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_745),
.B(n_570),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_798),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_705),
.B(n_394),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_726),
.B(n_606),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_763),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_710),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_737),
.B(n_759),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_772),
.B(n_394),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_709),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_783),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_771),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_800),
.B(n_824),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_771),
.Y(n_893)
);

AND2x6_ASAP7_75t_SL g894 ( 
.A(n_727),
.B(n_571),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_714),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_682),
.A2(n_338),
.B1(n_328),
.B2(n_325),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_795),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_737),
.B(n_629),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_776),
.B(n_393),
.C(n_389),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_772),
.B(n_262),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_759),
.B(n_629),
.Y(n_901)
);

AO221x1_ASAP7_75t_L g902 ( 
.A1(n_741),
.A2(n_685),
.B1(n_295),
.B2(n_299),
.C(n_277),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_694),
.B(n_649),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_694),
.B(n_293),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_729),
.A2(n_573),
.B(n_574),
.C(n_578),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_694),
.B(n_626),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_801),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_718),
.Y(n_908)
);

BUFx8_ASAP7_75t_L g909 ( 
.A(n_799),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_694),
.B(n_626),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_728),
.A2(n_732),
.B1(n_698),
.B2(n_720),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_762),
.B(n_626),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_783),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_728),
.A2(n_408),
.B1(n_410),
.B2(n_314),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_680),
.B(n_241),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_767),
.B(n_636),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_713),
.B(n_266),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_770),
.B(n_636),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_803),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_636),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_753),
.B(n_355),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_787),
.B(n_636),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_732),
.B(n_360),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_365),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_677),
.A2(n_406),
.B(n_450),
.C(n_449),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_709),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_699),
.B(n_788),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_699),
.B(n_375),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_802),
.B(n_398),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_764),
.B(n_585),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_783),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_693),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_795),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_809),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_695),
.B(n_241),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_810),
.B(n_420),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_823),
.B(n_652),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_788),
.B(n_296),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_697),
.A2(n_353),
.B1(n_301),
.B2(n_303),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_723),
.B(n_304),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_723),
.B(n_676),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_711),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_811),
.B(n_242),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_723),
.B(n_306),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_803),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_738),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_777),
.B(n_309),
.Y(n_947)
);

INVxp33_ASAP7_75t_L g948 ( 
.A(n_701),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_793),
.B(n_580),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_811),
.B(n_242),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_780),
.A2(n_312),
.B1(n_318),
.B2(n_320),
.Y(n_951)
);

AO221x1_ASAP7_75t_L g952 ( 
.A1(n_821),
.A2(n_361),
.B1(n_425),
.B2(n_426),
.C(n_429),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_826),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_820),
.B(n_322),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_791),
.B(n_805),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_684),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_828),
.B(n_323),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_784),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_805),
.B(n_324),
.Y(n_959)
);

AND2x6_ASAP7_75t_SL g960 ( 
.A(n_727),
.B(n_426),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_712),
.B(n_326),
.Y(n_961)
);

BUFx6f_ASAP7_75t_SL g962 ( 
.A(n_686),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_719),
.B(n_330),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_748),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_814),
.B(n_816),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_814),
.B(n_332),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_816),
.B(n_341),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_822),
.B(n_342),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_708),
.B(n_665),
.Y(n_969)
);

OAI22xp33_ASAP7_75t_L g970 ( 
.A1(n_689),
.A2(n_457),
.B1(n_429),
.B2(n_454),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_822),
.B(n_344),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_748),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_812),
.B(n_247),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_825),
.A2(n_457),
.B(n_436),
.C(n_454),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_707),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_782),
.A2(n_396),
.B(n_346),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_779),
.A2(n_444),
.B1(n_437),
.B2(n_438),
.Y(n_977)
);

BUFx5_ASAP7_75t_L g978 ( 
.A(n_738),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_827),
.B(n_806),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_808),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_754),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_769),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_718),
.A2(n_356),
.B1(n_359),
.B2(n_362),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_754),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_808),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_806),
.B(n_366),
.Y(n_986)
);

AO221x1_ASAP7_75t_L g987 ( 
.A1(n_821),
.A2(n_361),
.B1(n_425),
.B2(n_436),
.C(n_437),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_817),
.B(n_368),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_797),
.B(n_401),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_735),
.A2(n_403),
.B(n_371),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_769),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_817),
.B(n_372),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_785),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_751),
.B(n_374),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_757),
.B(n_381),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_794),
.Y(n_996)
);

INVx11_ASAP7_75t_L g997 ( 
.A(n_909),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_859),
.A2(n_792),
.B1(n_689),
.B2(n_812),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_955),
.A2(n_735),
.B(n_773),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_864),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_833),
.B(n_887),
.Y(n_1001)
);

BUFx8_ASAP7_75t_L g1002 ( 
.A(n_845),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_L g1003 ( 
.A1(n_833),
.A2(n_765),
.B1(n_781),
.B2(n_715),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_895),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_981),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_898),
.B(n_744),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_927),
.B(n_708),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_928),
.A2(n_739),
.B(n_736),
.C(n_830),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_907),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_955),
.A2(n_773),
.B(n_716),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_909),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_870),
.A2(n_739),
.B(n_736),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_901),
.B(n_744),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_923),
.A2(n_716),
.B(n_804),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_923),
.A2(n_870),
.B(n_911),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_903),
.A2(n_758),
.B(n_688),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_872),
.B(n_758),
.Y(n_1017)
);

AOI21x1_ASAP7_75t_L g1018 ( 
.A1(n_837),
.A2(n_756),
.B(n_755),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_927),
.B(n_708),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_837),
.A2(n_756),
.B(n_785),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_911),
.A2(n_689),
.B1(n_724),
.B2(n_779),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_841),
.B(n_721),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_883),
.B(n_743),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_868),
.B(n_804),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_980),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_907),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_849),
.A2(n_696),
.B(n_688),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_949),
.Y(n_1028)
);

CKINVDCx10_ASAP7_75t_R g1029 ( 
.A(n_845),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_908),
.B(n_714),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_906),
.A2(n_696),
.B(n_688),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_888),
.A2(n_790),
.B1(n_789),
.B2(n_796),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_886),
.B(n_715),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_865),
.B(n_915),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_910),
.A2(n_696),
.B(n_687),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_917),
.A2(n_804),
.B(n_790),
.C(n_687),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_920),
.A2(n_687),
.B(n_746),
.Y(n_1037)
);

AO32x2_ASAP7_75t_L g1038 ( 
.A1(n_896),
.A2(n_738),
.A3(n_796),
.B1(n_766),
.B2(n_19),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_873),
.A2(n_781),
.B1(n_760),
.B2(n_819),
.Y(n_1039)
);

BUFx4f_ASAP7_75t_L g1040 ( 
.A(n_842),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_956),
.B(n_724),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_922),
.A2(n_746),
.B(n_693),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_915),
.B(n_807),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_943),
.A2(n_433),
.B(n_248),
.C(n_249),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_956),
.B(n_724),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_935),
.A2(n_766),
.B1(n_796),
.B2(n_760),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_835),
.A2(n_813),
.B(n_807),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_935),
.B(n_807),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_979),
.A2(n_693),
.B(n_746),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_839),
.A2(n_813),
.B(n_807),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_852),
.B(n_752),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_962),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_854),
.B(n_813),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_854),
.B(n_813),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_941),
.A2(n_796),
.B1(n_738),
.B2(n_752),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_860),
.B(n_815),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_874),
.B(n_892),
.Y(n_1057)
);

O2A1O1Ixp5_ASAP7_75t_L g1058 ( 
.A1(n_917),
.A2(n_921),
.B(n_839),
.C(n_888),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_965),
.A2(n_746),
.B(n_693),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_948),
.B(n_848),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_941),
.A2(n_421),
.B1(n_248),
.B2(n_249),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_867),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_860),
.B(n_752),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_853),
.A2(n_829),
.B(n_386),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_928),
.A2(n_796),
.B1(n_738),
.B2(n_425),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_996),
.B(n_815),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_879),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_900),
.A2(n_361),
.B(n_16),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_950),
.A2(n_391),
.B1(n_407),
.B2(n_456),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_876),
.A2(n_421),
.B(n_456),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_985),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_989),
.B(n_819),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_950),
.A2(n_973),
.B(n_900),
.C(n_914),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_973),
.B(n_247),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_842),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_846),
.B(n_252),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_914),
.B(n_252),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_880),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_921),
.A2(n_453),
.B(n_452),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_855),
.B(n_253),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_880),
.B(n_438),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_899),
.B(n_253),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_851),
.A2(n_453),
.B1(n_452),
.B2(n_451),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_924),
.A2(n_451),
.B(n_448),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_969),
.B(n_958),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_856),
.B(n_255),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_946),
.B(n_82),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_995),
.A2(n_13),
.B(n_16),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_847),
.A2(n_937),
.B(n_916),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_939),
.B(n_255),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_880),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_919),
.A2(n_448),
.B(n_258),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_946),
.B(n_83),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_970),
.B(n_258),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_836),
.A2(n_259),
.B(n_260),
.C(n_263),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_919),
.A2(n_419),
.B(n_260),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_850),
.B(n_442),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_858),
.B(n_259),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_836),
.A2(n_424),
.B(n_264),
.C(n_268),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_847),
.A2(n_918),
.B(n_912),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_970),
.B(n_890),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_913),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_931),
.A2(n_402),
.B(n_413),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_861),
.B(n_263),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_885),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_847),
.A2(n_904),
.B(n_932),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_995),
.A2(n_430),
.B1(n_268),
.B2(n_272),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_983),
.B(n_264),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_966),
.A2(n_433),
.B(n_419),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_971),
.A2(n_434),
.B(n_424),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_986),
.A2(n_435),
.B(n_430),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_863),
.B(n_272),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_945),
.A2(n_439),
.B(n_435),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_866),
.A2(n_439),
.B(n_434),
.C(n_417),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_951),
.B(n_442),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_864),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_864),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_871),
.B(n_443),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_884),
.B(n_445),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_988),
.A2(n_445),
.B(n_227),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_992),
.A2(n_219),
.B(n_212),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_831),
.A2(n_209),
.B(n_205),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_974),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_1123)
);

INVxp67_ASAP7_75t_SL g1124 ( 
.A(n_885),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_832),
.A2(n_203),
.B(n_199),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_954),
.B(n_194),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_934),
.B(n_29),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_834),
.A2(n_185),
.B(n_180),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_840),
.A2(n_179),
.B(n_175),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_957),
.A2(n_893),
.B(n_933),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_953),
.B(n_30),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_869),
.A2(n_173),
.B(n_169),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_982),
.A2(n_162),
.B(n_160),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_875),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_991),
.A2(n_993),
.B(n_940),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_875),
.A2(n_882),
.B(n_940),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_891),
.A2(n_152),
.B1(n_145),
.B2(n_134),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_891),
.A2(n_893),
.B1(n_897),
.B2(n_933),
.Y(n_1138)
);

AND2x2_ASAP7_75t_SL g1139 ( 
.A(n_850),
.B(n_35),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_947),
.B(n_37),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_944),
.A2(n_133),
.B(n_121),
.Y(n_1141)
);

OAI321xp33_ASAP7_75t_L g1142 ( 
.A1(n_862),
.A2(n_37),
.A3(n_40),
.B1(n_41),
.B2(n_42),
.C(n_47),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_882),
.A2(n_118),
.B(n_116),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_929),
.B(n_41),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_944),
.A2(n_926),
.B(n_889),
.Y(n_1145)
);

OAI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_977),
.A2(n_50),
.B(n_51),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_936),
.B(n_50),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_947),
.B(n_53),
.Y(n_1148)
);

NOR2xp67_ASAP7_75t_L g1149 ( 
.A(n_975),
.B(n_99),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_930),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_838),
.A2(n_96),
.B(n_93),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_994),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_938),
.B(n_959),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_843),
.B(n_61),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_844),
.A2(n_61),
.B(n_62),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_977),
.B(n_62),
.C(n_63),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_942),
.A2(n_66),
.B(n_69),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_974),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_1158)
);

AND3x1_ASAP7_75t_L g1159 ( 
.A(n_905),
.B(n_71),
.C(n_74),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_946),
.B(n_877),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_994),
.A2(n_964),
.B(n_984),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_961),
.B(n_963),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_L g1163 ( 
.A1(n_959),
.A2(n_968),
.B(n_967),
.C(n_938),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_881),
.A2(n_968),
.B1(n_967),
.B2(n_972),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_976),
.A2(n_990),
.B(n_946),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_925),
.A2(n_878),
.B(n_902),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_978),
.B(n_952),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_978),
.B(n_987),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_978),
.B(n_962),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_978),
.A2(n_857),
.B(n_894),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_978),
.B(n_960),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_978),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_833),
.A2(n_868),
.B(n_950),
.C(n_943),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_833),
.B(n_887),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_981),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1173),
.A2(n_1001),
.B1(n_1174),
.B2(n_1153),
.Y(n_1176)
);

AOI221xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1073),
.A2(n_1146),
.B1(n_1021),
.B2(n_1077),
.C(n_1094),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1050),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1034),
.B(n_1023),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1009),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_998),
.A2(n_1108),
.B1(n_1139),
.B2(n_1057),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1015),
.A2(n_1024),
.B(n_999),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1015),
.A2(n_1140),
.B(n_1167),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_999),
.A2(n_1106),
.B(n_1010),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1010),
.A2(n_1017),
.B(n_1013),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1161),
.A2(n_1100),
.B(n_1037),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1004),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1058),
.A2(n_1163),
.B(n_1014),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1067),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1100),
.A2(n_1012),
.B(n_1042),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1165),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1175),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1030),
.B(n_1033),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1053),
.B(n_1054),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1006),
.A2(n_1130),
.B(n_1162),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1071),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1000),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1026),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1165),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1116),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1062),
.B(n_1097),
.Y(n_1202)
);

OAI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1101),
.A2(n_1156),
.B1(n_1078),
.B2(n_1091),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1157),
.A2(n_1088),
.B1(n_1068),
.B2(n_1150),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1089),
.A2(n_1014),
.B(n_1008),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1016),
.A2(n_1136),
.B(n_1035),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1089),
.A2(n_1027),
.B(n_1031),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1041),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1116),
.B(n_1000),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1142),
.A2(n_1123),
.B(n_1158),
.C(n_1152),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1145),
.A2(n_1135),
.B(n_1036),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1168),
.A2(n_1172),
.B(n_1032),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1055),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_SL g1214 ( 
.A1(n_1148),
.A2(n_1147),
.B(n_1144),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1081),
.B(n_1066),
.Y(n_1215)
);

NAND2x1_ASAP7_75t_L g1216 ( 
.A(n_1000),
.B(n_1117),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1138),
.A2(n_1164),
.B(n_1160),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1105),
.A2(n_1124),
.B(n_1126),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1160),
.A2(n_1132),
.B(n_1143),
.Y(n_1219)
);

AOI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1082),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1007),
.A2(n_1019),
.B(n_1064),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1041),
.B(n_1045),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1117),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1166),
.A2(n_1120),
.B(n_1116),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1070),
.A2(n_1166),
.B(n_1044),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1075),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1087),
.A2(n_1093),
.B(n_1154),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_SL g1228 ( 
.A1(n_1121),
.A2(n_1125),
.B(n_1129),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1229)
);

AOI21xp33_ASAP7_75t_L g1230 ( 
.A1(n_1060),
.A2(n_1099),
.B(n_1115),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1045),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1087),
.A2(n_1093),
.B(n_1169),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1056),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1102),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1114),
.A2(n_1083),
.B1(n_1131),
.B2(n_1127),
.C(n_1079),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1092),
.A2(n_1113),
.B(n_1096),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1111),
.A2(n_1084),
.B(n_1109),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1111),
.A2(n_1084),
.B(n_1109),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1086),
.A2(n_1098),
.B(n_1104),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1112),
.B(n_1119),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1118),
.B(n_1076),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1046),
.B(n_1069),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1121),
.A2(n_1151),
.B(n_1122),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1110),
.A2(n_1128),
.B(n_1125),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1072),
.A2(n_1090),
.B1(n_1171),
.B2(n_1003),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1122),
.A2(n_1129),
.B(n_1128),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1137),
.A2(n_1155),
.B(n_1110),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1134),
.Y(n_1248)
);

AOI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1149),
.A2(n_1051),
.B(n_1079),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1063),
.B(n_1170),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1065),
.A2(n_1061),
.B(n_1159),
.Y(n_1252)
);

AOI221x1_ASAP7_75t_L g1253 ( 
.A1(n_1103),
.A2(n_1039),
.B1(n_1038),
.B2(n_1095),
.C(n_1107),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1038),
.A2(n_1085),
.B(n_1040),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1038),
.A2(n_1040),
.A3(n_1002),
.B(n_1029),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1002),
.B(n_1011),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1052),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_997),
.A2(n_1047),
.B(n_1018),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1173),
.B(n_1073),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1005),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1173),
.A2(n_1015),
.B(n_1058),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1173),
.B(n_1001),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1265)
);

NOR2x1_ASAP7_75t_SL g1266 ( 
.A(n_1116),
.B(n_870),
.Y(n_1266)
);

AOI31xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1094),
.A2(n_914),
.A3(n_850),
.B(n_862),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1025),
.B(n_980),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1015),
.A2(n_887),
.B(n_1140),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1005),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1071),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1009),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1173),
.A2(n_1174),
.B(n_1001),
.C(n_1073),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1002),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1173),
.B(n_1073),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1173),
.A2(n_833),
.B1(n_1073),
.B2(n_1174),
.C(n_1001),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1173),
.A2(n_1073),
.B(n_1174),
.C(n_1001),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1028),
.B(n_956),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1173),
.A2(n_833),
.B(n_854),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1028),
.B(n_956),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1002),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1173),
.A2(n_1015),
.B(n_1058),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1297)
);

AOI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1173),
.A2(n_833),
.B(n_854),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_1116),
.B(n_1000),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1173),
.B(n_1073),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1071),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1067),
.Y(n_1304)
);

INVx5_ASAP7_75t_L g1305 ( 
.A(n_1000),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1028),
.B(n_854),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1000),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1173),
.A2(n_1015),
.B(n_1058),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1009),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1173),
.A2(n_1073),
.B(n_833),
.C(n_1001),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1173),
.A2(n_1015),
.B(n_1058),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1116),
.B(n_1000),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1173),
.A2(n_1073),
.B(n_833),
.C(n_1001),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1071),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1001),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1173),
.A2(n_1015),
.B(n_1058),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1047),
.A2(n_1018),
.B(n_1020),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1015),
.A2(n_1048),
.B(n_1043),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1001),
.B(n_1174),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1173),
.A2(n_833),
.B1(n_1174),
.B2(n_1001),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1201),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1199),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1193),
.A2(n_1267),
.B1(n_1263),
.B2(n_1318),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1202),
.B(n_1306),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1250),
.B(n_1222),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1197),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1250),
.B(n_1284),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1264),
.B(n_1265),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1273),
.Y(n_1333)
);

NOR2x1_ASAP7_75t_SL g1334 ( 
.A(n_1201),
.B(n_1305),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1180),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_L g1336 ( 
.A1(n_1286),
.A2(n_1298),
.B(n_1177),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1283),
.B(n_1285),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1193),
.B(n_1241),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1292),
.B(n_1297),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1302),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1305),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1182),
.A2(n_1184),
.B(n_1260),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1312),
.A2(n_1323),
.B1(n_1324),
.B2(n_1318),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1260),
.A2(n_1301),
.B(n_1279),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1226),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1279),
.A2(n_1301),
.B(n_1268),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1220),
.A2(n_1181),
.B1(n_1263),
.B2(n_1242),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1278),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1179),
.B(n_1176),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1250),
.B(n_1189),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1240),
.B(n_1215),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1281),
.B(n_1275),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1208),
.B(n_1231),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1317),
.B(n_1196),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1259),
.A2(n_1322),
.B(n_1270),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1245),
.A2(n_1251),
.B1(n_1233),
.B2(n_1281),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1275),
.B(n_1311),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1316),
.B(n_1282),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1269),
.B(n_1304),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1223),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1204),
.A2(n_1210),
.B1(n_1282),
.B2(n_1236),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1236),
.B(n_1225),
.C(n_1230),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1250),
.B(n_1284),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1274),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1239),
.B(n_1271),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1192),
.Y(n_1367)
);

OR2x6_ASAP7_75t_L g1368 ( 
.A(n_1234),
.B(n_1232),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1187),
.Y(n_1369)
);

INVx3_ASAP7_75t_SL g1370 ( 
.A(n_1257),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1309),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1287),
.B(n_1203),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1305),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1259),
.A2(n_1322),
.B(n_1268),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1287),
.B(n_1251),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1234),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1234),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1204),
.A2(n_1183),
.B1(n_1252),
.B2(n_1237),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1294),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1257),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1235),
.A2(n_1238),
.B1(n_1254),
.B2(n_1194),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1305),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1244),
.A2(n_1314),
.B(n_1295),
.C(n_1308),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1257),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1257),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1223),
.B(n_1198),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1261),
.B(n_1272),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1255),
.B(n_1198),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1209),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1248),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1255),
.B(n_1319),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1307),
.B(n_1216),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1262),
.B(n_1280),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1256),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1307),
.B(n_1258),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1229),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1255),
.B(n_1249),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1307),
.B(n_1266),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1300),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1246),
.A2(n_1224),
.B(n_1247),
.C(n_1195),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1212),
.B(n_1221),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1300),
.Y(n_1403)
);

AOI21xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1227),
.A2(n_1315),
.B(n_1188),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1315),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1280),
.B(n_1296),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1246),
.A2(n_1207),
.B(n_1224),
.C(n_1205),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1288),
.B(n_1296),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1195),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1217),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1219),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1289),
.B(n_1313),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1190),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1243),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1218),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1290),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1211),
.A2(n_1205),
.B(n_1185),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1218),
.B(n_1178),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1228),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1191),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1185),
.B(n_1207),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1200),
.A2(n_1186),
.B(n_1206),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1291),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1214),
.A2(n_1001),
.B1(n_1174),
.B2(n_1173),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1321),
.B(n_1320),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1214),
.B(n_1197),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1278),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1302),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1264),
.A2(n_1001),
.B1(n_1174),
.B2(n_1173),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1199),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1234),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1302),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1250),
.B(n_1222),
.Y(n_1436)
);

BUFx8_ASAP7_75t_SL g1437 ( 
.A(n_1278),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1264),
.B(n_1001),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1213),
.A2(n_1182),
.B(n_1184),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1197),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1199),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1199),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1199),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1264),
.B(n_1001),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1286),
.A2(n_1139),
.B1(n_1298),
.B2(n_1220),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1201),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1264),
.B(n_1001),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1199),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1264),
.A2(n_1001),
.B1(n_1174),
.B2(n_1173),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1234),
.B(n_1004),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1234),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1197),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1264),
.B(n_1001),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1180),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1305),
.B(n_1307),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1180),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1180),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1305),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1199),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1180),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1197),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1305),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1199),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1234),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1202),
.B(n_1306),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1187),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1264),
.B(n_1001),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1180),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1197),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1213),
.A2(n_1182),
.B(n_1184),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_SL g1471 ( 
.A1(n_1286),
.A2(n_1173),
.B(n_1073),
.C(n_1298),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1197),
.Y(n_1472)
);

OR2x6_ASAP7_75t_SL g1473 ( 
.A(n_1256),
.B(n_895),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1250),
.B(n_1222),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1264),
.A2(n_1001),
.B1(n_1174),
.B2(n_1173),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1199),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1187),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1196),
.B(n_980),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1278),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1197),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1193),
.B(n_1030),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1262),
.A2(n_1308),
.B(n_1295),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1339),
.B(n_1332),
.Y(n_1483)
);

INVx11_ASAP7_75t_L g1484 ( 
.A(n_1384),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1327),
.B(n_1348),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1363),
.A2(n_1445),
.B(n_1481),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1437),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1412),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1327),
.A2(n_1352),
.B1(n_1362),
.B2(n_1350),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1335),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1332),
.B(n_1337),
.Y(n_1491)
);

CKINVDCx11_ASAP7_75t_R g1492 ( 
.A(n_1349),
.Y(n_1492)
);

INVx11_ASAP7_75t_L g1493 ( 
.A(n_1430),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1357),
.A2(n_1372),
.B1(n_1328),
.B2(n_1465),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1407),
.A2(n_1374),
.B(n_1356),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1365),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1371),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1454),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1456),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1457),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1460),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1342),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1468),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1330),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1361),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1326),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1338),
.A2(n_1340),
.B1(n_1467),
.B2(n_1447),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1433),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1441),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1442),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1439),
.A2(n_1470),
.B(n_1366),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1340),
.B(n_1350),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1438),
.B(n_1444),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1443),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1448),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1438),
.A2(n_1444),
.B1(n_1467),
.B2(n_1453),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1459),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1342),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1463),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1447),
.B(n_1453),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1476),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_1360),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1361),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1330),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1362),
.A2(n_1353),
.B1(n_1391),
.B2(n_1359),
.Y(n_1527)
);

INVx4_ASAP7_75t_R g1528 ( 
.A(n_1369),
.Y(n_1528)
);

BUFx2_ASAP7_75t_R g1529 ( 
.A(n_1370),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1466),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1387),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1353),
.A2(n_1359),
.B1(n_1336),
.B2(n_1344),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1432),
.B(n_1449),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1342),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1417),
.A2(n_1344),
.B1(n_1383),
.B2(n_1480),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1461),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1469),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1336),
.A2(n_1475),
.B1(n_1358),
.B2(n_1355),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1358),
.A2(n_1378),
.B1(n_1399),
.B2(n_1429),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1399),
.A2(n_1429),
.B1(n_1482),
.B2(n_1375),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1401),
.A2(n_1343),
.B(n_1406),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1347),
.A2(n_1422),
.B(n_1411),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1370),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1429),
.A2(n_1482),
.B1(n_1478),
.B2(n_1397),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1379),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1427),
.A2(n_1385),
.B1(n_1394),
.B2(n_1345),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1341),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1342),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1431),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1477),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1450),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1406),
.A2(n_1408),
.B(n_1414),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_R g1554 ( 
.A(n_1380),
.B(n_1440),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1367),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1386),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1388),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1418),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1386),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1376),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1408),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1373),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1400),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1354),
.B(n_1435),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1333),
.A2(n_1480),
.B1(n_1452),
.B2(n_1472),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1403),
.Y(n_1566)
);

BUFx2_ASAP7_75t_SL g1567 ( 
.A(n_1351),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1405),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1329),
.A2(n_1474),
.B1(n_1436),
.B2(n_1402),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1404),
.A2(n_1366),
.B(n_1381),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1329),
.A2(n_1474),
.B1(n_1436),
.B2(n_1333),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1405),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1368),
.B(n_1423),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1415),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1331),
.A2(n_1364),
.B1(n_1368),
.B2(n_1393),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1473),
.A2(n_1346),
.B1(n_1464),
.B2(n_1451),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1376),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1393),
.B(n_1419),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1455),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1376),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1409),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1409),
.Y(n_1582)
);

AOI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1471),
.A2(n_1464),
.B1(n_1451),
.B2(n_1434),
.C1(n_1377),
.C2(n_1420),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1434),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1434),
.Y(n_1585)
);

INVx11_ASAP7_75t_L g1586 ( 
.A(n_1451),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1464),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1455),
.Y(n_1588)
);

AOI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1416),
.A2(n_1410),
.B(n_1426),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1413),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1428),
.A2(n_1423),
.B(n_1398),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1389),
.Y(n_1592)
);

BUFx8_ASAP7_75t_L g1593 ( 
.A(n_1398),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1428),
.A2(n_1425),
.B(n_1334),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1396),
.A2(n_1325),
.B1(n_1373),
.B2(n_1382),
.Y(n_1595)
);

CKINVDCx11_ASAP7_75t_R g1596 ( 
.A(n_1382),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1446),
.A2(n_1392),
.B1(n_1325),
.B2(n_1458),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1462),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1446),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1446),
.A2(n_1139),
.B1(n_1193),
.B2(n_640),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1458),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1462),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1335),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1335),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1335),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1327),
.B(n_1263),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1335),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1335),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1341),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1335),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1339),
.B(n_1332),
.Y(n_1611)
);

BUFx10_ASAP7_75t_L g1612 ( 
.A(n_1360),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1327),
.B(n_1263),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1327),
.B(n_1263),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1361),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1341),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1335),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1335),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1466),
.B(n_895),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1335),
.Y(n_1620)
);

OR2x6_ASAP7_75t_L g1621 ( 
.A(n_1368),
.B(n_1345),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1335),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1390),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1412),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1421),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1349),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1412),
.Y(n_1628)
);

AO21x1_ASAP7_75t_L g1629 ( 
.A1(n_1362),
.A2(n_1279),
.B(n_1260),
.Y(n_1629)
);

AOI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1424),
.A2(n_1279),
.B(n_1260),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1330),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1339),
.A2(n_1173),
.B1(n_1193),
.B2(n_1332),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1421),
.Y(n_1633)
);

AO21x1_ASAP7_75t_SL g1634 ( 
.A1(n_1336),
.A2(n_1378),
.B(n_1225),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1335),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1348),
.A2(n_1139),
.B1(n_1220),
.B2(n_1286),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1335),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1335),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1335),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1335),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1335),
.Y(n_1641)
);

BUFx2_ASAP7_75t_R g1642 ( 
.A(n_1437),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1412),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1488),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1548),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1600),
.A2(n_1636),
.B1(n_1485),
.B2(n_1613),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1495),
.B(n_1515),
.Y(n_1647)
);

NAND2x1_ASAP7_75t_L g1648 ( 
.A(n_1573),
.B(n_1621),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1520),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1624),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1624),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1591),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1551),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1573),
.B(n_1621),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1520),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1495),
.B(n_1515),
.Y(n_1656)
);

BUFx2_ASAP7_75t_SL g1657 ( 
.A(n_1552),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1623),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1522),
.B(n_1483),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1609),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1553),
.B(n_1591),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1628),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1537),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1606),
.B(n_1613),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1611),
.B(n_1616),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1643),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1606),
.B(n_1614),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1591),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1614),
.B(n_1557),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1558),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

AO21x2_ASAP7_75t_L g1672 ( 
.A1(n_1570),
.A2(n_1513),
.B(n_1589),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1537),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1507),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1507),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1561),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1553),
.A2(n_1542),
.B(n_1632),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1525),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1486),
.A2(n_1489),
.B(n_1536),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1574),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1553),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1520),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1485),
.B(n_1514),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1520),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1582),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1582),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1506),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1526),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1538),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1514),
.B(n_1527),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1525),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1615),
.Y(n_1694)
);

BUFx10_ASAP7_75t_L g1695 ( 
.A(n_1530),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1615),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1590),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1551),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1509),
.A2(n_1518),
.B(n_1547),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1594),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1581),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1625),
.B(n_1633),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1543),
.A2(n_1630),
.B(n_1496),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1531),
.B(n_1539),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1496),
.A2(n_1542),
.B(n_1578),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1581),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1621),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1545),
.B(n_1573),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1621),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1490),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1573),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1629),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1497),
.Y(n_1713)
);

BUFx12f_ASAP7_75t_L g1714 ( 
.A(n_1492),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1498),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1633),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1499),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1496),
.A2(n_1503),
.B(n_1627),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1500),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1550),
.B(n_1564),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1501),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1502),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1505),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1603),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1631),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1604),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_R g1727 ( 
.A(n_1492),
.B(n_1532),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1634),
.B(n_1533),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1605),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1607),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1608),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1610),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1594),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1617),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1618),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1620),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1634),
.B(n_1540),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1622),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1638),
.B(n_1639),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1640),
.B(n_1641),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1619),
.B(n_1530),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1503),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1633),
.B(n_1599),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1593),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1593),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1568),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1627),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1566),
.A2(n_1494),
.B(n_1572),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1627),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1508),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1510),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1556),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1575),
.B(n_1516),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1559),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1511),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1517),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1519),
.B(n_1523),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1555),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1601),
.A2(n_1602),
.B(n_1597),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1521),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1563),
.B(n_1569),
.Y(n_1763)
);

AO21x1_ASAP7_75t_L g1764 ( 
.A1(n_1576),
.A2(n_1562),
.B(n_1565),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1583),
.B(n_1585),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1535),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1535),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1549),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1664),
.B(n_1612),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1711),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1739),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1664),
.B(n_1612),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1660),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1680),
.A2(n_1571),
.B1(n_1592),
.B2(n_1538),
.C(n_1567),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1682),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1690),
.B(n_1612),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1682),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1700),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1701),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1667),
.B(n_1524),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1658),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1669),
.B(n_1524),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1654),
.B(n_1707),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1699),
.A2(n_1728),
.B1(n_1737),
.B2(n_1657),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1648),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1711),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1669),
.B(n_1549),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1684),
.B(n_1549),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1700),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1701),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1707),
.B(n_1580),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1738),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1700),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1665),
.Y(n_1795)
);

INVx5_ASAP7_75t_SL g1796 ( 
.A(n_1654),
.Y(n_1796)
);

OA211x2_ASAP7_75t_L g1797 ( 
.A1(n_1648),
.A2(n_1595),
.B(n_1584),
.C(n_1529),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1678),
.A2(n_1579),
.B(n_1562),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1709),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1761),
.B(n_1552),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1709),
.B(n_1577),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1692),
.B(n_1677),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1677),
.B(n_1579),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1647),
.B(n_1593),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1728),
.A2(n_1554),
.B(n_1598),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1725),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1710),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1710),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1656),
.B(n_1588),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1674),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1674),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1706),
.B(n_1560),
.Y(n_1812)
);

OR2x6_ASAP7_75t_L g1813 ( 
.A(n_1654),
.B(n_1504),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1737),
.B(n_1587),
.Y(n_1814)
);

OR2x2_ASAP7_75t_SL g1815 ( 
.A(n_1708),
.B(n_1504),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1706),
.B(n_1598),
.Y(n_1816)
);

AO31x2_ASAP7_75t_L g1817 ( 
.A1(n_1712),
.A2(n_1733),
.A3(n_1697),
.B(n_1670),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1713),
.B(n_1544),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1713),
.B(n_1717),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1717),
.B(n_1544),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1724),
.B(n_1562),
.Y(n_1821)
);

NAND2xp33_ASAP7_75t_R g1822 ( 
.A(n_1653),
.B(n_1642),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1675),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1653),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1724),
.B(n_1596),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1646),
.A2(n_1532),
.B1(n_1626),
.B2(n_1596),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1729),
.Y(n_1827)
);

NAND2xp33_ASAP7_75t_R g1828 ( 
.A(n_1698),
.B(n_1528),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1729),
.B(n_1626),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1731),
.B(n_1546),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1731),
.B(n_1546),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1734),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1652),
.B(n_1484),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1668),
.B(n_1484),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1739),
.B(n_1487),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1694),
.B(n_1586),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1675),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1740),
.B(n_1487),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1659),
.B(n_1586),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1740),
.B(n_1493),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1741),
.B(n_1644),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1776),
.B(n_1688),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_SL g1844 ( 
.A1(n_1774),
.A2(n_1727),
.B(n_1746),
.Y(n_1844)
);

OAI21xp33_ASAP7_75t_SL g1845 ( 
.A1(n_1800),
.A2(n_1805),
.B(n_1802),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1806),
.B(n_1689),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1826),
.A2(n_1704),
.B1(n_1645),
.B2(n_1755),
.C(n_1720),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1788),
.B(n_1661),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1779),
.B(n_1650),
.Y(n_1849)
);

NAND4xp25_ASAP7_75t_SL g1850 ( 
.A(n_1785),
.B(n_1764),
.C(n_1765),
.D(n_1712),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1791),
.B(n_1650),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_SL g1852 ( 
.A(n_1824),
.B(n_1714),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1782),
.B(n_1651),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1769),
.B(n_1657),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1771),
.B(n_1661),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1769),
.B(n_1662),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1772),
.B(n_1662),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1772),
.B(n_1780),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1803),
.B(n_1661),
.Y(n_1859)
);

NAND4xp25_ASAP7_75t_L g1860 ( 
.A(n_1795),
.B(n_1752),
.C(n_1755),
.D(n_1765),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1815),
.A2(n_1698),
.B1(n_1745),
.B2(n_1746),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1818),
.A2(n_1764),
.B1(n_1763),
.B2(n_1714),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1800),
.A2(n_1752),
.B(n_1742),
.Y(n_1863)
);

OA21x2_ASAP7_75t_L g1864 ( 
.A1(n_1790),
.A2(n_1705),
.B(n_1703),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1810),
.Y(n_1865)
);

OAI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1809),
.A2(n_1763),
.B(n_1671),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1773),
.A2(n_1722),
.B1(n_1723),
.B2(n_1730),
.C(n_1715),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1789),
.B(n_1718),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1833),
.A2(n_1825),
.B(n_1789),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1770),
.B(n_1672),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1770),
.B(n_1672),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1666),
.Y(n_1872)
);

OAI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1804),
.A2(n_1745),
.B1(n_1691),
.B2(n_1673),
.C(n_1663),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1798),
.B(n_1671),
.C(n_1756),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1842),
.B(n_1679),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1818),
.A2(n_1744),
.B(n_1743),
.Y(n_1876)
);

OA21x2_ASAP7_75t_L g1877 ( 
.A1(n_1790),
.A2(n_1705),
.B(n_1703),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1816),
.B(n_1749),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1787),
.B(n_1672),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1819),
.B(n_1679),
.Y(n_1880)
);

NOR3xp33_ASAP7_75t_SL g1881 ( 
.A(n_1822),
.B(n_1768),
.C(n_1767),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1829),
.A2(n_1744),
.B(n_1702),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1819),
.B(n_1696),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1833),
.B(n_1696),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1783),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1787),
.B(n_1799),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1811),
.B(n_1747),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1783),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1823),
.B(n_1749),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1838),
.B(n_1749),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1801),
.B(n_1719),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1801),
.B(n_1721),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1816),
.B(n_1726),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1815),
.A2(n_1673),
.B1(n_1663),
.B2(n_1691),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1825),
.B(n_1732),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1792),
.B(n_1829),
.C(n_1820),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1807),
.B(n_1808),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1820),
.A2(n_1735),
.B1(n_1751),
.B2(n_1753),
.C(n_1757),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_L g1899 ( 
.A(n_1840),
.B(n_1754),
.C(n_1716),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1807),
.B(n_1686),
.Y(n_1900)
);

OAI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1830),
.A2(n_1744),
.B1(n_1743),
.B2(n_1748),
.C(n_1750),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1830),
.B(n_1683),
.C(n_1750),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1808),
.B(n_1686),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1831),
.B(n_1683),
.C(n_1750),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1831),
.B(n_1754),
.C(n_1716),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_L g1906 ( 
.A(n_1786),
.B(n_1821),
.C(n_1812),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1827),
.B(n_1687),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1836),
.A2(n_1758),
.B1(n_1760),
.B2(n_1762),
.C(n_1741),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1827),
.B(n_1687),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1832),
.B(n_1676),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_L g1911 ( 
.A1(n_1814),
.A2(n_1762),
.B(n_1760),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1813),
.A2(n_1702),
.B(n_1761),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1832),
.B(n_1681),
.Y(n_1913)
);

NAND3xp33_ASAP7_75t_L g1914 ( 
.A(n_1786),
.B(n_1748),
.C(n_1766),
.Y(n_1914)
);

INVxp67_ASAP7_75t_SL g1915 ( 
.A(n_1889),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1878),
.B(n_1775),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1850),
.A2(n_1797),
.B1(n_1836),
.B2(n_1839),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1885),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1863),
.A2(n_1839),
.B1(n_1759),
.B2(n_1781),
.C(n_1793),
.Y(n_1919)
);

AND2x2_ASAP7_75t_SL g1920 ( 
.A(n_1862),
.B(n_1786),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1888),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1884),
.B(n_1817),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1897),
.Y(n_1923)
);

NOR2x1_ASAP7_75t_SL g1924 ( 
.A(n_1874),
.B(n_1813),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1868),
.B(n_1778),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1868),
.B(n_1778),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1900),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1878),
.B(n_1775),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1890),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1903),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1864),
.Y(n_1931)
);

INVx4_ASAP7_75t_L g1932 ( 
.A(n_1864),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1886),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1864),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1914),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1859),
.B(n_1784),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1848),
.B(n_1794),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1848),
.B(n_1794),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1855),
.B(n_1859),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1880),
.B(n_1883),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1877),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1907),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1909),
.Y(n_1943)
);

NAND2xp67_ASAP7_75t_L g1944 ( 
.A(n_1846),
.B(n_1841),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1862),
.A2(n_1847),
.B1(n_1844),
.B2(n_1908),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1877),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1910),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1887),
.B(n_1817),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1870),
.B(n_1777),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1875),
.B(n_1817),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1870),
.B(n_1777),
.Y(n_1951)
);

INVxp67_ASAP7_75t_L g1952 ( 
.A(n_1886),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1913),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1865),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1852),
.B(n_1695),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1871),
.B(n_1786),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1871),
.B(n_1786),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1849),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1879),
.B(n_1817),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1851),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1879),
.B(n_1817),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1872),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1931),
.Y(n_1963)
);

INVxp67_ASAP7_75t_L g1964 ( 
.A(n_1954),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1935),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1922),
.B(n_1891),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1956),
.B(n_1882),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1918),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1918),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1958),
.B(n_1895),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1921),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1956),
.B(n_1869),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1935),
.Y(n_1973)
);

OAI32xp33_ASAP7_75t_L g1974 ( 
.A1(n_1945),
.A2(n_1935),
.A3(n_1845),
.B1(n_1860),
.B2(n_1828),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1922),
.B(n_1892),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1921),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1956),
.B(n_1876),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1958),
.B(n_1866),
.Y(n_1978)
);

INVxp33_ASAP7_75t_L g1979 ( 
.A(n_1924),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1923),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1931),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1956),
.B(n_1796),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1931),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1923),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1927),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1956),
.B(n_1796),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1927),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1948),
.B(n_1950),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1930),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1937),
.B(n_1796),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1930),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1942),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1934),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1942),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1924),
.B(n_1902),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1943),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1948),
.B(n_1843),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1943),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1950),
.B(n_1853),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1937),
.B(n_1938),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1947),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1947),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1953),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1937),
.B(n_1796),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1953),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1960),
.B(n_1858),
.Y(n_2006)
);

INVxp33_ASAP7_75t_L g2007 ( 
.A(n_1955),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1938),
.B(n_1796),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1916),
.B(n_1893),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1938),
.B(n_1904),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1960),
.B(n_1911),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1949),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1949),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1949),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1916),
.B(n_1928),
.Y(n_2015)
);

NAND4xp25_ASAP7_75t_L g2016 ( 
.A(n_1945),
.B(n_1898),
.C(n_1867),
.D(n_1899),
.Y(n_2016)
);

INVx1_ASAP7_75t_SL g2017 ( 
.A(n_1940),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1919),
.B(n_1856),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1951),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1919),
.B(n_1857),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1963),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1968),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1965),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_2015),
.B(n_1929),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1964),
.B(n_1973),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1969),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2011),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1963),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_2015),
.B(n_1929),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1978),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_2017),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1977),
.B(n_1936),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1977),
.B(n_1939),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_2016),
.B(n_1896),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2018),
.B(n_2020),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1970),
.B(n_1944),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1967),
.B(n_1939),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1995),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_SL g2039 ( 
.A(n_1979),
.B(n_1917),
.C(n_1881),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1971),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1976),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1966),
.B(n_1928),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1980),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1985),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1981),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2007),
.A2(n_1920),
.B1(n_1917),
.B2(n_1861),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1995),
.A2(n_1920),
.B1(n_1797),
.B2(n_1894),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1995),
.B(n_1936),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1984),
.Y(n_2049)
);

OAI221xp5_ASAP7_75t_SL g2050 ( 
.A1(n_1974),
.A2(n_1873),
.B1(n_1901),
.B2(n_1912),
.C(n_1952),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1987),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1967),
.B(n_1939),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2009),
.B(n_1944),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2009),
.B(n_2006),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1981),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_2007),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1983),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1983),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1989),
.B(n_1991),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1992),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1994),
.B(n_1962),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2010),
.B(n_1925),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1996),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1998),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2001),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_2002),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2010),
.B(n_1925),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2003),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1974),
.B(n_1695),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2005),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1982),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1972),
.B(n_1925),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1972),
.B(n_1926),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1993),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2000),
.B(n_1926),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2026),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_2056),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2066),
.Y(n_2078)
);

OA21x2_ASAP7_75t_L g2079 ( 
.A1(n_2038),
.A2(n_1941),
.B(n_1934),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2055),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2034),
.A2(n_1920),
.B1(n_1979),
.B2(n_1982),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2035),
.B(n_1915),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2033),
.B(n_2000),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2055),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2055),
.Y(n_2085)
);

AND3x1_ASAP7_75t_L g2086 ( 
.A(n_2069),
.B(n_1841),
.C(n_1986),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2054),
.B(n_1997),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2026),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_2023),
.B(n_2025),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_2031),
.B(n_1695),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2033),
.B(n_1986),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2040),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_2048),
.B(n_1993),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2021),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2040),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2021),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2027),
.B(n_1915),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2038),
.B(n_1990),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2024),
.B(n_1997),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2028),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2030),
.B(n_1966),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2041),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2024),
.B(n_1975),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2062),
.B(n_1990),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2071),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2070),
.B(n_2044),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2041),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_2048),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_2036),
.B(n_2004),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2043),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2043),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2028),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2045),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2049),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2045),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_2071),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2049),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2078),
.Y(n_2118)
);

NAND3x1_ASAP7_75t_L g2119 ( 
.A(n_2089),
.B(n_2047),
.C(n_2053),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2108),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2077),
.Y(n_2121)
);

NOR2x1_ASAP7_75t_L g2122 ( 
.A(n_2077),
.B(n_2039),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_2108),
.Y(n_2123)
);

OAI21xp33_ASAP7_75t_L g2124 ( 
.A1(n_2081),
.A2(n_2050),
.B(n_2046),
.Y(n_2124)
);

OAI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_2105),
.A2(n_2029),
.B1(n_2042),
.B2(n_2048),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2082),
.A2(n_2059),
.B(n_2060),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_2078),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2083),
.Y(n_2128)
);

NAND3xp33_ASAP7_75t_SL g2129 ( 
.A(n_2105),
.B(n_2116),
.C(n_2097),
.Y(n_2129)
);

CKINVDCx16_ASAP7_75t_R g2130 ( 
.A(n_2090),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2086),
.A2(n_2032),
.B1(n_2022),
.B2(n_2051),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_2098),
.B(n_2032),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2076),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2086),
.A2(n_2032),
.B1(n_2051),
.B2(n_2063),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2076),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2136)
);

NAND4xp25_ASAP7_75t_L g2137 ( 
.A(n_2109),
.B(n_2106),
.C(n_2116),
.D(n_2101),
.Y(n_2137)
);

AO32x1_ASAP7_75t_L g2138 ( 
.A1(n_2080),
.A2(n_2064),
.A3(n_2063),
.B1(n_2065),
.B2(n_2068),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2097),
.B(n_2065),
.C(n_2064),
.Y(n_2139)
);

O2A1O1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_2106),
.A2(n_2029),
.B(n_2068),
.C(n_2057),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2101),
.B(n_2042),
.Y(n_2141)
);

OAI21xp33_ASAP7_75t_L g2142 ( 
.A1(n_2082),
.A2(n_2067),
.B(n_2061),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2091),
.B(n_2067),
.Y(n_2143)
);

OAI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2087),
.A2(n_2099),
.B1(n_2103),
.B2(n_2091),
.C(n_2104),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2083),
.B(n_2037),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2099),
.A2(n_2052),
.B1(n_2037),
.B2(n_1952),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2104),
.A2(n_2052),
.B(n_2072),
.Y(n_2147)
);

OAI21xp33_ASAP7_75t_L g2148 ( 
.A1(n_2087),
.A2(n_2103),
.B(n_2092),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2121),
.B(n_2088),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2118),
.Y(n_2150)
);

AND4x1_ASAP7_75t_L g2151 ( 
.A(n_2122),
.B(n_2092),
.C(n_2095),
.D(n_2088),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2123),
.B(n_2095),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2130),
.B(n_2137),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2136),
.B(n_2093),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2133),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_2132),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2132),
.B(n_2093),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2143),
.B(n_2128),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2122),
.B(n_2102),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2120),
.B(n_2102),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2148),
.B(n_2107),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2147),
.B(n_2093),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2135),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2127),
.B(n_2107),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2144),
.B(n_2110),
.Y(n_2165)
);

NOR3xp33_ASAP7_75t_SL g2166 ( 
.A(n_2129),
.B(n_2124),
.C(n_2125),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2119),
.A2(n_2093),
.B1(n_2117),
.B2(n_2114),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2138),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2138),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2126),
.B(n_2134),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2138),
.Y(n_2171)
);

AOI211xp5_ASAP7_75t_L g2172 ( 
.A1(n_2153),
.A2(n_2140),
.B(n_2139),
.C(n_2131),
.Y(n_2172)
);

OAI211xp5_ASAP7_75t_L g2173 ( 
.A1(n_2167),
.A2(n_2142),
.B(n_2141),
.C(n_2145),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_SL g2174 ( 
.A1(n_2153),
.A2(n_2146),
.B1(n_2079),
.B2(n_2114),
.Y(n_2174)
);

AOI221x1_ASAP7_75t_L g2175 ( 
.A1(n_2171),
.A2(n_2117),
.B1(n_2110),
.B2(n_2111),
.C(n_2084),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2166),
.A2(n_2111),
.B1(n_2115),
.B2(n_2112),
.Y(n_2176)
);

AOI221xp5_ASAP7_75t_L g2177 ( 
.A1(n_2170),
.A2(n_2115),
.B1(n_2113),
.B2(n_2112),
.C(n_2094),
.Y(n_2177)
);

OAI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2151),
.A2(n_2159),
.B(n_2165),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2159),
.A2(n_2079),
.B(n_2080),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2156),
.Y(n_2180)
);

O2A1O1Ixp33_ASAP7_75t_L g2181 ( 
.A1(n_2168),
.A2(n_2115),
.B(n_2113),
.C(n_2112),
.Y(n_2181)
);

OAI211xp5_ASAP7_75t_L g2182 ( 
.A1(n_2165),
.A2(n_2113),
.B(n_2100),
.C(n_2096),
.Y(n_2182)
);

O2A1O1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_2161),
.A2(n_2100),
.B(n_2096),
.C(n_2094),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2149),
.B(n_2094),
.Y(n_2184)
);

OAI21xp33_ASAP7_75t_SL g2185 ( 
.A1(n_2169),
.A2(n_2084),
.B(n_2080),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_2150),
.B(n_2072),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2152),
.Y(n_2187)
);

NOR3xp33_ASAP7_75t_L g2188 ( 
.A(n_2178),
.B(n_2164),
.C(n_2160),
.Y(n_2188)
);

NOR3x1_ASAP7_75t_L g2189 ( 
.A(n_2173),
.B(n_2163),
.C(n_2155),
.Y(n_2189)
);

OA22x2_ASAP7_75t_L g2190 ( 
.A1(n_2176),
.A2(n_2169),
.B1(n_2157),
.B2(n_2162),
.Y(n_2190)
);

NOR3xp33_ASAP7_75t_L g2191 ( 
.A(n_2172),
.B(n_2158),
.C(n_2162),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2180),
.B(n_2154),
.Y(n_2192)
);

NAND2x1p5_ASAP7_75t_L g2193 ( 
.A(n_2184),
.B(n_2157),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_2187),
.B(n_2154),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_2174),
.B(n_2084),
.Y(n_2195)
);

NOR3x1_ASAP7_75t_L g2196 ( 
.A(n_2182),
.B(n_1988),
.C(n_1905),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2186),
.B(n_2096),
.Y(n_2197)
);

OAI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2179),
.A2(n_1988),
.B1(n_1957),
.B2(n_2085),
.Y(n_2198)
);

NOR3x1_ASAP7_75t_L g2199 ( 
.A(n_2185),
.B(n_1906),
.C(n_1975),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_L g2200 ( 
.A(n_2181),
.B(n_2100),
.C(n_2085),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2177),
.B(n_2073),
.Y(n_2201)
);

NAND4xp25_ASAP7_75t_L g2202 ( 
.A(n_2175),
.B(n_2085),
.C(n_2073),
.D(n_2074),
.Y(n_2202)
);

NAND4xp75_ASAP7_75t_L g2203 ( 
.A(n_2189),
.B(n_2079),
.C(n_2183),
.D(n_2074),
.Y(n_2203)
);

AOI211xp5_ASAP7_75t_L g2204 ( 
.A1(n_2188),
.A2(n_2057),
.B(n_2058),
.C(n_2008),
.Y(n_2204)
);

NOR3xp33_ASAP7_75t_L g2205 ( 
.A(n_2192),
.B(n_2058),
.C(n_1837),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2191),
.A2(n_1932),
.B1(n_2075),
.B2(n_1961),
.C(n_1959),
.Y(n_2206)
);

NOR3xp33_ASAP7_75t_L g2207 ( 
.A(n_2194),
.B(n_1837),
.C(n_1835),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2195),
.A2(n_2079),
.B(n_2075),
.Y(n_2208)
);

NAND4xp25_ASAP7_75t_SL g2209 ( 
.A(n_2201),
.B(n_2008),
.C(n_2004),
.D(n_2013),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2197),
.A2(n_1932),
.B1(n_1959),
.B2(n_1961),
.C(n_2013),
.Y(n_2210)
);

AOI211xp5_ASAP7_75t_L g2211 ( 
.A1(n_2200),
.A2(n_1834),
.B(n_1835),
.C(n_1854),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2203),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2205),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2204),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2209),
.A2(n_2190),
.B1(n_2193),
.B2(n_2202),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2207),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2208),
.B(n_2196),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2211),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2206),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_2216),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2218),
.B(n_2199),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2212),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2215),
.B(n_2198),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_2214),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2213),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2217),
.B(n_2079),
.Y(n_2226)
);

OAI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_2223),
.A2(n_2219),
.B(n_2210),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2220),
.B(n_2012),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2221),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2225),
.B(n_2014),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2221),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_2229),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2231),
.Y(n_2233)
);

NAND5xp2_ASAP7_75t_L g2234 ( 
.A(n_2233),
.B(n_2227),
.C(n_2224),
.D(n_2222),
.E(n_2226),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2234),
.A2(n_2233),
.B1(n_2222),
.B2(n_2232),
.Y(n_2235)
);

AOI21xp33_ASAP7_75t_SL g2236 ( 
.A1(n_2234),
.A2(n_2232),
.B(n_2228),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2235),
.A2(n_2224),
.B1(n_2232),
.B2(n_2228),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2236),
.A2(n_2224),
.B1(n_2230),
.B2(n_1999),
.Y(n_2238)
);

CKINVDCx20_ASAP7_75t_R g2239 ( 
.A(n_2237),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2238),
.A2(n_1999),
.B(n_1835),
.Y(n_2240)
);

OAI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2239),
.A2(n_1835),
.B(n_1834),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2241),
.A2(n_2240),
.B1(n_2019),
.B2(n_1933),
.Y(n_2242)
);

AOI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2242),
.A2(n_1932),
.B1(n_1834),
.B2(n_1946),
.C(n_1934),
.Y(n_2243)
);

AOI211xp5_ASAP7_75t_L g2244 ( 
.A1(n_2243),
.A2(n_1655),
.B(n_1685),
.C(n_1649),
.Y(n_2244)
);


endmodule