module real_jpeg_26109_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_64),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_3),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_83),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_83),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_7),
.A2(n_71),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_132),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_132),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_11),
.B(n_107),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_11),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_78),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_11),
.B(n_42),
.C(n_56),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_11),
.B(n_152),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_181),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_11),
.B(n_28),
.C(n_47),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_11),
.A2(n_30),
.B(n_242),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_69),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_69),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_14),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_94)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_16),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_16),
.A2(n_155),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_113),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_112),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_66),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_23),
.A2(n_24),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_25),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_121),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_27),
.B(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_30),
.A2(n_32),
.B(n_34),
.Y(n_99)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_30),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_30),
.A2(n_157),
.B1(n_159),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_30),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_30),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_36),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_36),
.B(n_181),
.Y(n_266)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_40),
.A2(n_49),
.B1(n_91),
.B2(n_124),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_42),
.B(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_50),
.B1(n_52),
.B2(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_45),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_45),
.A2(n_52),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_49),
.A2(n_124),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_49),
.A2(n_177),
.B(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_49),
.B(n_181),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_52),
.B(n_178),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_53),
.B(n_66),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_54),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_54),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_54),
.A2(n_151),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_63),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_55),
.A2(n_127),
.B(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_60),
.B1(n_75),
.B2(n_76),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_59),
.A2(n_70),
.A3(n_76),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_60),
.B(n_75),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_60),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B(n_79),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_73),
.B1(n_78),
.B2(n_131),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_73),
.A2(n_80),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_106),
.B(n_110),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_77),
.A2(n_110),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_84),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B(n_95),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_91),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_91),
.A2(n_230),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_130),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_123),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_150),
.B1(n_152),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_166),
.B(n_290),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_164),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_138),
.B(n_164),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_143),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_145),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_161),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_161),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_159),
.A2(n_255),
.B(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_197),
.B(n_284),
.C(n_289),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_191),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_183),
.C(n_184),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_169),
.A2(n_170),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_183),
.B(n_184),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_278),
.B(n_283),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_231),
.B(n_277),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_220),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_220),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_217),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_203),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B(n_211),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_271),
.B(n_276),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_251),
.B(n_270),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_245),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_245),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_249),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_259),
.B(n_269),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_257),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_264),
.B(n_268),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);


endmodule