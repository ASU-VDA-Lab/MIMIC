module fake_jpeg_31195_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_21),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_46),
.A2(n_41),
.B1(n_30),
.B2(n_35),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_51),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_54),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_62),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_21),
.B(n_4),
.CON(n_68),
.SN(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_73),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_4),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_83),
.Y(n_133)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_89),
.B(n_111),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_91),
.A2(n_103),
.B1(n_109),
.B2(n_129),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_113),
.Y(n_140)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_102),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_50),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_30),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_116),
.B(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_83),
.B1(n_43),
.B2(n_42),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_67),
.B(n_39),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_39),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_35),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_61),
.B1(n_46),
.B2(n_53),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_144),
.Y(n_221)
);

AO22x2_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_79),
.B1(n_71),
.B2(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_138),
.B(n_151),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_81),
.B1(n_59),
.B2(n_84),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_139),
.A2(n_154),
.B1(n_100),
.B2(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_143),
.Y(n_208)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_88),
.B1(n_109),
.B2(n_91),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_145),
.B(n_181),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_61),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_148),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_149),
.B(n_152),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_70),
.B1(n_82),
.B2(n_74),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_175),
.B1(n_123),
.B2(n_93),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_34),
.B(n_33),
.C(n_23),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_20),
.B1(n_23),
.B2(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_159),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_82),
.B1(n_74),
.B2(n_72),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_99),
.B1(n_97),
.B2(n_106),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_87),
.B(n_86),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_166),
.Y(n_190)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_83),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_72),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_183),
.B1(n_7),
.B2(n_8),
.Y(n_216)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_101),
.A2(n_32),
.B1(n_42),
.B2(n_8),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_105),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.Y(n_191)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_124),
.B(n_5),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_5),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_7),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_5),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_112),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_12),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_94),
.C(n_134),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_138),
.C(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_128),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_128),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_209),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_99),
.B1(n_97),
.B2(n_104),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_197),
.A2(n_147),
.B1(n_173),
.B2(n_160),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_218),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_202),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_145),
.B(n_7),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_219),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_104),
.B(n_117),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_151),
.B(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_216),
.B1(n_226),
.B2(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_153),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_161),
.B(n_9),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_168),
.A2(n_144),
.B1(n_137),
.B2(n_138),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_137),
.B1(n_181),
.B2(n_144),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_189),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_206),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_137),
.B1(n_154),
.B2(n_138),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_243),
.B1(n_250),
.B2(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_251),
.C(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_169),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_239),
.A2(n_247),
.B1(n_257),
.B2(n_202),
.Y(n_270)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_139),
.B1(n_180),
.B2(n_162),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_147),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_210),
.B1(n_196),
.B2(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_192),
.C(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_221),
.A2(n_148),
.B1(n_165),
.B2(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_258),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_214),
.A2(n_216),
.B1(n_209),
.B2(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_174),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_261),
.Y(n_281)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_191),
.A2(n_12),
.A3(n_179),
.B1(n_203),
.B2(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_211),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_264),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_285),
.C(n_294),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_217),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_268),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_274),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_270),
.A2(n_237),
.B1(n_253),
.B2(n_242),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_211),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_218),
.C(n_224),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_276),
.B(n_284),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_229),
.A2(n_205),
.B1(n_185),
.B2(n_189),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_199),
.Y(n_278)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_245),
.B(n_213),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_212),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_249),
.A2(n_205),
.B1(n_204),
.B2(n_179),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_207),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_207),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_286),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_227),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_261),
.B(n_204),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_227),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_267),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_212),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_296),
.B(n_271),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_228),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_310),
.C(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_239),
.B1(n_231),
.B2(n_249),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_270),
.B1(n_281),
.B2(n_279),
.Y(n_325)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_231),
.A3(n_232),
.B1(n_243),
.B2(n_237),
.C(n_254),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_266),
.B1(n_286),
.B2(n_290),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_311),
.Y(n_329)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_255),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_237),
.B(n_238),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_238),
.C(n_258),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_256),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_280),
.C(n_275),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_303),
.C(n_297),
.Y(n_328)
);

AOI221xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_273),
.B1(n_292),
.B2(n_264),
.C(n_268),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_319),
.A2(n_276),
.B1(n_283),
.B2(n_266),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_330),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_326),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_334),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_300),
.B(n_263),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_332),
.B1(n_306),
.B2(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_309),
.B(n_248),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_336),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_293),
.Y(n_335)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_272),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_272),
.C(n_287),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_340),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_277),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_305),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_342),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_277),
.B1(n_287),
.B2(n_288),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_345),
.B(n_349),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_351),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_323),
.B(n_307),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_316),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_310),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_355),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_312),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_296),
.C(n_311),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_357),
.C(n_358),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_319),
.C(n_320),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_304),
.C(n_298),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_331),
.A2(n_298),
.B1(n_304),
.B2(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

OA21x2_ASAP7_75t_SL g363 ( 
.A1(n_360),
.A2(n_326),
.B(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_327),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_365),
.Y(n_382)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

OAI22x1_ASAP7_75t_L g366 ( 
.A1(n_359),
.A2(n_329),
.B1(n_325),
.B2(n_327),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_366),
.A2(n_342),
.B1(n_337),
.B2(n_308),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_346),
.B(n_321),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_371),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_321),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_322),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_352),
.A2(n_340),
.B(n_336),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_357),
.C(n_358),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_356),
.B(n_252),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_374),
.A2(n_344),
.B(n_347),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_385),
.C(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_355),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_380),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_377),
.A2(n_378),
.B(n_366),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_351),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_344),
.B1(n_235),
.B2(n_353),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_362),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_235),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_389),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_383),
.A2(n_364),
.B(n_361),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_378),
.B(n_220),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_381),
.A2(n_368),
.B(n_361),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_390),
.B(n_391),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_372),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_385),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_379),
.A2(n_370),
.B(n_215),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_393),
.B(n_381),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_397),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_375),
.C(n_391),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_220),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_394),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_401),
.B(n_402),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_398),
.B(n_220),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_403),
.A2(n_396),
.B(n_400),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_403),
.Y(n_406)
);

XNOR2x2_ASAP7_75t_SL g407 ( 
.A(n_406),
.B(n_405),
.Y(n_407)
);


endmodule