module real_jpeg_30079_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_0),
.A2(n_61),
.B1(n_62),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_0),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_138),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_138),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_138),
.Y(n_259)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_54),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_5),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_186),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_186),
.Y(n_272)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_57),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_9),
.B(n_44),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_44),
.B(n_224),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_184),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_9),
.A2(n_30),
.B(n_33),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_9),
.B(n_134),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_9),
.A2(n_84),
.B1(n_87),
.B2(n_272),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_63),
.Y(n_199)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_165),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_165),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_165),
.Y(n_264)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_48)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_98),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_81),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_21),
.A2(n_22),
.B1(n_71),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_22)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_24),
.A2(n_25),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_40),
.C(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_26),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_26),
.A2(n_32),
.B1(n_93),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_26),
.A2(n_36),
.B(n_94),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_26),
.A2(n_32),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_26),
.A2(n_76),
.B(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_26),
.A2(n_32),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_26),
.A2(n_32),
.B1(n_231),
.B2(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g220 ( 
.A1(n_28),
.A2(n_45),
.A3(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_29),
.B(n_222),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_29),
.A2(n_31),
.B(n_184),
.C(n_251),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_78),
.B(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_32),
.B(n_184),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_35),
.B(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B(n_52),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_41),
.A2(n_52),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_41),
.A2(n_108),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_53),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_42),
.A2(n_48),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_42),
.A2(n_48),
.B1(n_180),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_42),
.A2(n_48),
.B1(n_208),
.B2(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_44),
.B(n_58),
.Y(n_197)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_45),
.A2(n_66),
.B1(n_183),
.B2(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_70),
.B1(n_100),
.B2(n_112),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_64),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_60),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_56),
.A2(n_102),
.B1(n_137),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_56),
.A2(n_102),
.B1(n_164),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B(n_62),
.C(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_57),
.B(n_96),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_57),
.A2(n_65),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g183 ( 
.A(n_62),
.B(n_184),
.CON(n_183),
.SN(n_183)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_74),
.A2(n_110),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_82),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_91),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_95),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_83),
.A2(n_92),
.B1(n_121),
.B2(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B(n_89),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_84),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_84),
.A2(n_87),
.B1(n_156),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_84),
.A2(n_130),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_84),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_85),
.A2(n_90),
.B(n_158),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_85),
.A2(n_86),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_90),
.Y(n_130)
);

INVx11_ASAP7_75t_L g273 ( 
.A(n_86),
.Y(n_273)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_129),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_88),
.A2(n_127),
.B(n_199),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_111),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_144),
.B(n_319),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_140),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_117),
.B(n_140),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_123),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_122),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_123),
.A2(n_124),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_135),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_126),
.B(n_131),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_169),
.B(n_318),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_166),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_146),
.B(n_166),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_153),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_151),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_153),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.C(n_162),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_154),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_159),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_160),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_312),
.B(n_317),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_212),
.B(n_298),
.C(n_311),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_200),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_172),
.B(n_200),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_187),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_174),
.B(n_175),
.C(n_187),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_184),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_189),
.B(n_193),
.C(n_195),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_201),
.A2(n_202),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_297),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_290),
.B(n_296),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_242),
.B(n_289),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_233),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_216),
.B(n_233),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.C(n_229),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_218),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_240),
.C(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_283),
.B(n_288),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_260),
.B(n_282),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_268),
.B(n_281),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_266),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_280),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_309),
.B2(n_310),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_306),
.C(n_310),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule