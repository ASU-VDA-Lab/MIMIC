module fake_netlist_1_3697_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_2), .B(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NOR2x1_ASAP7_75t_L g13 ( .A(n_5), .B(n_4), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_0), .B(n_2), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_15), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_15), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_11), .B(n_14), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_11), .B(n_13), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
NOR2x1p5_ASAP7_75t_L g22 ( .A(n_20), .B(n_1), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_19), .B1(n_21), .B2(n_17), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_17), .B1(n_24), .B2(n_19), .C(n_6), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_29) );
AND3x4_ASAP7_75t_L g30 ( .A(n_29), .B(n_3), .C(n_7), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
BUFx6f_ASAP7_75t_L g32 ( .A(n_28), .Y(n_32) );
OAI221xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_27), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_32), .B1(n_30), .B2(n_33), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
endmodule