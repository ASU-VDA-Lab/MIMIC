module fake_jpeg_2236_n_478 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_478);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_478;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_49),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_39),
.B1(n_42),
.B2(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_20),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_66),
.Y(n_95)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_0),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_71),
.B(n_38),
.C(n_37),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_2),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_3),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_40),
.Y(n_137)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_30),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_17),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_92),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_96),
.B(n_128),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_107),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_39),
.B1(n_20),
.B2(n_22),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_114),
.B1(n_133),
.B2(n_135),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_145),
.C(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_18),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_108),
.B(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_52),
.A2(n_35),
.B1(n_44),
.B2(n_17),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_117),
.B1(n_142),
.B2(n_28),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_130),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_39),
.B1(n_26),
.B2(n_19),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_44),
.B1(n_35),
.B2(n_42),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_124),
.B(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_49),
.B(n_19),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_46),
.Y(n_130)
);

OR2x4_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_31),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_63),
.A2(n_26),
.B1(n_42),
.B2(n_46),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_47),
.A2(n_46),
.B1(n_45),
.B2(n_28),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_4),
.B(n_8),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_37),
.B1(n_45),
.B2(n_40),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_139),
.B(n_141),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_50),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_149),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_89),
.A2(n_45),
.B1(n_38),
.B2(n_37),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_15),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_33),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_154),
.Y(n_213)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_155),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_172),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_58),
.B1(n_68),
.B2(n_64),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_159),
.A2(n_202),
.B1(n_112),
.B2(n_119),
.Y(n_227)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_98),
.A2(n_53),
.B1(n_61),
.B2(n_60),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_163),
.A2(n_167),
.B1(n_186),
.B2(n_192),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_70),
.B1(n_56),
.B2(n_28),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_31),
.B1(n_43),
.B2(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_31),
.B1(n_43),
.B2(n_6),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_108),
.A2(n_43),
.B1(n_4),
.B2(n_6),
.Y(n_167)
);

OA22x2_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_43),
.B1(n_4),
.B2(n_7),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_168),
.A2(n_169),
.B(n_178),
.C(n_166),
.Y(n_251)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_169)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_194),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_189),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_95),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_119),
.B1(n_112),
.B2(n_116),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_9),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_104),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_180),
.A2(n_144),
.B1(n_143),
.B2(n_116),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_10),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_188),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_104),
.A2(n_139),
.B1(n_105),
.B2(n_138),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_11),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_194),
.Y(n_230)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_120),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_12),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_195),
.B(n_204),
.C(n_190),
.Y(n_255)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_12),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_199),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_93),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_127),
.A2(n_14),
.B1(n_15),
.B2(n_121),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_97),
.B(n_15),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_144),
.Y(n_235)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_113),
.A2(n_127),
.B1(n_102),
.B2(n_115),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_126),
.B1(n_132),
.B2(n_143),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_121),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_209),
.B(n_235),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_94),
.B(n_120),
.C(n_110),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_210),
.A2(n_228),
.B(n_191),
.C(n_193),
.D(n_176),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_94),
.B(n_110),
.Y(n_212)
);

OR2x2_ASAP7_75t_SL g279 ( 
.A(n_212),
.B(n_210),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_160),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_187),
.C(n_200),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_94),
.A3(n_147),
.B1(n_102),
.B2(n_115),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_201),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_162),
.A2(n_94),
.B(n_147),
.C(n_126),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_229),
.A2(n_214),
.B1(n_250),
.B2(n_253),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_175),
.A2(n_116),
.B(n_147),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_231),
.A2(n_217),
.B(n_209),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_233),
.A2(n_229),
.B1(n_213),
.B2(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_203),
.B(n_156),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_243),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_177),
.A2(n_156),
.B1(n_163),
.B2(n_192),
.Y(n_239)
);

AO21x2_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_246),
.B(n_253),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_164),
.B(n_177),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_215),
.B(n_225),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_184),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_183),
.B1(n_188),
.B2(n_186),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_170),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_195),
.B(n_168),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_195),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_169),
.B(n_196),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_280),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_262),
.A2(n_269),
.B(n_279),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_263),
.B(n_272),
.Y(n_316)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_265),
.Y(n_315)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_267),
.B(n_288),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_153),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_284),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_152),
.B(n_181),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_298),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_247),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_273),
.B(n_274),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_241),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_252),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_277),
.A2(n_286),
.B(n_207),
.Y(n_321)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_238),
.B(n_219),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_282),
.B(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_283),
.A2(n_292),
.B1(n_232),
.B2(n_250),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_208),
.B(n_220),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_217),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_254),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_240),
.A2(n_236),
.B1(n_223),
.B2(n_218),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_289),
.A2(n_294),
.B1(n_256),
.B2(n_281),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_220),
.B(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_240),
.A2(n_236),
.B1(n_218),
.B2(n_223),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_239),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_214),
.Y(n_298)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_207),
.Y(n_299)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

BUFx4f_ASAP7_75t_SL g300 ( 
.A(n_211),
.Y(n_300)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_259),
.A2(n_221),
.B1(n_232),
.B2(n_228),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_216),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_307),
.C(n_336),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_216),
.C(n_231),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_248),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_221),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_276),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_211),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_330),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_317),
.A2(n_322),
.B(n_333),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_207),
.B1(n_298),
.B2(n_280),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_318),
.A2(n_300),
.B1(n_278),
.B2(n_299),
.Y(n_370)
);

AOI221xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_339),
.B1(n_335),
.B2(n_316),
.C(n_314),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_257),
.A2(n_297),
.B(n_286),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_261),
.B(n_207),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_276),
.A2(n_257),
.B1(n_290),
.B2(n_283),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_269),
.B1(n_295),
.B2(n_300),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_259),
.A2(n_270),
.B1(n_264),
.B2(n_275),
.Y(n_333)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_282),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_261),
.B(n_289),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_294),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_325),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_359),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_353),
.B1(n_367),
.B2(n_369),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_268),
.Y(n_351)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_288),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_354),
.B(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_331),
.Y(n_355)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_356),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_322),
.A2(n_276),
.B1(n_285),
.B2(n_260),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_363),
.B1(n_370),
.B2(n_318),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_277),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_368),
.C(n_307),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_339),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_338),
.A2(n_267),
.B(n_277),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_338),
.B(n_339),
.Y(n_383)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_364),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_320),
.A2(n_276),
.B1(n_260),
.B2(n_270),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_371),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_301),
.B(n_271),
.C(n_279),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_314),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_306),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_363),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_384),
.B1(n_388),
.B2(n_394),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_301),
.C(n_324),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_385),
.C(n_390),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_328),
.B1(n_308),
.B2(n_311),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_324),
.C(n_321),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_325),
.Y(n_387)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_320),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_392),
.B1(n_391),
.B2(n_382),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_320),
.C(n_315),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_351),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_323),
.B1(n_312),
.B2(n_329),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_323),
.C(n_312),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_396),
.C(n_366),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_359),
.C(n_357),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_329),
.Y(n_398)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_385),
.B(n_354),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_383),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_404),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_382),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_403),
.B(n_417),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_344),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_408),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_374),
.B(n_345),
.C(n_344),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_411),
.C(n_414),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_378),
.A2(n_348),
.B1(n_369),
.B2(n_350),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_413),
.B1(n_372),
.B2(n_387),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_350),
.C(n_362),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_305),
.Y(n_412)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_386),
.A2(n_370),
.B1(n_346),
.B2(n_349),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_342),
.C(n_356),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_377),
.A2(n_355),
.B1(n_352),
.B2(n_346),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_415),
.A2(n_418),
.B1(n_420),
.B2(n_375),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_305),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_392),
.A2(n_391),
.B1(n_396),
.B2(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_372),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_424),
.B(n_436),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_432),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_428),
.C(n_431),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_388),
.Y(n_428)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_408),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_406),
.A2(n_375),
.B1(n_380),
.B2(n_394),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_410),
.A2(n_380),
.B1(n_397),
.B2(n_393),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_413),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_341),
.C(n_342),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_414),
.C(n_400),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_381),
.B1(n_393),
.B2(n_397),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_438),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_402),
.B(n_381),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_409),
.B(n_416),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_430),
.B(n_421),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_398),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_399),
.C(n_411),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_445),
.B(n_423),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_409),
.B(n_419),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_447),
.A2(n_450),
.B(n_451),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_329),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_449),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_341),
.C(n_334),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_425),
.A2(n_334),
.B(n_433),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_421),
.C(n_422),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_454),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_449),
.B(n_422),
.C(n_431),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_458),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_428),
.C(n_427),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_454),
.C(n_455),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_432),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_450),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_457),
.A2(n_453),
.B(n_452),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_465),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_467),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_447),
.B(n_441),
.Y(n_467)
);

OA21x2_ASAP7_75t_SL g468 ( 
.A1(n_462),
.A2(n_461),
.B(n_439),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_463),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_440),
.C(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_470),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_469),
.B(n_471),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_474),
.B(n_475),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_472),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_476),
.B(n_470),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_440),
.Y(n_478)
);


endmodule