module fake_jpeg_8690_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_24),
.B1(n_18),
.B2(n_23),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_22),
.B1(n_31),
.B2(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_35),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.C(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_16),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_67),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_74),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_31),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_25),
.B(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_25),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_72),
.B1(n_25),
.B2(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_22),
.B1(n_31),
.B2(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_31),
.B1(n_19),
.B2(n_27),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_57),
.B1(n_54),
.B2(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_87),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_69),
.C(n_63),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_73),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_43),
.C(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_79),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_79),
.B1(n_73),
.B2(n_63),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_113),
.B1(n_111),
.B2(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_40),
.C(n_37),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_11),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_7),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_98),
.B1(n_91),
.B2(n_82),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_107),
.B(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_81),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.C(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_80),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_97),
.Y(n_123)
);

OAI322xp33_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_100),
.A3(n_103),
.B1(n_107),
.B2(n_28),
.C1(n_9),
.C2(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_98),
.B1(n_84),
.B2(n_17),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_34),
.C(n_28),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_14),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_53),
.B1(n_68),
.B2(n_17),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_117),
.B1(n_127),
.B2(n_120),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_132),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_40),
.CI(n_37),
.CON(n_135),
.SN(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_142),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_126),
.C(n_116),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_118),
.C(n_119),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_145),
.C(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_68),
.C(n_53),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_28),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_156),
.Y(n_163)
);

AOI31xp67_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_135),
.A3(n_138),
.B(n_142),
.Y(n_154)
);

NAND4xp25_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_158),
.C(n_17),
.D(n_9),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_139),
.B1(n_137),
.B2(n_133),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_135),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_17),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_139),
.C(n_133),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_160),
.C(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.C(n_165),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_R g170 ( 
.A(n_164),
.B(n_3),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_1),
.C(n_2),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_157),
.C(n_158),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_163),
.B(n_3),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_168),
.B(n_4),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_1),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_4),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_4),
.C(n_5),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g172 ( 
.A(n_169),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_173),
.B(n_5),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_5),
.Y(n_177)
);


endmodule