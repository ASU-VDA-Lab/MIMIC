module fake_jpeg_5289_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_14),
.C(n_1),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_58),
.B1(n_39),
.B2(n_18),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_27),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_42),
.B(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_75),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_61),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_33),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_50),
.B1(n_59),
.B2(n_49),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_43),
.B1(n_51),
.B2(n_34),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_60),
.B(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_60),
.B1(n_45),
.B2(n_54),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_68),
.A3(n_77),
.B1(n_79),
.B2(n_76),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_98),
.B(n_70),
.C(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_92),
.B1(n_96),
.B2(n_107),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_106),
.B(n_17),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_54),
.B1(n_43),
.B2(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_34),
.B1(n_57),
.B2(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_44),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_84),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_33),
.B1(n_64),
.B2(n_31),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_64),
.B1(n_66),
.B2(n_20),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_68),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_73),
.C(n_70),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_28),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_16),
.B1(n_30),
.B2(n_25),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_19),
.B(n_16),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_110),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_117),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_127),
.B1(n_84),
.B2(n_15),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_106),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_123),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_97),
.B(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_93),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_85),
.C(n_83),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_17),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_129),
.B(n_100),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_75),
.B(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_64),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_92),
.B1(n_98),
.B2(n_89),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_130),
.B1(n_122),
.B2(n_116),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_141),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_136),
.C(n_142),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_137),
.B(n_145),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_129),
.A2(n_105),
.B(n_64),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_91),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_17),
.B(n_18),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_119),
.B1(n_118),
.B2(n_112),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_109),
.B1(n_118),
.B2(n_120),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_167),
.B1(n_169),
.B2(n_143),
.Y(n_176)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_115),
.C(n_117),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_162),
.C(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_145),
.B1(n_137),
.B2(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_118),
.C(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_93),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_149),
.B(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_66),
.C(n_30),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_131),
.B1(n_140),
.B2(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_182),
.B1(n_170),
.B2(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_136),
.C(n_135),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_135),
.B1(n_20),
.B2(n_25),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_1),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_2),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_3),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_161),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_181),
.B(n_155),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_200),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_171),
.B1(n_167),
.B2(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_173),
.B1(n_154),
.B2(n_188),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_183),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_164),
.B(n_158),
.C(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_193),
.B1(n_199),
.B2(n_178),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_206),
.B1(n_212),
.B2(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_179),
.Y(n_211)
);

OAI21x1_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_4),
.B(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_192),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_206),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_202),
.C(n_194),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_4),
.CI(n_5),
.CON(n_229),
.SN(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_196),
.C(n_24),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_24),
.B(n_22),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_228),
.B(n_22),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_4),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_230),
.A3(n_22),
.B1(n_19),
.B2(n_8),
.C1(n_9),
.C2(n_6),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_223),
.B1(n_222),
.B2(n_226),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_12),
.C1(n_13),
.C2(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_233),
.B1(n_19),
.B2(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_6),
.B1(n_9),
.B2(n_12),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_12),
.Y(n_238)
);


endmodule