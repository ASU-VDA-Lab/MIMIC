module real_jpeg_18845_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_0),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_0),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_1),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_53),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_53),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_21),
.B1(n_100),
.B2(n_104),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_4),
.B(n_184),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_196),
.A3(n_199),
.B1(n_202),
.B2(n_206),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_4),
.B(n_121),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_4),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_4),
.B(n_26),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_114),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_8),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_191),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_189),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_163),
.Y(n_12)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_13),
.B(n_163),
.Y(n_190)
);

XOR2x1_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_56),
.B1(n_108),
.B2(n_109),
.Y(n_14)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_37),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_18),
.B(n_38),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_21),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_R g156 ( 
.A(n_21),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_21),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_26),
.B(n_50),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_26),
.B(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_37),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_50),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_38),
.B(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_42),
.Y(n_176)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_49),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_82),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_57),
.A2(n_82),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_65),
.A3(n_68),
.B1(n_74),
.B2(n_80),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_119),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_80),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_88),
.B(n_98),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_85),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_89),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_89),
.B(n_150),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_97),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_98),
.A2(n_217),
.B(n_219),
.Y(n_216)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_142),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_128),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_121),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_121),
.B(n_129),
.Y(n_178)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_156),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_145),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_146),
.B(n_219),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.C(n_186),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_164),
.A2(n_165),
.B1(n_177),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_186),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_261),
.B(n_267),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_234),
.B(n_260),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_215),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_194),
.B(n_215),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_213),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_213),
.Y(n_258)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_228),
.Y(n_215)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_232),
.C(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_253),
.B(n_259),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_249),
.B(n_252),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_258),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);


endmodule