module fake_ibex_1724_n_1268 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_224, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_228, n_1268);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1268;

wire n_1084;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_242;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_1155;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_230;
wire n_917;
wire n_968;
wire n_1253;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_234;
wire n_973;
wire n_1038;
wire n_618;
wire n_662;
wire n_979;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_241;
wire n_231;
wire n_657;
wire n_1156;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1129;
wire n_1244;
wire n_449;
wire n_421;
wire n_738;
wire n_1217;
wire n_236;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1115;
wire n_998;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_996;
wire n_915;
wire n_1174;
wire n_542;
wire n_900;
wire n_377;
wire n_647;
wire n_317;
wire n_326;
wire n_270;
wire n_259;
wire n_339;
wire n_276;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_571;
wire n_229;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_277;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_237;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_302;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_232;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_239;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_243;
wire n_632;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_987;
wire n_750;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_238;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_233;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1016;
wire n_240;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_565;
wire n_1123;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_136),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_28),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_134),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_120),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_57),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_112),
.B(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_107),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_24),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_126),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_131),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_175),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_119),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_73),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_5),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_154),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_122),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_201),
.Y(n_253)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_189),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_92),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_90),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_108),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_168),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_203),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_37),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_57),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_106),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_170),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_160),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_143),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_207),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_118),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_R g284 ( 
.A(n_186),
.B(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_148),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_216),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_166),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_151),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_103),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_198),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_191),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_155),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_169),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_200),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_75),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_0),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_52),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_156),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_145),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_213),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_87),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_27),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_130),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_146),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_144),
.B(n_109),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_125),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_164),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_174),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_78),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_196),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_123),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_138),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_49),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_1),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_197),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_184),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_34),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_153),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_195),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_225),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_141),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_215),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_140),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_121),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_135),
.B(n_167),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_25),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_6),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_66),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_124),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_127),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_51),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_8),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_165),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_180),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_27),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_38),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_178),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_12),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_217),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_0),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_32),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_31),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_90),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_24),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_220),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_107),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_71),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_111),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_101),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_54),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_183),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_105),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_133),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_161),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_74),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_43),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_45),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_30),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_92),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_58),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_149),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_74),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_163),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_137),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_209),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_206),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_79),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_59),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_142),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_51),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_212),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_99),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_89),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_96),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_75),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_97),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_104),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_85),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_199),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_228),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_22),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_50),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_139),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_89),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_28),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_152),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_72),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_150),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_238),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_257),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_238),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_246),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_257),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_361),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_281),
.B(n_2),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_245),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_4),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_247),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_230),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_230),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_294),
.B(n_6),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g421 ( 
.A(n_300),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_258),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_294),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_258),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_309),
.B(n_7),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_273),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_229),
.B(n_8),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_300),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_298),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_245),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_308),
.A2(n_113),
.B(n_110),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_314),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_284),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_296),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_314),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_320),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_320),
.A2(n_115),
.B(n_114),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_324),
.B(n_9),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_330),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_331),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_9),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_344),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_249),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_348),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_350),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_249),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_11),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_256),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_381),
.A2(n_117),
.B(n_116),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_256),
.B(n_15),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_241),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_264),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_264),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_234),
.B(n_15),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_236),
.B(n_237),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_250),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_235),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_244),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_270),
.B(n_16),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_345),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_350),
.B(n_17),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_251),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_270),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_250),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_350),
.B(n_18),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_262),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_252),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_261),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_267),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_467),
.B(n_268),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_311),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_423),
.B(n_231),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_467),
.B(n_269),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_421),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_475),
.B(n_277),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_449),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_410),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_311),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_427),
.B(n_472),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_325),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_410),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_475),
.B(n_278),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_471),
.A2(n_266),
.B1(n_272),
.B2(n_259),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_404),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_455),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_471),
.A2(n_455),
.B1(n_416),
.B2(n_427),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_253),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_485),
.B(n_280),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_408),
.B(n_451),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_408),
.B(n_355),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_451),
.A2(n_232),
.B1(n_248),
.B2(n_239),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_254),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_481),
.B(n_468),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_481),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_417),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_L g538 ( 
.A1(n_413),
.A2(n_362),
.B1(n_367),
.B2(n_355),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_468),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_407),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_425),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_477),
.B(n_253),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_414),
.B(n_283),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_484),
.B(n_285),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_484),
.B(n_287),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_430),
.B(n_372),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_430),
.B(n_372),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_478),
.A2(n_292),
.B1(n_301),
.B2(n_299),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_429),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_414),
.B(n_260),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_453),
.B(n_384),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_434),
.B(n_375),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_460),
.B(n_377),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_474),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_482),
.B(n_313),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_486),
.B(n_289),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_443),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_437),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_479),
.B(n_384),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_439),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_438),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_440),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_466),
.B(n_291),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_415),
.A2(n_302),
.B1(n_303),
.B2(n_271),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_440),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_480),
.B(n_463),
.Y(n_579)
);

OA22x2_ASAP7_75t_L g580 ( 
.A1(n_413),
.A2(n_383),
.B1(n_400),
.B2(n_382),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_450),
.B(n_400),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_440),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_409),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_L g584 ( 
.A1(n_454),
.A2(n_302),
.B1(n_303),
.B2(n_271),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_474),
.A2(n_476),
.B1(n_420),
.B2(n_454),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_409),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_474),
.A2(n_232),
.B1(n_248),
.B2(n_239),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_466),
.B(n_304),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_456),
.B(n_310),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_418),
.B(n_388),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_422),
.A2(n_263),
.B1(n_275),
.B2(n_255),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_422),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_456),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_432),
.A2(n_328),
.B1(n_353),
.B2(n_332),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_585),
.A2(n_263),
.B1(n_275),
.B2(n_255),
.Y(n_598)
);

AND2x6_ASAP7_75t_SL g599 ( 
.A(n_579),
.B(n_531),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_459),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_509),
.Y(n_601)
);

CKINVDCx11_ASAP7_75t_R g602 ( 
.A(n_540),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_531),
.B(n_286),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_595),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_532),
.B(n_419),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_567),
.A2(n_516),
.B1(n_547),
.B2(n_559),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_493),
.B(n_363),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_581),
.B(n_570),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_366),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_526),
.B(n_365),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_380),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_535),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_595),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_552),
.B(n_424),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_504),
.A2(n_522),
.B1(n_503),
.B2(n_507),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_539),
.B(n_527),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_504),
.A2(n_441),
.B1(n_444),
.B2(n_433),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_522),
.A2(n_448),
.B1(n_457),
.B2(n_445),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_512),
.B(n_431),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_520),
.A2(n_295),
.B1(n_297),
.B2(n_286),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_431),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_538),
.B(n_584),
.C(n_577),
.Y(n_624)
);

BUFx6f_ASAP7_75t_SL g625 ( 
.A(n_531),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_564),
.B(n_435),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_583),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_590),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_592),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_SL g630 ( 
.A(n_563),
.B(n_555),
.C(n_515),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_518),
.A2(n_461),
.B1(n_465),
.B2(n_458),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_315),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_556),
.B(n_242),
.C(n_233),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_554),
.B(n_560),
.Y(n_635)
);

BUFx8_ASAP7_75t_L g636 ( 
.A(n_565),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_547),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_547),
.A2(n_356),
.B1(n_364),
.B2(n_359),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_561),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_243),
.Y(n_641)
);

BUFx4_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_530),
.A2(n_312),
.B1(n_357),
.B2(n_305),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_591),
.B(n_274),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_562),
.B(n_569),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_559),
.B(n_279),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_495),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_487),
.B(n_373),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_545),
.C(n_523),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_579),
.A2(n_297),
.B1(n_307),
.B2(n_295),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_531),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_533),
.B(n_316),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_494),
.B(n_318),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_579),
.A2(n_322),
.B1(n_327),
.B2(n_307),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_R g656 ( 
.A(n_573),
.B(n_322),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_596),
.B(n_290),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_579),
.A2(n_336),
.B1(n_398),
.B2(n_327),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_498),
.A2(n_462),
.B(n_442),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_501),
.B(n_293),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_580),
.A2(n_385),
.B1(n_389),
.B2(n_374),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_580),
.A2(n_393),
.B1(n_399),
.B2(n_391),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_514),
.B(n_319),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_543),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_498),
.A2(n_462),
.B(n_442),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_541),
.A2(n_398),
.B1(n_336),
.B2(n_288),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_542),
.A2(n_525),
.B1(n_558),
.B2(n_557),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_578),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_306),
.Y(n_671)
);

AND2x6_ASAP7_75t_SL g672 ( 
.A(n_523),
.B(n_305),
.Y(n_672)
);

INVx8_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_489),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_576),
.B(n_333),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_568),
.B(n_334),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_572),
.B(n_335),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_576),
.B(n_337),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_491),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_575),
.B(n_582),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_549),
.B(n_349),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_589),
.Y(n_682)
);

AND2x6_ASAP7_75t_SL g683 ( 
.A(n_589),
.B(n_312),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_491),
.B(n_352),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_499),
.B(n_386),
.Y(n_685)
);

INVxp33_ASAP7_75t_SL g686 ( 
.A(n_550),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_566),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_499),
.B(n_338),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_499),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_499),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_529),
.B(n_329),
.C(n_321),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_488),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_536),
.B(n_339),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_492),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_574),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_571),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_369),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_497),
.B(n_265),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_500),
.Y(n_699)
);

AND2x6_ASAP7_75t_SL g700 ( 
.A(n_505),
.B(n_357),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_508),
.B(n_276),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_511),
.B(n_282),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_513),
.B(n_378),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_517),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_519),
.B(n_379),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_524),
.B(n_341),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_635),
.B(n_342),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_600),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_624),
.A2(n_358),
.B1(n_401),
.B2(n_395),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_636),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_629),
.B(n_343),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_615),
.B(n_346),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_617),
.B(n_358),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_615),
.B(n_347),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_597),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_623),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_605),
.A2(n_403),
.B(n_317),
.C(n_340),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_626),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_639),
.B(n_351),
.Y(n_720)
);

BUFx8_ASAP7_75t_L g721 ( 
.A(n_625),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_646),
.B(n_387),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_636),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_666),
.B(n_20),
.Y(n_724)
);

OAI21xp33_ASAP7_75t_L g725 ( 
.A1(n_616),
.A2(n_397),
.B(n_534),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_597),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_638),
.A2(n_262),
.B1(n_452),
.B2(n_447),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_673),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_624),
.A2(n_452),
.B1(n_469),
.B2(n_240),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_650),
.A2(n_469),
.B1(n_546),
.B2(n_537),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_654),
.A2(n_551),
.B(n_553),
.C(n_548),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_22),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_648),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_610),
.B(n_23),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_601),
.B(n_23),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_652),
.B(n_606),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_622),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_695),
.B(n_620),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_630),
.B(n_26),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_603),
.B(n_26),
.Y(n_740)
);

BUFx4f_ASAP7_75t_L g741 ( 
.A(n_603),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_612),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_604),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_613),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_633),
.B(n_30),
.Y(n_745)
);

CKINVDCx10_ASAP7_75t_R g746 ( 
.A(n_642),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_621),
.A2(n_611),
.B(n_609),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_686),
.Y(n_749)
);

BUFx4f_ASAP7_75t_L g750 ( 
.A(n_649),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_33),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_655),
.B(n_35),
.Y(n_752)
);

AO21x1_ASAP7_75t_L g753 ( 
.A1(n_653),
.A2(n_588),
.B(n_483),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_598),
.A2(n_658),
.B1(n_662),
.B2(n_661),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_654),
.A2(n_483),
.B(n_37),
.C(n_38),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_687),
.B(n_483),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_676),
.A2(n_677),
.B(n_644),
.Y(n_757)
);

AO32x2_ASAP7_75t_L g758 ( 
.A1(n_668),
.A2(n_39),
.A3(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_662),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_663),
.B(n_46),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_696),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_602),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_599),
.B(n_47),
.Y(n_763)
);

INVx6_ASAP7_75t_L g764 ( 
.A(n_700),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

OR2x6_ASAP7_75t_SL g766 ( 
.A(n_656),
.B(n_48),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_647),
.B(n_50),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_628),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_631),
.B(n_52),
.Y(n_769)
);

BUFx4f_ASAP7_75t_L g770 ( 
.A(n_649),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_675),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_614),
.B(n_56),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_656),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_657),
.B(n_56),
.Y(n_774)
);

BUFx2_ASAP7_75t_SL g775 ( 
.A(n_695),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_697),
.A2(n_706),
.B(n_703),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_683),
.B(n_59),
.Y(n_777)
);

AO21x1_ASAP7_75t_L g778 ( 
.A1(n_697),
.A2(n_60),
.B(n_61),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_641),
.B(n_60),
.Y(n_779)
);

BUFx8_ASAP7_75t_SL g780 ( 
.A(n_672),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_618),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_678),
.B(n_62),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_634),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_693),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_634),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_660),
.B(n_70),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_618),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_693),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_619),
.B(n_76),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_682),
.B(n_77),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_619),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_645),
.B(n_77),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_640),
.Y(n_793)
);

INVx3_ASAP7_75t_SL g794 ( 
.A(n_696),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_679),
.B(n_80),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_664),
.A2(n_129),
.B(n_188),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_667),
.A2(n_128),
.B(n_187),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_669),
.A2(n_227),
.B(n_185),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_671),
.B(n_81),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_670),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_681),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_698),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_707),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_692),
.A2(n_181),
.B(n_179),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_699),
.A2(n_701),
.B(n_702),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_688),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_674),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_689),
.A2(n_91),
.B(n_93),
.C(n_94),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_684),
.B(n_685),
.C(n_690),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_694),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_748),
.B(n_704),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_810),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_711),
.B(n_705),
.Y(n_813)
);

BUFx4f_ASAP7_75t_SL g814 ( 
.A(n_810),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_719),
.B(n_95),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_794),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_SL g817 ( 
.A(n_762),
.B(n_98),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_753),
.A2(n_98),
.A3(n_100),
.B(n_101),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_742),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_714),
.B(n_100),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_728),
.B(n_102),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_710),
.B(n_788),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_765),
.B(n_768),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_733),
.B(n_723),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_754),
.B(n_708),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_778),
.A2(n_739),
.A3(n_731),
.B(n_755),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_767),
.A2(n_786),
.B(n_799),
.C(n_803),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_728),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_722),
.B(n_712),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_802),
.B(n_713),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_790),
.B(n_777),
.Y(n_831)
);

NOR2x1_ASAP7_75t_SL g832 ( 
.A(n_790),
.B(n_775),
.Y(n_832)
);

OAI22x1_ASAP7_75t_L g833 ( 
.A1(n_772),
.A2(n_763),
.B1(n_773),
.B2(n_766),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_728),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_752),
.B(n_741),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_802),
.B(n_715),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_790),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_749),
.B(n_734),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_709),
.A2(n_741),
.B1(n_791),
.B2(n_732),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_777),
.B(n_720),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_R g841 ( 
.A(n_764),
.B(n_743),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_777),
.A2(n_724),
.B1(n_764),
.B2(n_770),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_744),
.Y(n_843)
);

NOR4xp25_ASAP7_75t_L g844 ( 
.A(n_783),
.B(n_785),
.C(n_759),
.D(n_771),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_750),
.B(n_770),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_SL g846 ( 
.A1(n_769),
.A2(n_789),
.B(n_736),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_721),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_772),
.B(n_740),
.Y(n_848)
);

AO31x2_ASAP7_75t_L g849 ( 
.A1(n_806),
.A2(n_784),
.A3(n_808),
.B(n_727),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_751),
.A2(n_774),
.B1(n_787),
.B2(n_781),
.C(n_801),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_738),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_721),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_738),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_792),
.B(n_795),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_795),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_746),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_793),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_779),
.A2(n_725),
.B1(n_760),
.B2(n_782),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_716),
.B(n_726),
.Y(n_860)
);

AO31x2_ASAP7_75t_L g861 ( 
.A1(n_796),
.A2(n_797),
.A3(n_798),
.B(n_804),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_735),
.B(n_780),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_809),
.B(n_761),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_745),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_807),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_758),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_756),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_756),
.B(n_748),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_752),
.B(n_629),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_748),
.B(n_717),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_810),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_728),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_762),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_748),
.B(n_717),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_711),
.B(n_530),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_752),
.B(n_629),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_748),
.B(n_717),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_762),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_748),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_753),
.A2(n_776),
.A3(n_778),
.B(n_739),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_728),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_748),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_728),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_805),
.A2(n_665),
.B(n_659),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_728),
.B(n_748),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_748),
.Y(n_887)
);

AOI221xp5_ASAP7_75t_L g888 ( 
.A1(n_754),
.A2(n_624),
.B1(n_538),
.B2(n_584),
.C(n_661),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_748),
.B(n_717),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_752),
.B(n_629),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_737),
.B(n_556),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_747),
.A2(n_739),
.B(n_635),
.C(n_757),
.Y(n_892)
);

AO31x2_ASAP7_75t_L g893 ( 
.A1(n_753),
.A2(n_776),
.A3(n_778),
.B(n_739),
.Y(n_893)
);

AO22x2_ASAP7_75t_L g894 ( 
.A1(n_754),
.A2(n_651),
.B1(n_622),
.B2(n_530),
.Y(n_894)
);

AO31x2_ASAP7_75t_L g895 ( 
.A1(n_753),
.A2(n_776),
.A3(n_778),
.B(n_739),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_711),
.B(n_723),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_530),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_810),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_718),
.B(n_729),
.C(n_720),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_754),
.A2(n_530),
.B1(n_593),
.B2(n_622),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_748),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_748),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_733),
.B(n_711),
.Y(n_903)
);

INVx3_ASAP7_75t_SL g904 ( 
.A(n_762),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_748),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_747),
.A2(n_739),
.B(n_635),
.C(n_757),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_810),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_748),
.B(n_717),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_810),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_748),
.A2(n_788),
.B1(n_520),
.B2(n_637),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_748),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_728),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_794),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_748),
.B(n_717),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_748),
.B(n_717),
.Y(n_915)
);

OA22x2_ASAP7_75t_L g916 ( 
.A1(n_777),
.A2(n_643),
.B1(n_658),
.B2(n_655),
.Y(n_916)
);

AO21x2_ASAP7_75t_L g917 ( 
.A1(n_753),
.A2(n_730),
.B(n_665),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_748),
.B(n_717),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_748),
.B(n_717),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_794),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_748),
.B(n_717),
.Y(n_921)
);

NOR4xp25_ASAP7_75t_L g922 ( 
.A(n_783),
.B(n_785),
.C(n_754),
.D(n_718),
.Y(n_922)
);

OAI22x1_ASAP7_75t_L g923 ( 
.A1(n_710),
.A2(n_655),
.B1(n_658),
.B2(n_587),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_748),
.B(n_717),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_748),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_714),
.B(n_530),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_762),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_720),
.A2(n_539),
.B(n_629),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_748),
.B(n_717),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_810),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_748),
.B(n_717),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_748),
.B(n_717),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_748),
.B(n_717),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_748),
.B(n_717),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_810),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_711),
.B(n_723),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_754),
.A2(n_530),
.B1(n_593),
.B2(n_622),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_748),
.Y(n_938)
);

NOR2x1_ASAP7_75t_SL g939 ( 
.A(n_790),
.B(n_637),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_753),
.A2(n_730),
.B(n_665),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_748),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_752),
.B(n_629),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_748),
.B(n_717),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_752),
.B(n_629),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_810),
.Y(n_945)
);

AO31x2_ASAP7_75t_L g946 ( 
.A1(n_753),
.A2(n_776),
.A3(n_778),
.B(n_739),
.Y(n_946)
);

AO31x2_ASAP7_75t_L g947 ( 
.A1(n_753),
.A2(n_776),
.A3(n_778),
.B(n_739),
.Y(n_947)
);

AO31x2_ASAP7_75t_L g948 ( 
.A1(n_866),
.A2(n_867),
.A3(n_906),
.B(n_892),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_882),
.B(n_873),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_885),
.Y(n_950)
);

NAND2x1p5_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_873),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_882),
.Y(n_952)
);

OAI21x1_ASAP7_75t_SL g953 ( 
.A1(n_939),
.A2(n_832),
.B(n_837),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_814),
.Y(n_954)
);

OAI21x1_ASAP7_75t_SL g955 ( 
.A1(n_837),
.A2(n_855),
.B(n_839),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_833),
.B(n_935),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_854),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_838),
.A2(n_825),
.B(n_827),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_812),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_897),
.B(n_926),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_871),
.B(n_875),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_910),
.A2(n_899),
.B(n_836),
.Y(n_962)
);

INVx8_ASAP7_75t_L g963 ( 
.A(n_886),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_900),
.A2(n_937),
.B1(n_822),
.B2(n_894),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_888),
.B(n_908),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_915),
.B(n_918),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_929),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_894),
.A2(n_916),
.B1(n_831),
.B2(n_923),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_831),
.A2(n_942),
.B1(n_877),
.B2(n_870),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_872),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_880),
.B(n_887),
.Y(n_971)
);

INVx3_ASAP7_75t_SL g972 ( 
.A(n_852),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_901),
.Y(n_973)
);

OAI21x1_ASAP7_75t_SL g974 ( 
.A1(n_869),
.A2(n_889),
.B(n_878),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_830),
.A2(n_922),
.B(n_844),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_914),
.B(n_919),
.Y(n_976)
);

BUFx2_ASAP7_75t_R g977 ( 
.A(n_904),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_921),
.B(n_924),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_898),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_931),
.B(n_932),
.Y(n_980)
);

AO21x2_ASAP7_75t_L g981 ( 
.A1(n_917),
.A2(n_940),
.B(n_858),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_890),
.B(n_944),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_902),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_884),
.B(n_834),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_933),
.B(n_934),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_902),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_907),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_846),
.B(n_868),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_943),
.B(n_905),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_816),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_891),
.B(n_829),
.Y(n_991)
);

BUFx2_ASAP7_75t_SL g992 ( 
.A(n_909),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_864),
.A2(n_857),
.B(n_819),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_911),
.B(n_925),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_911),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_851),
.A2(n_853),
.B(n_843),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_925),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_945),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_850),
.A2(n_815),
.B(n_823),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_SL g1000 ( 
.A1(n_938),
.A2(n_941),
.B(n_821),
.Y(n_1000)
);

OA21x2_ASAP7_75t_L g1001 ( 
.A1(n_863),
.A2(n_947),
.B(n_946),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_913),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_811),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_845),
.B(n_884),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_920),
.B(n_860),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_848),
.B(n_835),
.Y(n_1006)
);

CKINVDCx11_ASAP7_75t_R g1007 ( 
.A(n_874),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_859),
.B(n_840),
.Y(n_1008)
);

AO21x2_ASAP7_75t_L g1009 ( 
.A1(n_881),
.A2(n_947),
.B(n_946),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_865),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

AO31x2_ASAP7_75t_L g1012 ( 
.A1(n_881),
.A2(n_893),
.A3(n_895),
.B(n_826),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_928),
.B(n_876),
.C(n_842),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_828),
.A2(n_912),
.B(n_895),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_930),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_893),
.A2(n_826),
.B(n_818),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_886),
.B(n_813),
.Y(n_1017)
);

OA21x2_ASAP7_75t_L g1018 ( 
.A1(n_861),
.A2(n_849),
.B(n_862),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_824),
.A2(n_903),
.B(n_849),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_813),
.A2(n_936),
.B(n_896),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_841),
.A2(n_817),
.B(n_936),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_896),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_847),
.A2(n_856),
.B(n_874),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_879),
.Y(n_1024)
);

INVx3_ASAP7_75t_SL g1025 ( 
.A(n_879),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_927),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_883),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_897),
.B(n_530),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_882),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_R g1030 ( 
.A(n_812),
.B(n_762),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_837),
.B(n_855),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_894),
.A2(n_752),
.B1(n_916),
.B2(n_888),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_816),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_866),
.A2(n_867),
.A3(n_906),
.B(n_892),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_894),
.A2(n_752),
.B1(n_916),
.B2(n_888),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_814),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_882),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_886),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_897),
.B(n_926),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_883),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_837),
.B(n_530),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_983),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_963),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_963),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_961),
.B(n_980),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_983),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1031),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_971),
.B(n_986),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_963),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_995),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_950),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_992),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_971),
.B(n_997),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_985),
.B(n_976),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_973),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_971),
.B(n_994),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_1017),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1039),
.B(n_978),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_958),
.B(n_975),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_949),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_993),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_954),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_965),
.B(n_989),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1014),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1039),
.B(n_991),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_948),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1032),
.A2(n_1035),
.B1(n_968),
.B2(n_991),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_968),
.B(n_964),
.Y(n_1068)
);

BUFx2_ASAP7_75t_SL g1069 ( 
.A(n_1017),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_951),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1031),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1034),
.Y(n_1072)
);

BUFx10_ASAP7_75t_L g1073 ( 
.A(n_954),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1010),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1038),
.B(n_996),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_966),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1034),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1034),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1034),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_952),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1018),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_1047),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1045),
.B(n_1015),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1056),
.B(n_1018),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1068),
.A2(n_1035),
.B1(n_1032),
.B2(n_1013),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1045),
.B(n_1015),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1042),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1056),
.B(n_1001),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1059),
.B(n_1063),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1059),
.B(n_1001),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1068),
.B(n_1054),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1042),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1075),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1051),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1054),
.B(n_1012),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1046),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1048),
.B(n_1016),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1048),
.B(n_1016),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1052),
.B(n_1020),
.C(n_990),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1053),
.B(n_1009),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1080),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1053),
.B(n_1009),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1067),
.A2(n_1041),
.B1(n_999),
.B2(n_982),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_1073),
.Y(n_1105)
);

BUFx2_ASAP7_75t_SL g1106 ( 
.A(n_1060),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1047),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1070),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_1050),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1065),
.A2(n_1028),
.B1(n_982),
.B2(n_957),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1071),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1061),
.A2(n_974),
.B(n_988),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1055),
.B(n_981),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1082),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1095),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1094),
.B(n_1064),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1088),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_1095),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1088),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1093),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1090),
.B(n_1066),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1090),
.B(n_1072),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1089),
.B(n_1077),
.Y(n_1123)
);

NAND2x1_ASAP7_75t_L g1124 ( 
.A(n_1107),
.B(n_1071),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1089),
.B(n_1078),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1082),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1085),
.B(n_1079),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1085),
.B(n_1081),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1091),
.B(n_1101),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1097),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1091),
.B(n_1101),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1109),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1094),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1103),
.B(n_1081),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1129),
.B(n_1096),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1117),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_1118),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1129),
.B(n_1103),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1117),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1118),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1119),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1119),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1116),
.B(n_1094),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1130),
.A2(n_1104),
.B(n_1102),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1115),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1131),
.B(n_1098),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1131),
.B(n_1098),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1114),
.B(n_1107),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1134),
.B(n_1113),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_SL g1150 ( 
.A(n_1114),
.B(n_1106),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1124),
.B(n_1107),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1116),
.B(n_1094),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1128),
.B(n_1099),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1128),
.B(n_1099),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_1115),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1120),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1154),
.B(n_1105),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1150),
.A2(n_1100),
.B(n_956),
.Y(n_1158)
);

OAI322xp33_ASAP7_75t_L g1159 ( 
.A1(n_1135),
.A2(n_1092),
.A3(n_1084),
.B1(n_1087),
.B2(n_1121),
.C1(n_1122),
.C2(n_1110),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1136),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1150),
.B(n_1105),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1153),
.B(n_1127),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1136),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1139),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1151),
.A2(n_1126),
.B(n_1114),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1138),
.B(n_1123),
.Y(n_1166)
);

AOI31xp33_ASAP7_75t_L g1167 ( 
.A1(n_1148),
.A2(n_1100),
.A3(n_1030),
.B(n_1074),
.Y(n_1167)
);

OAI31xp33_ASAP7_75t_L g1168 ( 
.A1(n_1148),
.A2(n_1086),
.A3(n_1108),
.B(n_1082),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1139),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1154),
.B(n_1135),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1138),
.B(n_1123),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1141),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1151),
.A2(n_1124),
.B(n_1112),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1141),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1142),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1146),
.B(n_1125),
.Y(n_1176)
);

OAI211xp5_ASAP7_75t_L g1177 ( 
.A1(n_1144),
.A2(n_998),
.B(n_979),
.C(n_1110),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1146),
.B(n_1125),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1142),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1168),
.B(n_1145),
.C(n_1144),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1167),
.A2(n_1151),
.B(n_1148),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1170),
.Y(n_1182)
);

AOI222xp33_ASAP7_75t_L g1183 ( 
.A1(n_1165),
.A2(n_1140),
.B1(n_1137),
.B2(n_1155),
.C1(n_1147),
.C2(n_1153),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1170),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1160),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1160),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1166),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1161),
.A2(n_1151),
.B1(n_1126),
.B2(n_1114),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1163),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1163),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1159),
.B(n_1155),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1164),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_1177),
.A2(n_1021),
.B(n_1022),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1164),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_1158),
.A2(n_1021),
.B(n_1022),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1175),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1157),
.A2(n_1092),
.B1(n_1151),
.B2(n_969),
.C(n_1149),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1166),
.B(n_1147),
.Y(n_1198)
);

OAI32xp33_ASAP7_75t_L g1199 ( 
.A1(n_1162),
.A2(n_1126),
.A3(n_1107),
.B1(n_1108),
.B2(n_1102),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1175),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1171),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1191),
.A2(n_1176),
.B1(n_1178),
.B2(n_1171),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1191),
.A2(n_1178),
.B(n_1176),
.Y(n_1203)
);

XOR2x2_ASAP7_75t_L g1204 ( 
.A(n_1181),
.B(n_972),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1183),
.A2(n_1173),
.B(n_1149),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1201),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1180),
.A2(n_1143),
.B1(n_1152),
.B2(n_1127),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1182),
.B(n_1140),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1185),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1197),
.B(n_1179),
.C(n_1172),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1184),
.B(n_1179),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1193),
.A2(n_1174),
.B(n_1169),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1203),
.A2(n_1188),
.B1(n_1187),
.B2(n_1195),
.Y(n_1213)
);

OAI211xp5_ASAP7_75t_L g1214 ( 
.A1(n_1207),
.A2(n_1007),
.B(n_1036),
.C(n_1199),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1211),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1205),
.A2(n_1210),
.B1(n_1202),
.B2(n_1206),
.C(n_1209),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1204),
.B(n_1187),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1208),
.A2(n_1200),
.B(n_1189),
.Y(n_1218)
);

OA22x2_ASAP7_75t_L g1219 ( 
.A1(n_1212),
.A2(n_1198),
.B1(n_1106),
.B2(n_972),
.Y(n_1219)
);

OAI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_1212),
.A2(n_1186),
.B1(n_1192),
.B2(n_1196),
.C(n_1194),
.Y(n_1220)
);

AND5x1_ASAP7_75t_L g1221 ( 
.A(n_1202),
.B(n_977),
.C(n_1188),
.D(n_1007),
.E(n_1112),
.Y(n_1221)
);

AOI211xp5_ASAP7_75t_L g1222 ( 
.A1(n_1203),
.A2(n_1199),
.B(n_1025),
.C(n_1026),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1202),
.B(n_1190),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1203),
.A2(n_1190),
.B1(n_1002),
.B2(n_1033),
.C(n_1024),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1204),
.A2(n_988),
.B(n_1019),
.Y(n_1225)
);

NAND4xp75_ASAP7_75t_L g1226 ( 
.A(n_1216),
.B(n_959),
.C(n_970),
.D(n_1044),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1215),
.B(n_1156),
.Y(n_1227)
);

NAND4xp75_ASAP7_75t_L g1228 ( 
.A(n_1217),
.B(n_1044),
.C(n_1049),
.D(n_1000),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1220),
.A2(n_998),
.B1(n_979),
.B2(n_1156),
.C(n_987),
.Y(n_1229)
);

NAND5xp2_ASAP7_75t_L g1230 ( 
.A(n_1214),
.B(n_1023),
.C(n_969),
.D(n_962),
.E(n_1025),
.Y(n_1230)
);

AOI211xp5_ASAP7_75t_L g1231 ( 
.A1(n_1225),
.A2(n_987),
.B(n_1062),
.C(n_960),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1224),
.A2(n_1143),
.B1(n_1152),
.B2(n_1133),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_L g1233 ( 
.A(n_1222),
.B(n_1062),
.C(n_1011),
.Y(n_1233)
);

NAND4xp25_ASAP7_75t_L g1234 ( 
.A(n_1213),
.B(n_1058),
.C(n_1108),
.D(n_1126),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1219),
.A2(n_1111),
.B1(n_1083),
.B2(n_1132),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1233),
.B(n_1221),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1229),
.B(n_1218),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_SL g1238 ( 
.A(n_1231),
.B(n_1223),
.C(n_1073),
.Y(n_1238)
);

OR5x1_ASAP7_75t_L g1239 ( 
.A(n_1234),
.B(n_1073),
.C(n_953),
.D(n_1069),
.E(n_1057),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_L g1240 ( 
.A(n_1226),
.B(n_1029),
.C(n_952),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_SL g1241 ( 
.A(n_1230),
.B(n_1006),
.C(n_957),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1228),
.B(n_1143),
.Y(n_1242)
);

NAND4xp75_ASAP7_75t_L g1243 ( 
.A(n_1232),
.B(n_1049),
.C(n_1008),
.D(n_1080),
.Y(n_1243)
);

NOR3xp33_ASAP7_75t_L g1244 ( 
.A(n_1235),
.B(n_1037),
.C(n_1029),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_L g1245 ( 
.A(n_1238),
.B(n_1037),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1237),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1236),
.B(n_1227),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1236),
.B(n_1070),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_R g1249 ( 
.A(n_1242),
.B(n_1005),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1244),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_L g1251 ( 
.A(n_1243),
.B(n_1005),
.C(n_1038),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1241),
.Y(n_1252)
);

OAI221xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1240),
.A2(n_1003),
.B1(n_1076),
.B2(n_1043),
.C(n_967),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1250),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1248),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1252),
.B(n_1239),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1246),
.B(n_1121),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1245),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1255),
.A2(n_1247),
.B1(n_1253),
.B2(n_1251),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1257),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1258),
.B(n_1253),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1259),
.A2(n_1254),
.B(n_1256),
.C(n_1261),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1262),
.B(n_1260),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1262),
.A2(n_1249),
.B(n_1005),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1263),
.A2(n_1004),
.B(n_984),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1265),
.B(n_1264),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1266),
.A2(n_955),
.B(n_1004),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_1004),
.B(n_1040),
.C(n_1027),
.Y(n_1268)
);


endmodule