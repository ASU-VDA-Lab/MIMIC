module fake_aes_4370_n_46 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_25;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_12), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_1), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
INVxp67_ASAP7_75t_SL g20 ( .A(n_11), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_0), .A2(n_5), .B1(n_10), .B2(n_6), .Y(n_21) );
INVx4_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_17), .B(n_1), .C(n_2), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_19), .B(n_3), .Y(n_25) );
NOR3xp33_ASAP7_75t_SL g26 ( .A(n_21), .B(n_3), .C(n_4), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_19), .B(n_6), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_15), .B1(n_18), .B2(n_13), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_15), .B1(n_18), .B2(n_13), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_24), .Y(n_31) );
OAI221xp5_ASAP7_75t_SL g32 ( .A1(n_30), .A2(n_25), .B1(n_13), .B2(n_26), .C(n_19), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_24), .Y(n_33) );
INVxp67_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_35), .Y(n_37) );
HB1xp67_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
O2A1O1Ixp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_32), .B(n_28), .C(n_21), .Y(n_39) );
OAI211xp5_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_23), .B(n_20), .C(n_29), .Y(n_40) );
OAI211xp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_20), .B(n_14), .C(n_22), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_38), .Y(n_42) );
OAI221xp5_ASAP7_75t_L g43 ( .A1(n_40), .A2(n_14), .B1(n_31), .B2(n_22), .C(n_7), .Y(n_43) );
HB1xp67_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
INVx2_ASAP7_75t_L g45 ( .A(n_42), .Y(n_45) );
AOI322xp5_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_7), .A3(n_9), .B1(n_22), .B2(n_41), .C1(n_43), .C2(n_45), .Y(n_46) );
endmodule