module fake_ariane_1202_n_759 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_759);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_759;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_557;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_458;
wire n_361;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_10),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_80),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_14),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_43),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_68),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_54),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_70),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_73),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_47),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_82),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_26),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_52),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_23),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

CKINVDCx11_ASAP7_75t_R g191 ( 
.A(n_53),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_9),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_23),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

BUFx8_ASAP7_75t_SL g198 ( 
.A(n_58),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_6),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_19),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_0),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_0),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_27),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_1),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_28),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_2),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_2),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_3),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_3),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_4),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_4),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_189),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_156),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_153),
.B(n_5),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_151),
.B(n_5),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

NOR2x1p5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_152),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_166),
.B1(n_159),
.B2(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_194),
.B1(n_193),
.B2(n_186),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_179),
.B1(n_177),
.B2(n_174),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_154),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_205),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_165),
.B1(n_171),
.B2(n_169),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_216),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_168),
.B1(n_164),
.B2(n_163),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_241),
.B1(n_236),
.B2(n_225),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_161),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_211),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_178),
.B1(n_161),
.B2(n_9),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_161),
.Y(n_264)
);

CKINVDCx6p67_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_178),
.B1(n_161),
.B2(n_10),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_178),
.B1(n_12),
.B2(n_13),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_178),
.B1(n_12),
.B2(n_13),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_178),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_208),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_224),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_227),
.A2(n_178),
.B1(n_18),
.B2(n_19),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_209),
.B(n_17),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_208),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_279)
);

OR2x6_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_22),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_282)
);

BUFx6f_ASAP7_75t_SL g283 ( 
.A(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

AO22x2_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_35),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_36),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_243),
.B(n_37),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_213),
.B1(n_212),
.B2(n_232),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

XOR2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_212),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_213),
.B(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_210),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

INVx3_ASAP7_75t_R g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

NAND2x1p5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_202),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_248),
.B(n_254),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_239),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_255),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_202),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_244),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_253),
.B(n_239),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_217),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_266),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_244),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_38),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_250),
.B(n_202),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_202),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_259),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_39),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_204),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_271),
.B(n_204),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_278),
.B(n_204),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_267),
.B(n_204),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_245),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_207),
.Y(n_351)
);

XNOR2x2_ASAP7_75t_SL g352 ( 
.A(n_285),
.B(n_210),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_272),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_260),
.B(n_210),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_207),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_358),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_206),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_206),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_210),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_349),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_207),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_207),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_40),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_299),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_215),
.B(n_210),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_294),
.A2(n_215),
.B(n_42),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_304),
.B(n_215),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_215),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_41),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_215),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_45),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_353),
.A2(n_46),
.B(n_48),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_50),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_51),
.B(n_55),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_56),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_57),
.B(n_59),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_323),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_313),
.B(n_60),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_139),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_61),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_317),
.B(n_318),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_138),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_333),
.B(n_63),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_303),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_330),
.B(n_64),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_333),
.B(n_65),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_137),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_335),
.B(n_66),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_310),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_348),
.B(n_340),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_310),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_337),
.B(n_136),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_305),
.B(n_67),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_331),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_417),
.Y(n_430)
);

NAND2x1_ASAP7_75t_SL g431 ( 
.A(n_420),
.B(n_331),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_372),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_298),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_367),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_311),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_376),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_298),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_334),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_385),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_320),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_326),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_349),
.Y(n_458)
);

NAND2x1p5_ASAP7_75t_L g459 ( 
.A(n_360),
.B(n_306),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_71),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_76),
.Y(n_461)
);

BUFx6f_ASAP7_75t_SL g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_421),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_77),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_78),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_81),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_365),
.B(n_83),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_363),
.B(n_84),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_85),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_407),
.B(n_86),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_407),
.B(n_87),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_363),
.B(n_427),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_419),
.B(n_88),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_363),
.B(n_89),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_374),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_411),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_411),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_436),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_436),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_481),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_429),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_419),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_451),
.A2(n_484),
.B1(n_462),
.B2(n_483),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_365),
.Y(n_495)
);

BUFx2_ASAP7_75t_SL g496 ( 
.A(n_437),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_448),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_455),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_464),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_439),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_454),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_474),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_439),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_430),
.B(n_412),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

BUFx8_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_463),
.Y(n_524)
);

CKINVDCx11_ASAP7_75t_R g525 ( 
.A(n_471),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_478),
.Y(n_526)
);

BUFx5_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_412),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_443),
.B1(n_484),
.B2(n_482),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_488),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_529),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_446),
.B1(n_449),
.B2(n_453),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_513),
.A2(n_449),
.B1(n_408),
.B2(n_383),
.Y(n_535)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_486),
.Y(n_536)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_488),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_502),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_525),
.A2(n_446),
.B1(n_471),
.B2(n_468),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_513),
.A2(n_522),
.B1(n_501),
.B2(n_500),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_508),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_509),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_490),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_500),
.A2(n_476),
.B1(n_475),
.B2(n_466),
.Y(n_547)
);

BUFx4f_ASAP7_75t_SL g548 ( 
.A(n_485),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_522),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_500),
.A2(n_479),
.B1(n_441),
.B2(n_396),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_528),
.A2(n_453),
.B1(n_371),
.B2(n_458),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_515),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_490),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_528),
.A2(n_458),
.B1(n_412),
.B2(n_402),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_522),
.A2(n_392),
.B1(n_387),
.B2(n_479),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_525),
.A2(n_395),
.B1(n_379),
.B2(n_384),
.Y(n_560)
);

CKINVDCx11_ASAP7_75t_R g561 ( 
.A(n_485),
.Y(n_561)
);

CKINVDCx6p67_ASAP7_75t_R g562 ( 
.A(n_489),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_504),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_495),
.A2(n_379),
.B1(n_384),
.B2(n_438),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_490),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_500),
.A2(n_523),
.B1(n_512),
.B2(n_510),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_500),
.A2(n_523),
.B1(n_512),
.B2(n_527),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_487),
.B(n_441),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_535),
.A2(n_547),
.B(n_409),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_532),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_539),
.A2(n_494),
.B(n_403),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_559),
.A2(n_512),
.B1(n_523),
.B2(n_496),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_539),
.A2(n_493),
.B1(n_492),
.B2(n_379),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_559),
.A2(n_493),
.B1(n_384),
.B2(n_416),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_550),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_569),
.B(n_516),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_534),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_543),
.B(n_519),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_537),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_542),
.A2(n_403),
.B(n_413),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_533),
.A2(n_493),
.B1(n_401),
.B2(n_392),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_555),
.A2(n_523),
.B1(n_504),
.B2(n_480),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_554),
.A2(n_401),
.B1(n_479),
.B2(n_527),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_486),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_563),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_530),
.A2(n_523),
.B1(n_480),
.B2(n_391),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

OAI222xp33_ASAP7_75t_L g596 ( 
.A1(n_558),
.A2(n_526),
.B1(n_400),
.B2(n_423),
.C1(n_419),
.C2(n_362),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_554),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_542),
.B(n_498),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_560),
.A2(n_401),
.B1(n_527),
.B2(n_400),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_564),
.A2(n_527),
.B1(n_364),
.B2(n_373),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_548),
.B(n_536),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_540),
.B(n_503),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_546),
.A2(n_527),
.B1(n_472),
.B2(n_418),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_546),
.A2(n_527),
.B1(n_472),
.B2(n_393),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_548),
.A2(n_527),
.B1(n_373),
.B2(n_364),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_568),
.A2(n_388),
.B(n_459),
.Y(n_610)
);

OAI21xp33_ASAP7_75t_L g611 ( 
.A1(n_566),
.A2(n_431),
.B(n_406),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_567),
.A2(n_373),
.B1(n_375),
.B2(n_364),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_549),
.Y(n_614)
);

AOI222xp33_ASAP7_75t_L g615 ( 
.A1(n_561),
.A2(n_427),
.B1(n_489),
.B2(n_499),
.C1(n_378),
.C2(n_404),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_544),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_503),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_589),
.A2(n_557),
.B1(n_499),
.B2(n_508),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_581),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_SL g621 ( 
.A(n_615),
.B(n_459),
.C(n_427),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_578),
.B(n_498),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_SL g623 ( 
.A(n_570),
.B(n_405),
.C(n_544),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_574),
.A2(n_398),
.B1(n_423),
.B2(n_399),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_605),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_398),
.B1(n_423),
.B2(n_399),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_572),
.A2(n_508),
.B1(n_562),
.B2(n_557),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_598),
.A2(n_508),
.B1(n_467),
.B2(n_473),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_585),
.B(n_498),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_579),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_595),
.B(n_521),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_584),
.A2(n_391),
.B1(n_426),
.B2(n_511),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_582),
.B(n_505),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_598),
.A2(n_467),
.B1(n_473),
.B2(n_461),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_611),
.A2(n_398),
.B1(n_399),
.B2(n_375),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_590),
.A2(n_575),
.B1(n_607),
.B2(n_588),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_SL g638 ( 
.A1(n_610),
.A2(n_410),
.B1(n_404),
.B2(n_361),
.C(n_359),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_593),
.A2(n_391),
.B1(n_426),
.B2(n_511),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_595),
.B(n_521),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_601),
.A2(n_391),
.B1(n_511),
.B2(n_452),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_594),
.A2(n_461),
.B1(n_375),
.B2(n_521),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_606),
.A2(n_399),
.B1(n_410),
.B2(n_368),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_580),
.B(n_520),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_597),
.A2(n_511),
.B1(n_452),
.B2(n_457),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_613),
.A2(n_505),
.B1(n_520),
.B2(n_518),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_613),
.A2(n_518),
.B1(n_382),
.B2(n_386),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_597),
.B(n_361),
.C(n_399),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_614),
.B(n_591),
.C(n_616),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_573),
.A2(n_442),
.B1(n_428),
.B2(n_450),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_612),
.A2(n_425),
.B(n_432),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_576),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_583),
.A2(n_521),
.B1(n_514),
.B2(n_428),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_609),
.A2(n_477),
.B1(n_457),
.B2(n_452),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_576),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_L g656 ( 
.A1(n_638),
.A2(n_599),
.B(n_616),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_625),
.B(n_599),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_627),
.A2(n_604),
.B(n_618),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_SL g659 ( 
.A(n_623),
.B(n_583),
.C(n_617),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_620),
.B(n_608),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_636),
.A2(n_592),
.B1(n_577),
.B2(n_596),
.C(n_608),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_622),
.B(n_603),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_652),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_649),
.B(n_603),
.C(n_602),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_637),
.B(n_600),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_630),
.B(n_600),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_653),
.B(n_600),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_652),
.B(n_600),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_636),
.A2(n_643),
.B1(n_632),
.B2(n_628),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_600),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_577),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_571),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_633),
.B(n_571),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_631),
.B(n_521),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_640),
.B(n_514),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_643),
.B(n_514),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_514),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_648),
.B(n_397),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_619),
.B(n_440),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_663),
.B(n_634),
.C(n_635),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_650),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_657),
.B(n_621),
.Y(n_682)
);

AOI211xp5_ASAP7_75t_L g683 ( 
.A1(n_669),
.A2(n_642),
.B(n_639),
.C(n_641),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_667),
.B(n_677),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_659),
.B(n_646),
.C(n_651),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_668),
.B(n_654),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_666),
.B(n_672),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_672),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_676),
.A2(n_647),
.B1(n_624),
.B2(n_626),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_676),
.A2(n_399),
.B1(n_642),
.B2(n_397),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_660),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_658),
.B(n_442),
.C(n_440),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_656),
.B(n_477),
.C(n_457),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_691),
.B(n_665),
.Y(n_694)
);

NAND4xp75_ASAP7_75t_SL g695 ( 
.A(n_686),
.B(n_675),
.C(n_679),
.D(n_667),
.Y(n_695)
);

XNOR2x2_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_661),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_688),
.B(n_662),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_687),
.Y(n_698)
);

NAND4xp75_ASAP7_75t_L g699 ( 
.A(n_681),
.B(n_679),
.C(n_673),
.D(n_675),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g700 ( 
.A(n_684),
.B(n_685),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_684),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_684),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_682),
.Y(n_703)
);

XOR2x2_ASAP7_75t_L g704 ( 
.A(n_700),
.B(n_693),
.Y(n_704)
);

XOR2x2_ASAP7_75t_L g705 ( 
.A(n_696),
.B(n_683),
.Y(n_705)
);

NOR2x1_ASAP7_75t_L g706 ( 
.A(n_695),
.B(n_680),
.Y(n_706)
);

OAI22x1_ASAP7_75t_L g707 ( 
.A1(n_702),
.A2(n_664),
.B1(n_671),
.B2(n_683),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_703),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_708),
.Y(n_709)
);

OA22x2_ASAP7_75t_L g710 ( 
.A1(n_707),
.A2(n_703),
.B1(n_701),
.B2(n_698),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_705),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_704),
.Y(n_713)
);

OA22x2_ASAP7_75t_L g714 ( 
.A1(n_712),
.A2(n_701),
.B1(n_697),
.B2(n_695),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_709),
.Y(n_716)
);

OAI322xp33_ASAP7_75t_L g717 ( 
.A1(n_710),
.A2(n_694),
.A3(n_678),
.B1(n_674),
.B2(n_699),
.C1(n_692),
.C2(n_690),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_713),
.B1(n_709),
.B2(n_689),
.Y(n_718)
);

OA22x2_ASAP7_75t_L g719 ( 
.A1(n_715),
.A2(n_716),
.B1(n_717),
.B2(n_432),
.Y(n_719)
);

AO22x1_ASAP7_75t_SL g720 ( 
.A1(n_718),
.A2(n_716),
.B1(n_92),
.B2(n_93),
.Y(n_720)
);

BUFx8_ASAP7_75t_L g721 ( 
.A(n_719),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_SL g722 ( 
.A1(n_718),
.A2(n_470),
.B(n_397),
.C(n_377),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_720),
.Y(n_723)
);

AOI31xp33_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_386),
.A3(n_382),
.B(n_369),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_722),
.B(n_470),
.C(n_369),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_477),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_721),
.B(n_477),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_721),
.A2(n_397),
.B1(n_366),
.B2(n_381),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_720),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_723),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_729),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_457),
.B1(n_452),
.B2(n_96),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_724),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_725),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_728),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

NAND4xp25_ASAP7_75t_L g737 ( 
.A(n_731),
.B(n_727),
.C(n_94),
.D(n_98),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_734),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_732),
.A2(n_366),
.B1(n_381),
.B2(n_101),
.Y(n_739)
);

AOI211xp5_ASAP7_75t_SL g740 ( 
.A1(n_733),
.A2(n_366),
.B(n_381),
.C(n_102),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_735),
.B1(n_366),
.B2(n_381),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_738),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_739),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_737),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_740),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_742),
.B1(n_743),
.B2(n_744),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_741),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_745),
.A2(n_366),
.B1(n_381),
.B2(n_103),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_742),
.A2(n_366),
.B1(n_381),
.B2(n_104),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_366),
.B1(n_381),
.B2(n_105),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_747),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_750),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_752),
.A2(n_746),
.B1(n_748),
.B2(n_749),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_91),
.B1(n_100),
.B2(n_106),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_753),
.Y(n_755)
);

AOI211xp5_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_751),
.B(n_754),
.C(n_109),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_756),
.Y(n_757)
);

AOI221xp5_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.C(n_111),
.Y(n_758)
);

AOI211xp5_ASAP7_75t_L g759 ( 
.A1(n_758),
.A2(n_112),
.B(n_116),
.C(n_119),
.Y(n_759)
);


endmodule