module real_aes_8091_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
NAND3xp33_ASAP7_75t_SL g734 ( .A(n_0), .B(n_83), .C(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g474 ( .A(n_1), .Y(n_474) );
INVx1_ASAP7_75t_L g253 ( .A(n_2), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_3), .A2(n_36), .B1(n_172), .B2(n_502), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g160 ( .A1(n_4), .A2(n_161), .B(n_162), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_5), .B(n_159), .Y(n_451) );
AND2x6_ASAP7_75t_L g134 ( .A(n_6), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_7), .A2(n_229), .B(n_230), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_8), .B(n_37), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_8), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g169 ( .A(n_9), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_10), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g131 ( .A(n_11), .Y(n_131) );
INVx1_ASAP7_75t_L g470 ( .A(n_12), .Y(n_470) );
INVx1_ASAP7_75t_L g235 ( .A(n_13), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_14), .B(n_137), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_15), .B(n_127), .Y(n_479) );
AO32x2_ASAP7_75t_L g499 ( .A1(n_16), .A2(n_126), .A3(n_159), .B1(n_462), .B2(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_17), .B(n_172), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_18), .B(n_180), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_19), .B(n_127), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_20), .A2(n_50), .B1(n_172), .B2(n_502), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_21), .B(n_161), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_22), .A2(n_74), .B1(n_137), .B2(n_172), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_23), .B(n_172), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_24), .B(n_157), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_25), .A2(n_233), .B(n_234), .C(n_236), .Y(n_232) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_26), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_27), .B(n_174), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_28), .B(n_167), .Y(n_254) );
AOI222xp33_ASAP7_75t_L g116 ( .A1(n_29), .A2(n_97), .B1(n_117), .B2(n_718), .C1(n_721), .C2(n_722), .Y(n_116) );
INVx1_ASAP7_75t_L g145 ( .A(n_30), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_31), .B(n_174), .Y(n_496) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_33), .B(n_172), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_34), .B(n_174), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_35), .A2(n_134), .B(n_146), .C(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g733 ( .A(n_37), .Y(n_733) );
INVx1_ASAP7_75t_L g143 ( .A(n_38), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_39), .B(n_167), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_40), .A2(n_118), .B1(n_119), .B2(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_40), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_41), .Y(n_108) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_42), .A2(n_100), .B1(n_730), .B2(n_738), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_43), .B(n_172), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_44), .A2(n_84), .B1(n_197), .B2(n_502), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_45), .B(n_172), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_46), .B(n_172), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_47), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_48), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_49), .B(n_161), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_51), .A2(n_60), .B1(n_137), .B2(n_172), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_52), .A2(n_137), .B1(n_140), .B2(n_146), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_53), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_54), .B(n_172), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_55), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_56), .B(n_172), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_57), .A2(n_166), .B(n_168), .C(n_171), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_58), .Y(n_210) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
INVx1_ASAP7_75t_L g135 ( .A(n_61), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_62), .B(n_172), .Y(n_475) );
INVx1_ASAP7_75t_L g130 ( .A(n_63), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_64), .Y(n_106) );
AO32x2_ASAP7_75t_L g519 ( .A1(n_65), .A2(n_159), .A3(n_215), .B1(n_462), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g459 ( .A(n_66), .Y(n_459) );
INVx1_ASAP7_75t_L g491 ( .A(n_67), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_68), .A2(n_171), .B(n_180), .C(n_181), .Y(n_179) );
INVxp67_ASAP7_75t_L g182 ( .A(n_69), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_70), .B(n_137), .Y(n_492) );
INVx1_ASAP7_75t_L g737 ( .A(n_71), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_72), .Y(n_154) );
INVx1_ASAP7_75t_L g203 ( .A(n_73), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_75), .A2(n_134), .B(n_146), .C(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_76), .B(n_502), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_77), .B(n_137), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_78), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_80), .B(n_180), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_81), .B(n_137), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_82), .A2(n_134), .B(n_146), .C(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g111 ( .A(n_83), .B(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g433 ( .A(n_83), .B(n_113), .Y(n_433) );
INVx2_ASAP7_75t_L g717 ( .A(n_83), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_85), .A2(n_98), .B1(n_137), .B2(n_138), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_86), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_87), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_88), .A2(n_134), .B(n_146), .C(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_89), .Y(n_225) );
INVx1_ASAP7_75t_L g178 ( .A(n_90), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_91), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_92), .B(n_193), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_93), .B(n_137), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_94), .B(n_159), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_95), .A2(n_161), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_96), .B(n_737), .Y(n_736) );
CKINVDCx16_ASAP7_75t_R g721 ( .A(n_97), .Y(n_721) );
BUFx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_106), .B1(n_116), .B2(n_725), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_107), .A2(n_726), .B(n_728), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g729 ( .A(n_111), .Y(n_729) );
NOR2x2_ASAP7_75t_L g724 ( .A(n_112), .B(n_717), .Y(n_724) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g716 ( .A(n_113), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_431), .B1(n_434), .B2(n_714), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_119), .A2(n_431), .B1(n_719), .B2(n_720), .Y(n_718) );
AND3x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_356), .C(n_405), .Y(n_119) );
NOR3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_263), .C(n_301), .Y(n_120) );
OAI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_184), .B1(n_238), .B2(n_244), .C1(n_258), .C2(n_261), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_155), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_123), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_123), .B(n_306), .Y(n_397) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g274 ( .A(n_124), .B(n_175), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_124), .B(n_156), .Y(n_282) );
AND2x2_ASAP7_75t_L g317 ( .A(n_124), .B(n_294), .Y(n_317) );
OR2x2_ASAP7_75t_L g341 ( .A(n_124), .B(n_156), .Y(n_341) );
OR2x2_ASAP7_75t_L g349 ( .A(n_124), .B(n_248), .Y(n_349) );
AND2x2_ASAP7_75t_L g352 ( .A(n_124), .B(n_175), .Y(n_352) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g246 ( .A(n_125), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g260 ( .A(n_125), .B(n_175), .Y(n_260) );
AND2x2_ASAP7_75t_L g310 ( .A(n_125), .B(n_248), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_125), .B(n_156), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_125), .B(n_409), .Y(n_430) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_132), .B(n_153), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_126), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g198 ( .A(n_126), .Y(n_198) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_126), .A2(n_249), .B(n_256), .Y(n_248) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_127), .Y(n_159) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_128), .B(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
OAI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_136), .B1(n_149), .B2(n_150), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_163), .B(n_164), .C(n_165), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_133), .A2(n_164), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_133), .A2(n_164), .B(n_231), .C(n_232), .Y(n_230) );
INVx4_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_134), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g161 ( .A(n_134), .B(n_151), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_134), .A2(n_443), .B(n_446), .Y(n_442) );
BUFx3_ASAP7_75t_L g462 ( .A(n_134), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_134), .A2(n_469), .B(n_473), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_134), .A2(n_490), .B(n_493), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_134), .A2(n_506), .B(n_510), .Y(n_505) );
INVx2_ASAP7_75t_L g255 ( .A(n_137), .Y(n_255) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
INVx1_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_140) );
INVx2_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx4_ASAP7_75t_L g233 ( .A(n_141), .Y(n_233) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
AND2x2_ASAP7_75t_L g151 ( .A(n_142), .B(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx3_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
INVx1_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
INVx5_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
BUFx3_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
INVx1_ASAP7_75t_L g502 ( .A(n_147), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_150), .A2(n_203), .B(n_204), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_150), .A2(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g449 ( .A(n_152), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_155), .A2(n_349), .B(n_350), .C(n_353), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_155), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_155), .B(n_293), .Y(n_415) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_175), .Y(n_155) );
AND2x2_ASAP7_75t_SL g259 ( .A(n_156), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g273 ( .A(n_156), .Y(n_273) );
AND2x2_ASAP7_75t_L g300 ( .A(n_156), .B(n_294), .Y(n_300) );
INVx1_ASAP7_75t_SL g308 ( .A(n_156), .Y(n_308) );
AND2x2_ASAP7_75t_L g331 ( .A(n_156), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g409 ( .A(n_156), .Y(n_409) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_160), .B(n_173), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g199 ( .A(n_158), .B(n_200), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_158), .B(n_462), .C(n_481), .Y(n_480) );
AO21x1_ASAP7_75t_L g525 ( .A1(n_158), .A2(n_481), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_159), .A2(n_176), .B(n_183), .Y(n_175) );
OA21x2_ASAP7_75t_L g441 ( .A1(n_159), .A2(n_442), .B(n_451), .Y(n_441) );
BUFx2_ASAP7_75t_L g229 ( .A(n_161), .Y(n_229) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_166), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_166), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_167), .A2(n_450), .B1(n_482), .B2(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_167), .A2(n_450), .B1(n_501), .B2(n_503), .Y(n_500) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_167), .A2(n_170), .B1(n_521), .B2(n_522), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_170), .B(n_182), .Y(n_181) );
INVx5_ASAP7_75t_L g193 ( .A(n_170), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_SL g490 ( .A1(n_171), .A2(n_193), .B(n_491), .C(n_492), .Y(n_490) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_172), .Y(n_222) );
INVx1_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
INVx2_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_174), .A2(n_228), .B(n_237), .Y(n_227) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_174), .A2(n_489), .B(n_496), .Y(n_488) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_505), .B(n_513), .Y(n_504) );
BUFx2_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
INVx1_ASAP7_75t_L g307 ( .A(n_175), .Y(n_307) );
INVx3_ASAP7_75t_L g332 ( .A(n_175), .Y(n_332) );
INVx1_ASAP7_75t_L g509 ( .A(n_180), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_184), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_212), .Y(n_184) );
INVx1_ASAP7_75t_L g328 ( .A(n_185), .Y(n_328) );
OAI32xp33_ASAP7_75t_L g334 ( .A1(n_185), .A2(n_273), .A3(n_335), .B1(n_336), .B2(n_337), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_185), .A2(n_339), .B1(n_342), .B2(n_347), .Y(n_338) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g276 ( .A(n_186), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g354 ( .A(n_186), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g424 ( .A(n_186), .B(n_370), .Y(n_424) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_201), .Y(n_186) );
AND2x2_ASAP7_75t_L g239 ( .A(n_187), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
INVx1_ASAP7_75t_L g288 ( .A(n_187), .Y(n_288) );
OR2x2_ASAP7_75t_L g296 ( .A(n_187), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g303 ( .A(n_187), .B(n_277), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_187), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_187), .B(n_242), .Y(n_324) );
INVx3_ASAP7_75t_L g346 ( .A(n_187), .Y(n_346) );
AND2x2_ASAP7_75t_L g371 ( .A(n_187), .B(n_243), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_187), .B(n_336), .Y(n_419) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
AOI21xp5_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_190), .B(n_198), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_195), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_193), .A2(n_253), .B(n_254), .C(n_255), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_193), .A2(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g450 ( .A(n_193), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_193), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_195), .A2(n_206), .B(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g236 ( .A(n_197), .Y(n_236) );
INVx1_ASAP7_75t_L g208 ( .A(n_198), .Y(n_208) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_198), .A2(n_454), .B(n_463), .Y(n_453) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_198), .A2(n_468), .B(n_476), .Y(n_467) );
INVx2_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
AND2x2_ASAP7_75t_L g375 ( .A(n_201), .B(n_213), .Y(n_375) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_208), .B(n_209), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_211), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_211), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g417 ( .A(n_212), .Y(n_417) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx1_ASAP7_75t_L g262 ( .A(n_213), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_213), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_213), .B(n_243), .Y(n_297) );
AND2x2_ASAP7_75t_L g355 ( .A(n_213), .B(n_278), .Y(n_355) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g241 ( .A(n_214), .Y(n_241) );
AND2x2_ASAP7_75t_L g268 ( .A(n_214), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g277 ( .A(n_214), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_214), .B(n_243), .Y(n_343) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_222), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_226), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_226), .B(n_243), .Y(n_336) );
AND2x2_ASAP7_75t_L g345 ( .A(n_226), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g370 ( .A(n_226), .Y(n_370) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g242 ( .A(n_227), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g278 ( .A(n_227), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_233), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g472 ( .A(n_233), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_233), .A2(n_494), .B(n_495), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_238), .A2(n_248), .B1(n_407), .B2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_240), .A2(n_351), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_241), .B(n_346), .Y(n_363) );
INVx1_ASAP7_75t_L g388 ( .A(n_241), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_242), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g315 ( .A(n_242), .B(n_268), .Y(n_315) );
INVx2_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
INVx1_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_244), .A2(n_396), .B1(n_413), .B2(n_416), .C(n_418), .Y(n_412) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g283 ( .A(n_245), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_245), .B(n_294), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_246), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g337 ( .A(n_246), .B(n_283), .Y(n_337) );
INVx3_ASAP7_75t_SL g378 ( .A(n_246), .Y(n_378) );
AND2x2_ASAP7_75t_L g322 ( .A(n_247), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g351 ( .A(n_247), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_247), .B(n_260), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_247), .B(n_306), .Y(n_392) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g294 ( .A(n_248), .Y(n_294) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_248), .A2(n_320), .A3(n_342), .B1(n_390), .B2(n_392), .C1(n_393), .C2(n_394), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_255), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_259), .A2(n_262), .B(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_SL g339 ( .A(n_260), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g361 ( .A(n_260), .B(n_273), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_260), .B(n_300), .Y(n_376) );
INVxp67_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_262), .A2(n_334), .B(n_338), .C(n_348), .Y(n_333) );
OAI221xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_272), .B1(n_275), .B2(n_279), .C(n_284), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g287 ( .A(n_271), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g404 ( .A(n_271), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_272), .A2(n_421), .B1(n_426), .B2(n_427), .C(n_429), .Y(n_420) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_273), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g320 ( .A(n_273), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_273), .B(n_351), .Y(n_358) );
AND2x2_ASAP7_75t_L g400 ( .A(n_273), .B(n_378), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_274), .B(n_299), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_274), .A2(n_286), .B1(n_396), .B2(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g426 ( .A(n_274), .B(n_294), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g403 ( .A(n_277), .Y(n_403) );
AND2x2_ASAP7_75t_L g428 ( .A(n_277), .B(n_371), .Y(n_428) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_SL g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g292 ( .A(n_282), .B(n_293), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_291), .B1(n_295), .B2(n_298), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g359 ( .A(n_287), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_287), .B(n_327), .Y(n_394) );
AOI322xp5_ASAP7_75t_L g318 ( .A1(n_289), .A2(n_319), .A3(n_321), .B1(n_322), .B2(n_324), .C1(n_325), .C2(n_329), .Y(n_318) );
INVxp67_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_292), .A2(n_297), .B1(n_314), .B2(n_316), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_293), .B(n_306), .Y(n_393) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_294), .B(n_332), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_294), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g390 ( .A(n_296), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND3xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_318), .C(n_333), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_309), .B2(n_311), .C(n_313), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_305), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g319 ( .A(n_310), .B(n_320), .Y(n_319) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_312), .Y(n_391) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_317), .B(n_331), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_320), .B(n_378), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_321), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g396 ( .A(n_324), .Y(n_396) );
AND2x2_ASAP7_75t_L g411 ( .A(n_324), .B(n_388), .Y(n_411) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_335), .A2(n_406), .B(n_412), .C(n_420), .Y(n_405) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g374 ( .A(n_345), .B(n_375), .Y(n_374) );
NAND2x1_ASAP7_75t_SL g416 ( .A(n_346), .B(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_349), .Y(n_386) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
AND2x2_ASAP7_75t_L g385 ( .A(n_355), .B(n_371), .Y(n_385) );
NOR5xp2_ASAP7_75t_L g356 ( .A(n_357), .B(n_372), .C(n_389), .D(n_395), .E(n_398), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_360), .B2(n_362), .C(n_364), .Y(n_357) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_361), .B(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_371), .B(n_388), .Y(n_387) );
OAI221xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_376), .B1(n_377), .B2(n_379), .C(n_382), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
AOI211xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_401), .B(n_403), .C(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
CKINVDCx14_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g719 ( .A(n_434), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_435), .B(n_638), .Y(n_434) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_596), .Y(n_435) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_437), .B(n_536), .C(n_572), .D(n_586), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_484), .B1(n_514), .B2(n_523), .C(n_527), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_438), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_464), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_452), .Y(n_440) );
AND2x2_ASAP7_75t_L g533 ( .A(n_441), .B(n_453), .Y(n_533) );
INVx3_ASAP7_75t_L g541 ( .A(n_441), .Y(n_541) );
AND2x2_ASAP7_75t_L g595 ( .A(n_441), .B(n_467), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_441), .B(n_466), .Y(n_631) );
AND2x2_ASAP7_75t_L g689 ( .A(n_441), .B(n_551), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_450), .Y(n_446) );
INVx2_ASAP7_75t_L g460 ( .A(n_449), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_450), .A2(n_460), .B(n_474), .C(n_475), .Y(n_473) );
AND2x2_ASAP7_75t_L g524 ( .A(n_452), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g538 ( .A(n_452), .B(n_467), .Y(n_538) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_453), .B(n_467), .Y(n_553) );
AND2x2_ASAP7_75t_L g565 ( .A(n_453), .B(n_541), .Y(n_565) );
OR2x2_ASAP7_75t_L g567 ( .A(n_453), .B(n_525), .Y(n_567) );
AND2x2_ASAP7_75t_L g602 ( .A(n_453), .B(n_525), .Y(n_602) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_453), .Y(n_647) );
INVx1_ASAP7_75t_L g655 ( .A(n_453), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B(n_462), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_464), .A2(n_573), .B1(n_577), .B2(n_581), .C(n_582), .Y(n_572) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g532 ( .A(n_465), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_477), .Y(n_465) );
INVx2_ASAP7_75t_L g531 ( .A(n_466), .Y(n_531) );
AND2x2_ASAP7_75t_L g584 ( .A(n_466), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g603 ( .A(n_466), .B(n_541), .Y(n_603) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g666 ( .A(n_467), .B(n_541), .Y(n_666) );
AND2x2_ASAP7_75t_L g588 ( .A(n_477), .B(n_533), .Y(n_588) );
OAI322xp33_ASAP7_75t_L g656 ( .A1(n_477), .A2(n_612), .A3(n_657), .B1(n_659), .B2(n_662), .C1(n_664), .C2(n_668), .Y(n_656) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_478), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
AND2x2_ASAP7_75t_L g661 ( .A(n_478), .B(n_541), .Y(n_661) );
AND2x2_ASAP7_75t_L g693 ( .A(n_478), .B(n_565), .Y(n_693) );
OR2x2_ASAP7_75t_L g696 ( .A(n_478), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g526 ( .A(n_479), .Y(n_526) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
INVx1_ASAP7_75t_L g709 ( .A(n_486), .Y(n_709) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g516 ( .A(n_487), .B(n_504), .Y(n_516) );
INVx2_ASAP7_75t_L g549 ( .A(n_487), .Y(n_549) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g571 ( .A(n_488), .Y(n_571) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_488), .Y(n_579) );
OR2x2_ASAP7_75t_L g703 ( .A(n_488), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g528 ( .A(n_497), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g568 ( .A(n_497), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g620 ( .A(n_497), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
AND2x2_ASAP7_75t_L g517 ( .A(n_498), .B(n_518), .Y(n_517) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_498), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g629 ( .A(n_498), .B(n_519), .Y(n_629) );
OR2x2_ASAP7_75t_L g637 ( .A(n_498), .B(n_571), .Y(n_637) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g546 ( .A(n_499), .Y(n_546) );
AND2x2_ASAP7_75t_L g556 ( .A(n_499), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g580 ( .A(n_499), .B(n_504), .Y(n_580) );
AND2x2_ASAP7_75t_L g644 ( .A(n_499), .B(n_519), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_504), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_504), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g557 ( .A(n_504), .Y(n_557) );
INVx1_ASAP7_75t_L g562 ( .A(n_504), .Y(n_562) );
AND2x2_ASAP7_75t_L g574 ( .A(n_504), .B(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_504), .Y(n_652) );
INVx1_ASAP7_75t_L g704 ( .A(n_504), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
AND2x2_ASAP7_75t_L g681 ( .A(n_515), .B(n_590), .Y(n_681) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g608 ( .A(n_517), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g707 ( .A(n_517), .B(n_642), .Y(n_707) );
INVx1_ASAP7_75t_L g529 ( .A(n_518), .Y(n_529) );
AND2x2_ASAP7_75t_L g555 ( .A(n_518), .B(n_549), .Y(n_555) );
BUFx2_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_519), .Y(n_535) );
INVx1_ASAP7_75t_L g545 ( .A(n_519), .Y(n_545) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_523), .B(n_530), .Y(n_683) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI32xp33_ASAP7_75t_L g527 ( .A1(n_524), .A2(n_528), .A3(n_530), .B1(n_532), .B2(n_534), .Y(n_527) );
AND2x2_ASAP7_75t_L g667 ( .A(n_524), .B(n_540), .Y(n_667) );
AND2x2_ASAP7_75t_L g705 ( .A(n_524), .B(n_603), .Y(n_705) );
INVx1_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_529), .B(n_591), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_530), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_530), .B(n_533), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_530), .B(n_602), .Y(n_684) );
OR2x2_ASAP7_75t_L g698 ( .A(n_530), .B(n_567), .Y(n_698) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g625 ( .A(n_531), .B(n_533), .Y(n_625) );
OR2x2_ASAP7_75t_L g634 ( .A(n_531), .B(n_621), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_533), .B(n_584), .Y(n_606) );
INVx2_ASAP7_75t_L g621 ( .A(n_535), .Y(n_621) );
OR2x2_ASAP7_75t_L g636 ( .A(n_535), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_652), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_535), .A2(n_628), .B(n_709), .C(n_710), .Y(n_708) );
OAI321xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_542), .A3(n_547), .B1(n_550), .B2(n_554), .C(n_558), .Y(n_536) );
INVx1_ASAP7_75t_L g649 ( .A(n_537), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g660 ( .A(n_538), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g612 ( .A(n_540), .Y(n_612) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_541), .B(n_655), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_542), .A2(n_680), .B1(n_682), .B2(n_684), .C(n_685), .Y(n_679) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g617 ( .A(n_544), .B(n_591), .Y(n_617) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_545), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g590 ( .A(n_546), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_547), .A2(n_588), .B(n_633), .C(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g599 ( .A(n_549), .B(n_556), .Y(n_599) );
BUFx2_ASAP7_75t_L g609 ( .A(n_549), .Y(n_609) );
INVx1_ASAP7_75t_L g624 ( .A(n_549), .Y(n_624) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OR2x2_ASAP7_75t_L g630 ( .A(n_552), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g713 ( .A(n_552), .Y(n_713) );
INVx1_ASAP7_75t_L g706 ( .A(n_553), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g559 ( .A(n_555), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g663 ( .A(n_555), .B(n_580), .Y(n_663) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_563), .B1(n_566), .B2(n_568), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_560), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g628 ( .A(n_561), .B(n_629), .Y(n_628) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_562), .B(n_571), .Y(n_591) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g583 ( .A(n_565), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g593 ( .A(n_567), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_570), .A2(n_688), .B1(n_690), .B2(n_691), .C(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g576 ( .A(n_571), .Y(n_576) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_571), .Y(n_642) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_574), .B(n_693), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_575), .A2(n_580), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_578), .B(n_588), .Y(n_685) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g654 ( .A(n_579), .Y(n_654) );
AND2x2_ASAP7_75t_L g613 ( .A(n_580), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g702 ( .A(n_580), .Y(n_702) );
INVx1_ASAP7_75t_L g618 ( .A(n_583), .Y(n_618) );
INVx1_ASAP7_75t_L g673 ( .A(n_584), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B1(n_592), .B2(n_593), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_590), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_591), .B(n_629), .Y(n_695) );
OR2x2_ASAP7_75t_L g668 ( .A(n_592), .B(n_621), .Y(n_668) );
INVx1_ASAP7_75t_L g607 ( .A(n_593), .Y(n_607) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_595), .B(n_646), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_615), .C(n_626), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_604), .C(n_610), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_599), .A2(n_670), .B1(n_674), .B2(n_677), .C(n_679), .Y(n_669) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g611 ( .A(n_602), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g665 ( .A(n_602), .B(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_603), .A2(n_651), .B(n_653), .C(n_655), .Y(n_650) );
INVx2_ASAP7_75t_L g697 ( .A(n_603), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_608), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g676 ( .A(n_609), .B(n_629), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_618), .B(n_619), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_622), .B(n_625), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_620), .B(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_625), .B(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B(n_632), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g653 ( .A(n_629), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND4x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_669), .C(n_686), .D(n_708), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_656), .Y(n_639) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_645), .B(n_648), .C(n_650), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_644), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_655), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g690 ( .A(n_665), .Y(n_690) );
INVx2_ASAP7_75t_SL g678 ( .A(n_666), .Y(n_678) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g691 ( .A(n_676), .Y(n_691) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_694), .Y(n_686) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
OAI221xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g720 ( .A(n_715), .Y(n_720) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
BUFx4f_ASAP7_75t_SL g738 ( .A(n_731), .Y(n_738) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
endmodule