module real_jpeg_11265_n_13 (n_5, n_4, n_8, n_0, n_12, n_57, n_1, n_11, n_2, n_56, n_6, n_7, n_55, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_57;
input n_1;
input n_11;
input n_2;
input n_56;
input n_6;
input n_7;
input n_55;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_49;
wire n_52;
wire n_31;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_27;
wire n_30;
wire n_16;
wire n_15;

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_55),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_3),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_56),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_12),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI221xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_20),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_18),
.B2(n_50),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g50 ( 
.A1(n_20),
.A2(n_37),
.A3(n_46),
.B1(n_48),
.B2(n_51),
.C1(n_52),
.C2(n_53),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_32),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_24),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_32),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_35),
.B(n_36),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);


endmodule