module fake_ariane_1433_n_1211 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1211);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1211;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_1167;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_670;
wire n_607;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_1131;
wire n_1187;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_790;
wire n_207;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_779;
wire n_336;
wire n_754;
wire n_731;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1201;
wire n_1107;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_218;
wire n_1099;
wire n_271;
wire n_1153;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_1207;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_1074;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_206;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_1121;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_1194;
wire n_907;
wire n_225;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_888;
wire n_845;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_571;
wire n_414;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_609;
wire n_212;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_171;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_215;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_213;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_999;
wire n_967;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_204;
wire n_615;
wire n_1070;
wire n_1027;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_1102;
wire n_360;
wire n_1101;
wire n_975;
wire n_1129;
wire n_1189;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_1011;
wire n_211;
wire n_642;
wire n_978;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_54),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_56),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_45),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_33),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_20),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_39),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_136),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_79),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_32),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_84),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_24),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_167),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_66),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_48),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_26),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_65),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_52),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_80),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_103),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_185),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_190),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_183),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_195),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_203),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_221),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_171),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_233),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_258),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_230),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_230),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_232),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_231),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_231),
.B(n_208),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_245),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_243),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_238),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_229),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_229),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_293),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_266),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_272),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_260),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_304),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_267),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_307),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_292),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_298),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_288),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_290),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_281),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_273),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_294),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_312),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_329),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_331),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_315),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_262),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_308),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_308),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_262),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_310),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_336),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_318),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_342),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_320),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_321),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_302),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_313),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_348),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_321),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_323),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_332),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_332),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_273),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_353),
.B1(n_324),
.B2(n_323),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

AOI22x1_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_334),
.B1(n_176),
.B2(n_177),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_337),
.B(n_309),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_376),
.A2(n_325),
.B1(n_324),
.B2(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_335),
.B1(n_349),
.B2(n_319),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_335),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_345),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_299),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_338),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_341),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_363),
.Y(n_424)
);

BUFx8_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_372),
.B(n_341),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_366),
.A2(n_325),
.B1(n_299),
.B2(n_298),
.Y(n_428)
);

CKINVDCx8_ASAP7_75t_R g429 ( 
.A(n_375),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_291),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_392),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g433 ( 
.A(n_357),
.B(n_296),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_296),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_398),
.A2(n_287),
.B1(n_279),
.B2(n_346),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_343),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_387),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_389),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_395),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_265),
.Y(n_453)
);

OAI22x1_ASAP7_75t_SL g454 ( 
.A1(n_381),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_374),
.A2(n_173),
.B1(n_179),
.B2(n_186),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_369),
.B(n_265),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_354),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_179),
.Y(n_462)
);

BUFx12f_ASAP7_75t_L g463 ( 
.A(n_359),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_368),
.B(n_191),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_359),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_359),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_368),
.B(n_175),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_354),
.B(n_223),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_368),
.B(n_180),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g471 ( 
.A(n_359),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_368),
.B(n_181),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_410),
.B(n_401),
.C(n_431),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_399),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_424),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_434),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_424),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_434),
.B(n_202),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_465),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_465),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_441),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_276),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_411),
.B(n_432),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_463),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_463),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_416),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_277),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_425),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_186),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_283),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_411),
.B(n_196),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_196),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_425),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_473),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_425),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_437),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_429),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_400),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_429),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_421),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_458),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_421),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_426),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_426),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_467),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_500),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_524),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_441),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_513),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_520),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_528),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_506),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_520),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_477),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_528),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_477),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_480),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_489),
.B(n_420),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_480),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_497),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_482),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_505),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_516),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_516),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_482),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_484),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_484),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_490),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_R g558 ( 
.A(n_526),
.B(n_490),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_509),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_524),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_491),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_491),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_492),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_492),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_521),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_537),
.Y(n_569)
);

INVxp33_ASAP7_75t_L g570 ( 
.A(n_561),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_475),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_545),
.B(n_489),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_531),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_533),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_550),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_537),
.B(n_481),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_550),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_536),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_534),
.A2(n_428),
.B1(n_501),
.B2(n_455),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_568),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_550),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_558),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_536),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_532),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_562),
.B(n_479),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_SL g593 ( 
.A(n_541),
.B(n_501),
.C(n_430),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_539),
.A2(n_481),
.B1(n_474),
.B2(n_489),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_543),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_483),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_560),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_535),
.B(n_452),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_560),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_544),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_540),
.B(n_450),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_567),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_546),
.B(n_448),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_549),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_551),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

OAI21xp33_ASAP7_75t_SL g615 ( 
.A1(n_552),
.A2(n_450),
.B(n_446),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_553),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_538),
.A2(n_427),
.B1(n_438),
.B2(n_515),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_SL g619 ( 
.A1(n_538),
.A2(n_494),
.B(n_493),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_548),
.B(n_522),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_557),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_563),
.B(n_441),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_555),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_556),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_417),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_565),
.B(n_452),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_559),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_541),
.Y(n_631)
);

INVx4_ASAP7_75t_SL g632 ( 
.A(n_545),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_545),
.A2(n_436),
.B1(n_411),
.B2(n_432),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_541),
.B(n_443),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_537),
.B(n_456),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_541),
.B(n_443),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_537),
.B(n_495),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_537),
.B(n_510),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_537),
.B(n_452),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_537),
.B(n_441),
.Y(n_642)
);

NAND2x1p5_ASAP7_75t_L g643 ( 
.A(n_545),
.B(n_476),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_537),
.B(n_442),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_537),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_531),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_541),
.B(n_444),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_531),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_545),
.A2(n_432),
.B1(n_445),
.B2(n_412),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_531),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_569),
.B(n_512),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_593),
.B(n_444),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_623),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_588),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_596),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_610),
.B(n_466),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_637),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_645),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_638),
.B(n_517),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_617),
.A2(n_470),
.B1(n_472),
.B2(n_468),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_590),
.B(n_459),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_573),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_583),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_634),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_631),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_580),
.A2(n_499),
.B1(n_487),
.B2(n_504),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_632),
.B(n_507),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_623),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_598),
.B(n_518),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_619),
.B(n_197),
.C(n_189),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_613),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_592),
.B(n_521),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_616),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_579),
.B(n_525),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_577),
.B(n_507),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_629),
.B(n_525),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_623),
.B(n_466),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_587),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_636),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_579),
.B(n_527),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_632),
.B(n_527),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_571),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_582),
.B(n_423),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_623),
.A2(n_469),
.B1(n_470),
.B2(n_468),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_592),
.B(n_414),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_632),
.B(n_478),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_571),
.Y(n_695)
);

CKINVDCx6p67_ASAP7_75t_R g696 ( 
.A(n_631),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_588),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_630),
.B(n_423),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_623),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_629),
.B(n_503),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_630),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_601),
.B(n_423),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_614),
.B(n_523),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_633),
.A2(n_445),
.B1(n_454),
.B2(n_468),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_609),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_623),
.Y(n_706)
);

BUFx4f_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_650),
.A2(n_472),
.B1(n_470),
.B2(n_453),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_609),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_648),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_589),
.B(n_488),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_589),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_649),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_589),
.B(n_488),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_651),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_614),
.B(n_420),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_589),
.B(n_488),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_600),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_647),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_600),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_600),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_611),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_611),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_596),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_635),
.B(n_519),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_614),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_587),
.B(n_223),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_631),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_612),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_575),
.B(n_488),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_570),
.B(n_462),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_612),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_570),
.B(n_496),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_622),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_659),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_705),
.Y(n_740)
);

AND2x2_ASAP7_75t_SL g741 ( 
.A(n_683),
.B(n_605),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_710),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_669),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_683),
.B(n_601),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_721),
.B(n_604),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_665),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_724),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_668),
.B(n_627),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_660),
.B(n_639),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_699),
.B(n_627),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_668),
.B(n_622),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_653),
.B(n_639),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_707),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_658),
.B(n_604),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_699),
.B(n_620),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_662),
.B(n_642),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_661),
.B(n_578),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_664),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_666),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_661),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_699),
.B(n_577),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_676),
.B(n_605),
.C(n_642),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_667),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_670),
.A2(n_663),
.B1(n_709),
.B2(n_676),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_657),
.B(n_730),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_625),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_700),
.B(n_644),
.C(n_615),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_653),
.B(n_618),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_687),
.B(n_625),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_699),
.B(n_626),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_SL g772 ( 
.A(n_655),
.B(n_626),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_663),
.A2(n_595),
.B1(n_572),
.B2(n_472),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_704),
.A2(n_572),
.B1(n_486),
.B2(n_628),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_675),
.B(n_618),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_709),
.A2(n_451),
.B1(n_442),
.B2(n_643),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_720),
.B(n_621),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_673),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_677),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_687),
.B(n_624),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_690),
.B(n_695),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_684),
.B(n_578),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_675),
.B(n_602),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_679),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_689),
.B(n_643),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_697),
.B(n_0),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_685),
.B(n_602),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_707),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_711),
.B(n_606),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_654),
.B(n_698),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_689),
.B(n_641),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_725),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_735),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_691),
.B(n_656),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_714),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_655),
.B(n_606),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_716),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_727),
.B(n_0),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_726),
.B(n_641),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_693),
.B(n_606),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_726),
.B(n_641),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_719),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_738),
.B(n_1),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_703),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_703),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_702),
.B(n_575),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_669),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_717),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_702),
.B(n_575),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_760),
.B(n_701),
.Y(n_812)
);

AO22x2_ASAP7_75t_L g813 ( 
.A1(n_740),
.A2(n_574),
.B1(n_581),
.B2(n_576),
.Y(n_813)
);

NOR2x1p5_ASAP7_75t_L g814 ( 
.A(n_760),
.B(n_696),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_793),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_805),
.B(n_729),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_746),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_759),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_764),
.A2(n_572),
.B1(n_734),
.B2(n_700),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_794),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_763),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_742),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_757),
.B(n_694),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_806),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_747),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_741),
.B(n_791),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_771),
.Y(n_827)
);

OR2x6_ASAP7_75t_SL g828 ( 
.A(n_764),
.B(n_669),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_810),
.B(n_729),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_778),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_745),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_779),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_784),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_796),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_798),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_757),
.B(n_674),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_758),
.B(n_686),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_788),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_754),
.B(n_731),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_768),
.B(n_717),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_803),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_766),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_739),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_768),
.B(n_686),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_808),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_775),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_801),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_762),
.A2(n_692),
.B1(n_572),
.B2(n_681),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_782),
.B(n_674),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_775),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_781),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_783),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_752),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_761),
.B(n_706),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_752),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_750),
.B(n_720),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_782),
.B(n_706),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_783),
.B(n_737),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_773),
.A2(n_692),
.B1(n_572),
.B2(n_464),
.Y(n_859)
);

INVx4_ASAP7_75t_SL g860 ( 
.A(n_797),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_787),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_787),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_790),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_772),
.B(n_672),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_790),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_756),
.A2(n_574),
.B1(n_581),
.B2(n_576),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_795),
.Y(n_867)
);

OR2x2_ASAP7_75t_SL g868 ( 
.A(n_767),
.B(n_749),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_743),
.Y(n_869)
);

AO22x2_ASAP7_75t_L g870 ( 
.A1(n_776),
.A2(n_599),
.B1(n_603),
.B2(n_594),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_776),
.A2(n_572),
.B1(n_681),
.B2(n_682),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_797),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_797),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_774),
.A2(n_464),
.B1(n_418),
.B2(n_422),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_809),
.B(n_736),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_807),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_753),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_780),
.B(n_682),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_744),
.B(n_672),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_811),
.B(n_736),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_748),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_751),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_753),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_755),
.B(n_720),
.Y(n_884)
);

AO22x2_ASAP7_75t_L g885 ( 
.A1(n_769),
.A2(n_599),
.B1(n_603),
.B2(n_594),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_792),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_753),
.B(n_694),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_867),
.B(n_786),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_812),
.B(n_770),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_824),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_853),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_877),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_842),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_853),
.B(n_804),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_855),
.B(n_777),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_868),
.A2(n_799),
.B1(n_785),
.B2(n_688),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_855),
.B(n_733),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_708),
.Y(n_898)
);

NOR2x2_ASAP7_75t_L g899 ( 
.A(n_828),
.B(n_765),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_837),
.B(n_708),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_876),
.B(n_680),
.C(n_712),
.Y(n_901)
);

AO22x1_ASAP7_75t_L g902 ( 
.A1(n_887),
.A2(n_789),
.B1(n_722),
.B2(n_723),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_823),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_824),
.Y(n_904)
);

INVx5_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_831),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_854),
.B(n_713),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_852),
.B(n_713),
.Y(n_908)
);

BUFx12f_ASAP7_75t_SL g909 ( 
.A(n_836),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_826),
.A2(n_223),
.B(n_800),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_813),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_813),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_861),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_862),
.B(n_722),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_860),
.B(n_723),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_863),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_865),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_839),
.B(n_789),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_819),
.A2(n_208),
.B(n_200),
.C(n_201),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_881),
.A2(n_206),
.B(n_207),
.C(n_198),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_869),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_878),
.B(n_882),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_840),
.B(n_585),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_816),
.B(n_585),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_829),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_829),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_860),
.B(n_836),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_846),
.B(n_585),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_817),
.Y(n_929)
);

AND2x4_ASAP7_75t_SL g930 ( 
.A(n_849),
.B(n_789),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_813),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_818),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_SL g933 ( 
.A(n_814),
.B(n_802),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_847),
.B(n_586),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_821),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_850),
.B(n_586),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_887),
.A2(n_586),
.B1(n_640),
.B2(n_469),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_840),
.B(n_640),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_896),
.A2(n_854),
.B(n_880),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_925),
.B(n_844),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_927),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_913),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_937),
.B(n_864),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_926),
.B(n_843),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_896),
.A2(n_880),
.B(n_856),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_894),
.B(n_895),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_906),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_920),
.A2(n_884),
.B(n_885),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_922),
.A2(n_871),
.B1(n_879),
.B2(n_848),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_902),
.A2(n_907),
.B(n_895),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_894),
.B(n_886),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_903),
.B(n_875),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_888),
.B(n_827),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_916),
.B(n_830),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_919),
.A2(n_833),
.B(n_834),
.C(n_832),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_910),
.A2(n_885),
.B1(n_851),
.B2(n_870),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_905),
.B(n_860),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_917),
.B(n_835),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_921),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_891),
.B(n_841),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_890),
.A2(n_885),
.B(n_883),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_924),
.A2(n_872),
.B(n_873),
.C(n_858),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_933),
.A2(n_884),
.B(n_879),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_938),
.B(n_866),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_927),
.A2(n_870),
.B(n_857),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_900),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_905),
.A2(n_857),
.B(n_849),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_905),
.A2(n_866),
.B(n_864),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_905),
.A2(n_866),
.B(n_718),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_910),
.A2(n_715),
.B(n_874),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_938),
.B(n_815),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_929),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_892),
.B(n_820),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_899),
.A2(n_859),
.B(n_845),
.C(n_214),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_924),
.A2(n_914),
.B(n_908),
.Y(n_975)
);

CKINVDCx10_ASAP7_75t_R g976 ( 
.A(n_918),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_904),
.A2(n_822),
.B(n_838),
.C(n_825),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_914),
.A2(n_859),
.B(n_640),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_928),
.B(n_936),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_932),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_908),
.A2(n_823),
.B(n_887),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_928),
.A2(n_823),
.B(n_502),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_936),
.B(n_823),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_496),
.B1(n_508),
.B2(n_498),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_909),
.B(n_607),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_889),
.B(n_607),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_901),
.A2(n_897),
.B(n_923),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_911),
.A2(n_215),
.B(n_224),
.C(n_212),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_892),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_935),
.A2(n_226),
.B(n_225),
.Y(n_990)
);

AND2x2_ASAP7_75t_SL g991 ( 
.A(n_930),
.B(n_204),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_898),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_934),
.B(n_227),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_915),
.A2(n_228),
.B(n_219),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_915),
.A2(n_219),
.B(n_204),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_892),
.B(n_496),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_912),
.B(n_1),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_931),
.A2(n_469),
.B(n_213),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_922),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_896),
.A2(n_469),
.B(n_213),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_896),
.A2(n_210),
.B(n_220),
.C(n_218),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_911),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_939),
.B(n_496),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_946),
.B(n_2),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_950),
.B(n_496),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_999),
.B(n_498),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_963),
.B(n_498),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_985),
.B(n_498),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_985),
.B(n_498),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_941),
.B(n_442),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_981),
.B(n_508),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_945),
.B(n_508),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_941),
.B(n_508),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_987),
.B(n_508),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_952),
.B(n_442),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_SL g1016 ( 
.A(n_966),
.B(n_989),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_967),
.B(n_511),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_965),
.B(n_511),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_975),
.B(n_511),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_968),
.B(n_951),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1000),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1003),
.A2(n_974),
.B1(n_959),
.B2(n_956),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_1016),
.B(n_962),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_1004),
.B(n_1000),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_1014),
.B(n_979),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_1005),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1006),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1012),
.B(n_948),
.C(n_990),
.Y(n_1028)
);

INVx3_ASAP7_75t_SL g1029 ( 
.A(n_1007),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1019),
.A2(n_949),
.B1(n_983),
.B2(n_953),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_1011),
.A2(n_961),
.B(n_964),
.C(n_960),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1017),
.A2(n_992),
.B1(n_943),
.B2(n_982),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1018),
.A2(n_997),
.B(n_957),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1013),
.B(n_942),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_1008),
.A2(n_993),
.B(n_994),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1015),
.B(n_972),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_1009),
.B(n_991),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1010),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_1016),
.B(n_978),
.C(n_984),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_1020),
.A2(n_977),
.B(n_988),
.C(n_970),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_1016),
.B(n_980),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1016),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1004),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1004),
.B(n_944),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1020),
.A2(n_995),
.B(n_955),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1021),
.A2(n_998),
.B(n_969),
.Y(n_1046)
);

BUFx4_ASAP7_75t_SL g1047 ( 
.A(n_1042),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_1024),
.B(n_947),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1043),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_1023),
.A2(n_973),
.B(n_943),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1044),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_1038),
.B(n_1026),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_1048),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_1050),
.B(n_1035),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1051),
.B(n_1024),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_1053),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1054),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1057),
.A2(n_1048),
.B1(n_1047),
.B2(n_1029),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_1052),
.B(n_1046),
.Y(n_1060)
);

INVx3_ASAP7_75t_SL g1061 ( 
.A(n_1059),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_1060),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1062),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1061),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_1064),
.A2(n_1056),
.B(n_1058),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1066),
.B(n_1057),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1065),
.B(n_1056),
.Y(n_1068)
);

NAND2xp33_ASAP7_75t_SL g1069 ( 
.A(n_1067),
.B(n_1039),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_1068),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1070),
.B(n_1049),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_1070),
.A2(n_1045),
.B(n_1040),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1071),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1072),
.B(n_1073),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1073),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_1026),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1075),
.B(n_1026),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_1076),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1080),
.Y(n_1081)
);

CKINVDCx8_ASAP7_75t_R g1082 ( 
.A(n_1079),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_1022),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_199),
.C(n_1031),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1083),
.B(n_1041),
.Y(n_1085)
);

AOI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_1030),
.B1(n_1032),
.B2(n_1027),
.C1(n_1036),
.C2(n_1034),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1027),
.B1(n_1025),
.B2(n_1033),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1037),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1088),
.B(n_2),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1087),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1088),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1091),
.B(n_3),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1090),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_SL g1094 ( 
.A(n_1089),
.B(n_976),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1093),
.B(n_1002),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1095),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_1092),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1097),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_R g1100 ( 
.A(n_1098),
.B(n_210),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_3),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_218),
.B1(n_220),
.B2(n_194),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1102),
.B(n_4),
.Y(n_1103)
);

OAI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_192),
.B1(n_193),
.B2(n_419),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_209),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1106),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_4),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1106),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_1107),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1109),
.A2(n_209),
.B(n_270),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1108),
.B(n_5),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1110),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_7),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1113),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1114),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1115),
.B(n_1111),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_1116),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1118),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_271),
.B(n_270),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1119),
.B(n_271),
.C(n_209),
.Y(n_1121)
);

OAI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_209),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_996),
.B1(n_418),
.B2(n_943),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_418),
.B1(n_9),
.B2(n_10),
.Y(n_1124)
);

XNOR2x1_ASAP7_75t_L g1125 ( 
.A(n_1124),
.B(n_8),
.Y(n_1125)
);

OAI21xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1123),
.A2(n_8),
.B(n_11),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1124),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1125),
.A2(n_433),
.B1(n_958),
.B2(n_954),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1126),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1127),
.B(n_12),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1129),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_998),
.B1(n_295),
.B2(n_285),
.C(n_283),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1131),
.A2(n_1128),
.B1(n_971),
.B2(n_940),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1134),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_453),
.B1(n_422),
.B2(n_461),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_13),
.C(n_14),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_SL g1138 ( 
.A(n_1136),
.B(n_15),
.C(n_16),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1138),
.B(n_16),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1137),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1139),
.A2(n_1140),
.B1(n_18),
.B2(n_19),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1142),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1142),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1143),
.B(n_17),
.C(n_20),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_1147)
);

NAND4xp25_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_21),
.C(n_23),
.D(n_25),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1146),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1150),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_SL g1152 ( 
.A(n_1149),
.B(n_1148),
.C(n_27),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1152),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_28),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1154),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1156)
);

INVxp67_ASAP7_75t_SL g1157 ( 
.A(n_1156),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1157),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1159)
);

AOI31xp33_ASAP7_75t_L g1160 ( 
.A1(n_1158),
.A2(n_34),
.A3(n_35),
.B(n_36),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1159),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_35),
.B(n_36),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1159),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1159),
.B(n_37),
.C(n_38),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1161),
.A2(n_1163),
.B1(n_1164),
.B2(n_1162),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1161),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1161),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1161),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1166),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1167),
.Y(n_1170)
);

XNOR2xp5_ASAP7_75t_L g1171 ( 
.A(n_1168),
.B(n_37),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_1165),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1170),
.A2(n_38),
.B(n_39),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1171),
.A2(n_41),
.B(n_42),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1169),
.A2(n_41),
.B(n_43),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1169),
.B(n_44),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1169),
.A2(n_46),
.B(n_47),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1169),
.A2(n_49),
.B(n_50),
.Y(n_1178)
);

OAI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_1169),
.A2(n_51),
.B(n_53),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1169),
.B(n_55),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1169),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1169),
.A2(n_57),
.B(n_58),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1169),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1183)
);

XNOR2xp5_ASAP7_75t_L g1184 ( 
.A(n_1172),
.B(n_63),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1181),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1178),
.Y(n_1186)
);

AOI222xp33_ASAP7_75t_L g1187 ( 
.A1(n_1179),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.C1(n_77),
.C2(n_81),
.Y(n_1187)
);

AOI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_1174),
.A2(n_82),
.B(n_83),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1183),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1176),
.A2(n_1180),
.B1(n_1175),
.B2(n_1177),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1182),
.B(n_89),
.Y(n_1191)
);

AOI222xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1173),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.C1(n_93),
.C2(n_94),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1190),
.A2(n_986),
.B(n_97),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1187),
.B(n_96),
.Y(n_1194)
);

OAI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1188),
.A2(n_1184),
.B1(n_1185),
.B2(n_1186),
.C1(n_1192),
.C2(n_1191),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1189),
.A2(n_98),
.B(n_99),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1190),
.B(n_100),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_SL g1198 ( 
.A1(n_1190),
.A2(n_101),
.B(n_104),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1190),
.B(n_105),
.C(n_106),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1195),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1197),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1199),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1198),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_1203)
);

AOI322xp5_ASAP7_75t_L g1204 ( 
.A1(n_1202),
.A2(n_1194),
.A3(n_1193),
.B1(n_1196),
.B2(n_125),
.C1(n_126),
.C2(n_127),
.Y(n_1204)
);

OAI332xp33_ASAP7_75t_L g1205 ( 
.A1(n_1200),
.A2(n_121),
.A3(n_122),
.B1(n_124),
.B2(n_130),
.B3(n_131),
.C1(n_135),
.C2(n_137),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1204),
.A2(n_1201),
.B(n_1203),
.Y(n_1206)
);

OAI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1206),
.A2(n_1205),
.B1(n_139),
.B2(n_141),
.C(n_144),
.Y(n_1207)
);

NOR3xp33_ASAP7_75t_L g1208 ( 
.A(n_1207),
.B(n_138),
.C(n_145),
.Y(n_1208)
);

AOI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.C1(n_154),
.C2(n_155),
.Y(n_1209)
);

AOI211xp5_ASAP7_75t_L g1210 ( 
.A1(n_1209),
.A2(n_156),
.B(n_158),
.C(n_160),
.Y(n_1210)
);

AOI211xp5_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_161),
.B(n_162),
.C(n_164),
.Y(n_1211)
);


endmodule