module real_jpeg_6391_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_89),
.B1(n_189),
.B2(n_193),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_1),
.A2(n_89),
.B1(n_175),
.B2(n_327),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_1),
.A2(n_89),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_3),
.A2(n_59),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_78),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_78),
.B1(n_136),
.B2(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_4),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_152),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_90),
.B1(n_152),
.B2(n_211),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_4),
.A2(n_37),
.B1(n_152),
.B2(n_251),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_91),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_5),
.A2(n_199),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_5),
.A2(n_65),
.B1(n_199),
.B2(n_305),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_5),
.A2(n_199),
.B1(n_222),
.B2(n_405),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_53),
.B1(n_142),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_244),
.C(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_6),
.B(n_138),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_29),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_6),
.B(n_83),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_6),
.B(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_7),
.A2(n_66),
.B1(n_108),
.B2(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_7),
.A2(n_30),
.B1(n_74),
.B2(n_108),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_7),
.A2(n_108),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_9),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_10),
.Y(n_378)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_53),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_12),
.A2(n_264),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_12),
.A2(n_264),
.B1(n_353),
.B2(n_357),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_12),
.A2(n_117),
.B1(n_264),
.B2(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_13),
.Y(n_375)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_15),
.A2(n_45),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_15),
.A2(n_45),
.B1(n_251),
.B2(n_272),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_16),
.A2(n_36),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_227),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_225),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_203),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_20),
.B(n_203),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_121),
.C(n_167),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_21),
.A2(n_22),
.B1(n_121),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_84),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_23),
.A2(n_24),
.B(n_86),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B1(n_86),
.B2(n_120),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_24),
.A2(n_43),
.B1(n_120),
.B2(n_423),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_25),
.A2(n_35),
.B1(n_170),
.B2(n_178),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_25),
.A2(n_249),
.B(n_254),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_25),
.A2(n_237),
.B(n_254),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_25),
.A2(n_385),
.B1(n_386),
.B2(n_389),
.Y(n_384)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_26),
.B(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_26),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_26),
.A2(n_28),
.B1(n_326),
.B2(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_26),
.A2(n_255),
.B1(n_390),
.B2(n_429),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_39),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_40),
.Y(n_282)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_41),
.Y(n_272)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_43),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_56),
.B1(n_77),
.B2(n_83),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_44),
.A2(n_56),
.B1(n_83),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g328 ( 
.A1(n_47),
.A2(n_314),
.A3(n_329),
.B1(n_333),
.B2(n_336),
.Y(n_328)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_48),
.Y(n_263)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_49),
.Y(n_163)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_50),
.Y(n_414)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_51),
.Y(n_186)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_51),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_51),
.Y(n_338)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_55),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_56),
.A2(n_77),
.B1(n_83),
.B2(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_56),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_56),
.B(n_239),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_59),
.B(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_62),
.Y(n_244)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_68),
.A2(n_261),
.B(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_83),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_83),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_106),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_94),
.B(n_107),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_94),
.Y(n_209)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_103),
.B2(n_105),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_97),
.B(n_311),
.Y(n_379)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_100),
.Y(n_321)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_102),
.Y(n_312)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_104),
.Y(n_356)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_104),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_106),
.A2(n_209),
.B(n_432),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_109),
.Y(n_382)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_112),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_113),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_113),
.A2(n_397),
.B(n_401),
.Y(n_396)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_121),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_159),
.B(n_166),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_160),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_138),
.B1(n_146),
.B2(n_153),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_124),
.A2(n_309),
.B(n_318),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_124),
.B(n_359),
.Y(n_358)
);

AOI22x1_ASAP7_75t_L g435 ( 
.A1(n_124),
.A2(n_138),
.B1(n_359),
.B2(n_436),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_124),
.A2(n_318),
.B(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_125),
.A2(n_147),
.B1(n_188),
.B2(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_125),
.A2(n_195),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_125),
.A2(n_195),
.B1(n_352),
.B2(n_404),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_138),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_136),
.Y(n_357)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_138),
.Y(n_195)
);

AO22x2_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_141),
.Y(n_335)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g222 ( 
.A(n_148),
.Y(n_222)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_149),
.A2(n_373),
.A3(n_376),
.B1(n_379),
.B2(n_380),
.Y(n_372)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_166),
.B(n_204),
.CI(n_205),
.CON(n_203),
.SN(n_203)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_167),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_187),
.C(n_196),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_168),
.B(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_181),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_169),
.B(n_181),
.Y(n_446)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_170),
.Y(n_429)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_178),
.A2(n_277),
.B(n_283),
.Y(n_276)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_182),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_183),
.Y(n_306)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_186),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_187),
.B(n_196),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_188),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_194),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_195),
.B(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_195),
.A2(n_352),
.B(n_358),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B(n_202),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_197),
.A2(n_198),
.B1(n_209),
.B2(n_432),
.Y(n_431)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_202),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g479 ( 
.A(n_203),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_214),
.B2(n_224),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_209),
.B(n_237),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_223),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_236),
.B(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_216),
.A2(n_217),
.B1(n_261),
.B2(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_216),
.A2(n_238),
.B(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_216),
.A2(n_217),
.B1(n_408),
.B2(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_217),
.A2(n_265),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI311xp33_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_417),
.A3(n_455),
.B1(n_473),
.C1(n_474),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_366),
.B(n_416),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_343),
.B(n_365),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_298),
.B(n_342),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_268),
.B(n_297),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_247),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_235),
.A2(n_241),
.B1(n_242),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_SL g309 ( 
.A1(n_237),
.A2(n_310),
.B(n_313),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_237),
.B(n_381),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_SL g397 ( 
.A1(n_237),
.A2(n_380),
.B(n_398),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_258),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_259),
.C(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_256),
.A2(n_283),
.B(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_266),
.B2(n_267),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_286),
.B(n_296),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B(n_285),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_284),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_294),
.Y(n_296)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_300),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_323),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_307),
.B2(n_308),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_307),
.C(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_335),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_344),
.B(n_345),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_364),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_349),
.C(n_364),
.Y(n_367)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_360),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_361),
.C(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_367),
.B(n_368),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_394),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_383),
.B2(n_384),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_383),
.Y(n_450)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_391),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_391),
.B(n_392),
.C(n_394),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_402),
.B2(n_415),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_403),
.C(n_407),
.Y(n_464)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_407),
.Y(n_402)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_440),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_SL g474 ( 
.A1(n_418),
.A2(n_440),
.B(n_475),
.C(n_478),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_437),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_437),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.C(n_424),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_422),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.C(n_435),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_428),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_430),
.A2(n_431),
.B1(n_435),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_435),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_453),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_453),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.C(n_447),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_442),
.A2(n_443),
.B1(n_446),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_450),
.C(n_451),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_448),
.A2(n_449),
.B1(n_451),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_451),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_468),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_457),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

NOR2x1_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_465),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_465),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.C(n_464),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_462),
.A2(n_463),
.B1(n_464),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_464),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_470),
.Y(n_476)
);


endmodule