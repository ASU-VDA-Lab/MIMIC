module real_aes_4448_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_1218, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_1217, n_169, n_242, n_308, n_1219, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_1220, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_1216, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_1218;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_1217;
input n_169;
input n_242;
input n_308;
input n_1219;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_1220;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_1216;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1205;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_792;
wire n_386;
wire n_905;
wire n_673;
wire n_518;
wire n_1192;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_1200;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_364;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1123;
wire n_593;
wire n_1137;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_958;
wire n_677;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_1199;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_1213;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_1182;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_369;
wire n_1070;
wire n_1189;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_1210;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_973;
wire n_455;
wire n_725;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1207;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1196;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_1167;
wire n_1100;
wire n_1174;
wire n_688;
wire n_1193;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_363;
wire n_449;
wire n_607;
wire n_417;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_1198;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_1212;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1202;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_1179;
wire n_1201;
wire n_569;
wire n_997;
wire n_563;
wire n_1203;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1014;
wire n_1028;
wire n_1187;
wire n_366;
wire n_727;
wire n_1083;
wire n_649;
wire n_397;
wire n_749;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_377;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_710;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1209;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_1214;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_1208;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_503;
wire n_459;
wire n_558;
wire n_1015;
wire n_1172;
wire n_863;
wire n_998;
wire n_1175;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_1190;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1159;
wire n_1156;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_1211;
wire n_650;
wire n_743;
wire n_646;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_601;
wire n_500;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_1101;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_0), .A2(n_220), .B1(n_550), .B2(n_731), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_1), .A2(n_313), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g854 ( .A(n_2), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_3), .A2(n_263), .B1(n_742), .B2(n_743), .Y(n_866) );
INVx1_ASAP7_75t_L g500 ( .A(n_4), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_5), .A2(n_245), .B1(n_583), .B2(n_589), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_6), .A2(n_177), .B1(n_412), .B2(n_649), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_7), .A2(n_295), .B1(n_483), .B2(n_540), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_8), .A2(n_284), .B1(n_626), .B2(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_9), .A2(n_139), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_10), .A2(n_199), .B1(n_742), .B2(n_943), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_11), .A2(n_275), .B1(n_495), .B2(n_496), .C(n_499), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_12), .A2(n_76), .B1(n_542), .B2(n_543), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_13), .A2(n_224), .B1(n_577), .B2(n_586), .Y(n_932) );
INVx1_ASAP7_75t_L g857 ( .A(n_14), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_15), .A2(n_287), .B1(n_542), .B2(n_548), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_16), .A2(n_18), .B1(n_548), .B2(n_550), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_17), .A2(n_73), .B1(n_517), .B2(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_19), .B(n_387), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_20), .A2(n_129), .B1(n_576), .B2(n_577), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g892 ( .A1(n_21), .A2(n_412), .B(n_893), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_22), .A2(n_229), .B1(n_742), .B2(n_743), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_23), .A2(n_330), .B1(n_966), .B2(n_970), .Y(n_965) );
INVx1_ASAP7_75t_L g750 ( .A(n_24), .Y(n_750) );
INVx1_ASAP7_75t_L g852 ( .A(n_25), .Y(n_852) );
AOI221x1_ASAP7_75t_L g813 ( .A1(n_26), .A2(n_89), .B1(n_641), .B2(n_690), .C(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_27), .A2(n_342), .B1(n_508), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_28), .A2(n_278), .B1(n_517), .B2(n_518), .Y(n_697) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_29), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_30), .A2(n_36), .B1(n_550), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g650 ( .A(n_31), .Y(n_650) );
INVx1_ASAP7_75t_L g919 ( .A(n_32), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_33), .A2(n_357), .B1(n_557), .B2(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_34), .A2(n_266), .B1(n_517), .B2(n_518), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_35), .A2(n_47), .B1(n_608), .B2(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g924 ( .A(n_37), .Y(n_924) );
AOI21xp33_ASAP7_75t_L g951 ( .A1(n_38), .A2(n_594), .B(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g599 ( .A(n_39), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_40), .A2(n_144), .B1(n_479), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_41), .A2(n_236), .B1(n_692), .B2(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_42), .A2(n_286), .B1(n_411), .B2(n_416), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_43), .A2(n_109), .B1(n_579), .B2(n_580), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_44), .B(n_647), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_45), .A2(n_296), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_46), .A2(n_288), .B1(n_407), .B2(n_610), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_48), .A2(n_215), .B1(n_630), .B2(n_742), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_49), .A2(n_55), .B1(n_661), .B2(n_731), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_50), .A2(n_127), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_51), .A2(n_328), .B1(n_452), .B2(n_460), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_52), .A2(n_234), .B1(n_539), .B2(n_540), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_53), .A2(n_218), .B1(n_548), .B2(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_54), .A2(n_344), .B1(n_706), .B2(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_56), .A2(n_329), .B1(n_595), .B2(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_57), .A2(n_427), .B(n_431), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_58), .B(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_59), .A2(n_137), .B1(n_771), .B2(n_772), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_60), .A2(n_354), .B1(n_476), .B2(n_546), .Y(n_545) );
OA22x2_ASAP7_75t_L g385 ( .A1(n_61), .A2(n_154), .B1(n_386), .B2(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g423 ( .A(n_61), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_62), .A2(n_135), .B1(n_579), .B2(n_580), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_63), .A2(n_178), .B1(n_554), .B2(n_555), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_64), .A2(n_194), .B1(n_993), .B2(n_1006), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_65), .A2(n_309), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_66), .A2(n_108), .B1(n_555), .B2(n_891), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_67), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_68), .A2(n_175), .B1(n_973), .B2(n_976), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_69), .A2(n_143), .B1(n_557), .B2(n_1190), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_70), .A2(n_350), .B1(n_576), .B2(n_742), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_71), .A2(n_209), .B1(n_483), .B2(n_540), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_72), .B(n_554), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_74), .A2(n_302), .B1(n_461), .B2(n_540), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_75), .B(n_169), .Y(n_370) );
INVx1_ASAP7_75t_L g393 ( .A(n_75), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g424 ( .A1(n_75), .A2(n_154), .B(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_77), .A2(n_323), .B1(n_476), .B2(n_546), .Y(n_803) );
AO221x2_ASAP7_75t_L g991 ( .A1(n_78), .A2(n_331), .B1(n_973), .B2(n_980), .C(n_992), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_79), .A2(n_246), .B1(n_461), .B2(n_542), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_80), .A2(n_244), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_81), .A2(n_253), .B1(n_476), .B2(n_546), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_82), .A2(n_208), .B1(n_476), .B2(n_479), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_83), .A2(n_170), .B1(n_495), .B2(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_84), .A2(n_317), .B1(n_976), .B2(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_85), .A2(n_337), .B1(n_966), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_86), .A2(n_211), .B1(n_453), .B2(n_520), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g560 ( .A1(n_87), .A2(n_495), .B(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g969 ( .A(n_88), .B(n_262), .Y(n_969) );
INVx1_ASAP7_75t_L g975 ( .A(n_88), .Y(n_975) );
HB1xp67_ASAP7_75t_L g1213 ( .A(n_88), .Y(n_1213) );
AO22x1_ASAP7_75t_L g992 ( .A1(n_90), .A2(n_174), .B1(n_970), .B2(n_993), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_91), .A2(n_281), .B1(n_476), .B2(n_546), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_92), .A2(n_150), .B1(n_557), .B2(n_610), .Y(n_664) );
AO22x1_ASAP7_75t_L g541 ( .A1(n_93), .A2(n_306), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g989 ( .A1(n_94), .A2(n_124), .B1(n_982), .B2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_95), .A2(n_168), .B1(n_645), .B2(n_1192), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_96), .A2(n_114), .B1(n_626), .B2(n_818), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_97), .A2(n_142), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_98), .A2(n_310), .B1(n_558), .B2(n_693), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_99), .A2(n_112), .B1(n_407), .B2(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_100), .B(n_428), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_101), .A2(n_210), .B1(n_555), .B2(n_557), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_102), .A2(n_136), .B1(n_521), .B2(n_731), .Y(n_863) );
INVx1_ASAP7_75t_L g654 ( .A(n_103), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_104), .A2(n_190), .B1(n_508), .B2(n_630), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_105), .A2(n_319), .B1(n_543), .B2(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_106), .A2(n_118), .B1(n_504), .B2(n_539), .Y(n_662) );
INVx1_ASAP7_75t_L g968 ( .A(n_107), .Y(n_968) );
AND2x4_ASAP7_75t_L g971 ( .A(n_107), .B(n_366), .Y(n_971) );
INVx1_ASAP7_75t_SL g988 ( .A(n_107), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_110), .A2(n_340), .B1(n_504), .B2(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_111), .B(n_428), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_113), .B(n_592), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_115), .A2(n_792), .B(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_116), .A2(n_149), .B1(n_966), .B2(n_970), .Y(n_1014) );
AOI33xp33_ASAP7_75t_R g1198 ( .A1(n_117), .A2(n_243), .A3(n_409), .B1(n_419), .B2(n_1199), .B3(n_1220), .Y(n_1198) );
INVx1_ASAP7_75t_L g762 ( .A(n_119), .Y(n_762) );
INVx1_ASAP7_75t_L g878 ( .A(n_120), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_121), .A2(n_315), .B1(n_583), .B2(n_586), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_122), .A2(n_257), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_123), .A2(n_256), .B1(n_517), .B2(n_518), .Y(n_779) );
AO22x1_ASAP7_75t_L g506 ( .A1(n_125), .A2(n_308), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_126), .A2(n_232), .B1(n_381), .B2(n_405), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_128), .A2(n_214), .B1(n_486), .B2(n_507), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_130), .A2(n_248), .B1(n_649), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_131), .A2(n_159), .B1(n_483), .B2(n_615), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_132), .A2(n_252), .B1(n_577), .B2(n_582), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_133), .A2(n_180), .B1(n_647), .B2(n_649), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_134), .A2(n_223), .B1(n_686), .B2(n_688), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_138), .A2(n_291), .B1(n_594), .B2(n_597), .C(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_140), .A2(n_334), .B1(n_776), .B2(n_777), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_141), .A2(n_279), .B1(n_382), .B2(n_608), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_145), .B(n_428), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_146), .A2(n_267), .B1(n_504), .B2(n_520), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_147), .A2(n_294), .B1(n_476), .B2(n_546), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_148), .A2(n_348), .B1(n_504), .B2(n_520), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_151), .A2(n_165), .B1(n_542), .B2(n_630), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_152), .A2(n_322), .B1(n_498), .B2(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g404 ( .A(n_153), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_153), .B(n_203), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_153), .B(n_421), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_154), .B(n_274), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_155), .A2(n_217), .B1(n_1003), .B2(n_1094), .Y(n_1093) );
XNOR2x1_ASAP7_75t_L g572 ( .A(n_156), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g939 ( .A(n_157), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_158), .A2(n_164), .B1(n_505), .B2(n_508), .Y(n_695) );
INVx1_ASAP7_75t_L g908 ( .A(n_160), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_161), .B(n_594), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_162), .A2(n_167), .B1(n_483), .B2(n_615), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_163), .A2(n_173), .B1(n_576), .B2(n_585), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_166), .A2(n_270), .B1(n_548), .B2(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_169), .B(n_397), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_171), .A2(n_332), .B1(n_507), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_172), .A2(n_314), .B1(n_686), .B2(n_688), .Y(n_768) );
XNOR2x1_ASAP7_75t_L g678 ( .A(n_175), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_176), .A2(n_356), .B1(n_475), .B2(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g913 ( .A(n_179), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_181), .Y(n_829) );
INVx1_ASAP7_75t_L g953 ( .A(n_182), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_183), .A2(n_222), .B1(n_476), .B2(n_546), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_184), .B(n_514), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_185), .A2(n_349), .B1(n_576), .B2(n_577), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_186), .A2(n_324), .B1(n_557), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_187), .A2(n_359), .B1(n_557), .B2(n_558), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_188), .A2(n_226), .B1(n_582), .B2(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g847 ( .A(n_189), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_191), .A2(n_352), .B1(n_594), .B2(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g918 ( .A(n_192), .Y(n_918) );
INVx1_ASAP7_75t_L g605 ( .A(n_193), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_195), .A2(n_307), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_196), .A2(n_239), .B1(n_482), .B2(n_485), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_197), .A2(n_271), .B1(n_582), .B2(n_585), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_198), .A2(n_230), .B1(n_973), .B2(n_980), .Y(n_979) );
XOR2x2_ASAP7_75t_L g1185 ( .A(n_198), .B(n_1186), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_198), .A2(n_1205), .B1(n_1207), .B2(n_1211), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_200), .A2(n_269), .B1(n_576), .B2(n_597), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_201), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_202), .B(n_682), .Y(n_769) );
INVx1_ASAP7_75t_L g391 ( .A(n_203), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_204), .A2(n_343), .B1(n_579), .B2(n_580), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_205), .A2(n_321), .B1(n_557), .B2(n_752), .Y(n_796) );
INVx1_ASAP7_75t_L g492 ( .A(n_206), .Y(n_492) );
OAI222xp33_ASAP7_75t_L g509 ( .A1(n_206), .A2(n_510), .B1(n_516), .B2(n_519), .C1(n_1216), .C2(n_1217), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_206), .B(n_519), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_207), .Y(n_831) );
INVx1_ASAP7_75t_L g736 ( .A(n_212), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_212), .A2(n_303), .B1(n_973), .B2(n_976), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_213), .A2(n_341), .B1(n_582), .B2(n_583), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_216), .A2(n_241), .B1(n_486), .B2(n_507), .Y(n_698) );
XNOR2x1_ASAP7_75t_L g377 ( .A(n_219), .B(n_378), .Y(n_377) );
XNOR2x2_ASAP7_75t_SL g529 ( .A(n_219), .B(n_378), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_219), .A2(n_254), .B1(n_973), .B2(n_976), .Y(n_972) );
INVx1_ASAP7_75t_L g643 ( .A(n_221), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_225), .B(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_227), .A2(n_280), .B1(n_539), .B2(n_801), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_228), .A2(n_247), .B1(n_495), .B2(n_641), .C(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_231), .A2(n_298), .B1(n_973), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_233), .A2(n_292), .B1(n_970), .B2(n_993), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_235), .A2(n_347), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_237), .A2(n_326), .B1(n_966), .B2(n_982), .Y(n_981) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_238), .A2(n_535), .B(n_566), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_238), .B(n_538), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_240), .A2(n_325), .B1(n_592), .B2(n_597), .C(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_242), .A2(n_250), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g894 ( .A(n_249), .Y(n_894) );
INVx1_ASAP7_75t_L g441 ( .A(n_251), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_255), .A2(n_285), .B1(n_483), .B2(n_540), .Y(n_862) );
INVx1_ASAP7_75t_L g668 ( .A(n_258), .Y(n_668) );
INVx1_ASAP7_75t_L g787 ( .A(n_259), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_259), .B(n_802), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_260), .A2(n_639), .B(n_642), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_261), .A2(n_301), .B1(n_504), .B2(n_520), .Y(n_696) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_262), .Y(n_371) );
AND2x4_ASAP7_75t_L g974 ( .A(n_262), .B(n_975), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_264), .A2(n_273), .B1(n_585), .B2(n_586), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_265), .Y(n_826) );
XNOR2x1_ASAP7_75t_L g600 ( .A(n_268), .B(n_601), .Y(n_600) );
AOI211x1_ASAP7_75t_L g904 ( .A1(n_272), .A2(n_905), .B(n_907), .C(n_915), .Y(n_904) );
INVx1_ASAP7_75t_L g402 ( .A(n_274), .Y(n_402) );
INVxp67_ASAP7_75t_L g440 ( .A(n_274), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_276), .A2(n_351), .B1(n_465), .B2(n_470), .Y(n_464) );
INVx1_ASAP7_75t_L g562 ( .A(n_277), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_282), .A2(n_318), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g366 ( .A(n_283), .Y(n_366) );
INVx1_ASAP7_75t_SL g812 ( .A(n_289), .Y(n_812) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_289), .B(n_838), .C(n_839), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_290), .A2(n_335), .B1(n_412), .B2(n_416), .Y(n_795) );
INVx1_ASAP7_75t_L g849 ( .A(n_293), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_297), .A2(n_299), .B1(n_589), .B2(n_595), .Y(n_928) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_300), .A2(n_597), .B(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_304), .A2(n_320), .B1(n_382), .B2(n_555), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_305), .A2(n_316), .B1(n_597), .B2(n_706), .Y(n_927) );
INVx1_ASAP7_75t_L g794 ( .A(n_311), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_312), .B(n_514), .Y(n_1193) );
XOR2xp5_ASAP7_75t_L g700 ( .A(n_317), .B(n_701), .Y(n_700) );
XOR2xp5_ASAP7_75t_L g755 ( .A(n_317), .B(n_701), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_327), .A2(n_333), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g733 ( .A(n_331), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_336), .A2(n_355), .B1(n_592), .B2(n_645), .Y(n_929) );
AO22x2_ASAP7_75t_L g841 ( .A1(n_338), .A2(n_842), .B1(n_843), .B2(n_844), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_338), .Y(n_842) );
AND2x2_ASAP7_75t_L g814 ( .A(n_339), .B(n_772), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_345), .A2(n_1208), .B1(n_1209), .B2(n_1210), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_345), .Y(n_1208) );
INVx1_ASAP7_75t_L g917 ( .A(n_346), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_353), .A2(n_358), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_372), .B(n_958), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
BUFx4_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .C(n_371), .Y(n_363) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_364), .B(n_1202), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_364), .B(n_1203), .Y(n_1206) );
AOI21xp5_ASAP7_75t_L g1214 ( .A1(n_364), .A2(n_371), .B(n_988), .Y(n_1214) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AO21x1_ASAP7_75t_L g1212 ( .A1(n_365), .A2(n_1213), .B(n_1214), .Y(n_1212) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g967 ( .A(n_366), .B(n_968), .Y(n_967) );
AND3x4_ASAP7_75t_L g987 ( .A(n_366), .B(n_974), .C(n_988), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_367), .B(n_1203), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_368), .A2(n_447), .B(n_448), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g1203 ( .A(n_371), .Y(n_1203) );
XNOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_757), .Y(n_372) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_674), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_530), .B1(n_672), .B2(n_673), .Y(n_374) );
INVx1_ASAP7_75t_L g673 ( .A(n_375), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_489), .B1(n_490), .B2(n_529), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_450), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_410), .C(n_426), .Y(n_379) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g848 ( .A(n_382), .Y(n_848) );
BUFx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_383), .Y(n_495) );
INVx1_ASAP7_75t_L g687 ( .A(n_383), .Y(n_687) );
BUFx3_ASAP7_75t_L g891 ( .A(n_383), .Y(n_891) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_394), .Y(n_383) );
AND2x4_ASAP7_75t_L g413 ( .A(n_384), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g592 ( .A(n_384), .B(n_414), .Y(n_592) );
AND2x4_ASAP7_75t_L g597 ( .A(n_384), .B(n_394), .Y(n_597) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
AND2x2_ASAP7_75t_L g409 ( .A(n_385), .B(n_389), .Y(n_409) );
AND2x2_ASAP7_75t_L g438 ( .A(n_385), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g456 ( .A(n_385), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_386), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp33_ASAP7_75t_L g390 ( .A(n_387), .B(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g397 ( .A(n_387), .Y(n_397) );
NAND2xp33_ASAP7_75t_L g403 ( .A(n_387), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
AND2x4_ASAP7_75t_L g455 ( .A(n_388), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_391), .B(n_423), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_393), .A2(n_425), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g408 ( .A(n_394), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g477 ( .A(n_394), .B(n_455), .Y(n_477) );
AND2x4_ASAP7_75t_L g579 ( .A(n_394), .B(n_455), .Y(n_579) );
AND2x4_ASAP7_75t_L g589 ( .A(n_394), .B(n_409), .Y(n_589) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_399), .Y(n_394) );
INVx2_ASAP7_75t_L g415 ( .A(n_395), .Y(n_415) );
AND2x2_ASAP7_75t_L g434 ( .A(n_395), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g468 ( .A(n_395), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_397), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g421 ( .A(n_397), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_398), .B(n_420), .C(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g414 ( .A(n_399), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_406), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_408), .Y(n_557) );
INVx2_ASAP7_75t_L g637 ( .A(n_408), .Y(n_637) );
AND2x2_ASAP7_75t_L g430 ( .A(n_409), .B(n_414), .Y(n_430) );
AND2x2_ASAP7_75t_L g467 ( .A(n_409), .B(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g472 ( .A(n_409), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g549 ( .A(n_409), .B(n_468), .Y(n_549) );
AND2x4_ASAP7_75t_L g576 ( .A(n_409), .B(n_468), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_409), .B(n_457), .Y(n_577) );
AND2x2_ASAP7_75t_L g594 ( .A(n_409), .B(n_414), .Y(n_594) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g514 ( .A(n_413), .Y(n_514) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_413), .Y(n_554) );
INVx2_ASAP7_75t_L g648 ( .A(n_413), .Y(n_648) );
BUFx8_ASAP7_75t_SL g690 ( .A(n_413), .Y(n_690) );
INVx2_ASAP7_75t_L g767 ( .A(n_413), .Y(n_767) );
AND2x4_ASAP7_75t_L g418 ( .A(n_414), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g480 ( .A(n_414), .B(n_455), .Y(n_480) );
AND2x4_ASAP7_75t_L g580 ( .A(n_414), .B(n_455), .Y(n_580) );
AND2x4_ASAP7_75t_L g595 ( .A(n_414), .B(n_419), .Y(n_595) );
INVx1_ASAP7_75t_L g916 ( .A(n_416), .Y(n_916) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g608 ( .A(n_417), .Y(n_608) );
INVx3_ASAP7_75t_L g649 ( .A(n_417), .Y(n_649) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_418), .Y(n_515) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_418), .Y(n_555) );
AND2x4_ASAP7_75t_L g463 ( .A(n_419), .B(n_457), .Y(n_463) );
AND2x4_ASAP7_75t_L g488 ( .A(n_419), .B(n_468), .Y(n_488) );
AND2x4_ASAP7_75t_L g585 ( .A(n_419), .B(n_468), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_419), .B(n_457), .Y(n_586) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_424), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g607 ( .A(n_429), .Y(n_607) );
INVx2_ASAP7_75t_L g641 ( .A(n_429), .Y(n_641) );
INVx2_ASAP7_75t_L g910 ( .A(n_429), .Y(n_910) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g498 ( .A(n_430), .Y(n_498) );
INVx2_ASAP7_75t_L g684 ( .A(n_430), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_441), .B(n_442), .Y(n_431) );
INVx2_ASAP7_75t_L g512 ( .A(n_432), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_432), .A2(n_643), .B(n_644), .Y(n_642) );
INVx4_ASAP7_75t_L g692 ( .A(n_432), .Y(n_692) );
INVx2_ASAP7_75t_L g752 ( .A(n_432), .Y(n_752) );
INVx2_ASAP7_75t_L g771 ( .A(n_432), .Y(n_771) );
INVx5_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_433), .Y(n_558) );
BUFx2_ASAP7_75t_L g610 ( .A(n_433), .Y(n_610) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_433), .Y(n_1190) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_438), .Y(n_433) );
AND2x4_ASAP7_75t_L g590 ( .A(n_434), .B(n_438), .Y(n_590) );
AND2x2_ASAP7_75t_L g706 ( .A(n_434), .B(n_438), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g447 ( .A(n_436), .Y(n_447) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_444), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g693 ( .A(n_444), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_444), .B(n_894), .Y(n_893) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g773 ( .A(n_445), .Y(n_773) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_446), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_464), .C(n_474), .D(n_481), .Y(n_450) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_454), .Y(n_540) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_454), .Y(n_615) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
AND2x4_ASAP7_75t_L g484 ( .A(n_455), .B(n_468), .Y(n_484) );
AND2x4_ASAP7_75t_L g582 ( .A(n_455), .B(n_468), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_455), .B(n_473), .Y(n_583) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g473 ( .A(n_458), .Y(n_473) );
INVx1_ASAP7_75t_L g469 ( .A(n_459), .Y(n_469) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g505 ( .A(n_462), .Y(n_505) );
INVx5_ASAP7_75t_L g543 ( .A(n_462), .Y(n_543) );
INVx3_ASAP7_75t_L g743 ( .A(n_462), .Y(n_743) );
INVx1_ASAP7_75t_L g777 ( .A(n_462), .Y(n_777) );
INVx2_ASAP7_75t_L g943 ( .A(n_462), .Y(n_943) );
INVx6_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx12f_ASAP7_75t_L g630 ( .A(n_463), .Y(n_630) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_466), .Y(n_781) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx8_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_468), .Y(n_1199) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx12f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_472), .Y(n_508) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_472), .Y(n_742) );
BUFx3_ASAP7_75t_L g776 ( .A(n_472), .Y(n_776) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx12f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
INVx3_ASAP7_75t_L g746 ( .A(n_477), .Y(n_746) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx5_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
INVx1_ASAP7_75t_L g627 ( .A(n_480), .Y(n_627) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx12f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_484), .Y(n_520) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_484), .Y(n_539) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g521 ( .A(n_487), .Y(n_521) );
INVx4_ASAP7_75t_L g550 ( .A(n_487), .Y(n_550) );
INVx4_ASAP7_75t_L g632 ( .A(n_487), .Y(n_632) );
INVx2_ASAP7_75t_SL g661 ( .A(n_487), .Y(n_661) );
INVx1_ASAP7_75t_L g782 ( .A(n_487), .Y(n_782) );
INVx1_ASAP7_75t_L g801 ( .A(n_487), .Y(n_801) );
INVx8_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_522), .Y(n_490) );
AOI21x1_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_509), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_501), .Y(n_493) );
BUFx2_ASAP7_75t_L g523 ( .A(n_494), .Y(n_523) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g856 ( .A1(n_497), .A2(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g527 ( .A(n_503), .B(n_516), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_506), .Y(n_528) );
INVx1_ASAP7_75t_L g526 ( .A(n_510), .Y(n_526) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
NAND4xp75_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .C(n_527), .D(n_528), .Y(n_522) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g672 ( .A(n_530), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_619), .B2(n_671), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OA22x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_570), .B1(n_571), .B2(n_618), .Y(n_532) );
INVx2_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_551), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .C(n_544), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_541), .B(n_559), .C(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_544), .B(n_552), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx4f_ASAP7_75t_L g731 ( .A(n_549), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_559), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx2_ASAP7_75t_L g853 ( .A(n_554), .Y(n_853) );
INVx3_ASAP7_75t_L g855 ( .A(n_555), .Y(n_855) );
INVx3_ASAP7_75t_L g850 ( .A(n_557), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_563), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g726 ( .A(n_563), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_563), .B(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_563), .B(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_563), .B(n_953), .Y(n_952) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_564), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g645 ( .A(n_564), .Y(n_645) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_564), .Y(n_669) );
INVx2_ASAP7_75t_SL g708 ( .A(n_564), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_600), .Y(n_571) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_572), .A2(n_652), .B1(n_653), .B2(n_670), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_572), .Y(n_652) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_587), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .C(n_581), .D(n_584), .Y(n_574) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .C(n_593), .D(n_596), .Y(n_587) );
INVx2_ASAP7_75t_L g832 ( .A(n_589), .Y(n_832) );
INVx4_ASAP7_75t_L g825 ( .A(n_590), .Y(n_825) );
INVx2_ASAP7_75t_L g827 ( .A(n_595), .Y(n_827) );
INVx2_ASAP7_75t_L g830 ( .A(n_597), .Y(n_830) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_602), .B(n_611), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .C(n_609), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .C(n_616), .D(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g671 ( .A(n_619), .Y(n_671) );
XNOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_651), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
XOR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_650), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_633), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .C(n_629), .D(n_631), .Y(n_623) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_638), .C(n_646), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g688 ( .A(n_636), .Y(n_688) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g670 ( .A(n_653), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND4xp75_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .C(n_663), .D(n_666), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g859 ( .A(n_669), .Y(n_859) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AO22x1_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_716), .B2(n_756), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AO22x2_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_699), .B1(n_714), .B2(n_715), .Y(n_677) );
INVx2_ASAP7_75t_L g714 ( .A(n_678), .Y(n_714) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_694), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .C(n_689), .D(n_691), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g1192 ( .A(n_684), .Y(n_1192) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g792 ( .A(n_687), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .C(n_697), .D(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g715 ( .A(n_699), .Y(n_715) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_709), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .C(n_705), .D(n_707), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .C(n_712), .D(n_713), .Y(n_709) );
INVx2_ASAP7_75t_SL g756 ( .A(n_716), .Y(n_756) );
XNOR2x1_ASAP7_75t_L g716 ( .A(n_717), .B(n_734), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
XOR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_733), .Y(n_719) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_727), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .C(n_724), .D(n_725), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .C(n_730), .D(n_732), .Y(n_727) );
XNOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_754), .Y(n_734) );
XNOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_747), .Y(n_737) );
NAND4xp25_ASAP7_75t_SL g738 ( .A(n_739), .B(n_740), .C(n_741), .D(n_744), .Y(n_738) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g818 ( .A(n_746), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .C(n_753), .Y(n_747) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_872), .B2(n_873), .Y(n_757) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_783), .B1(n_870), .B2(n_871), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_761), .Y(n_870) );
XNOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_774), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_765), .B(n_768), .C(n_769), .D(n_770), .Y(n_764) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
OAI21xp5_ASAP7_75t_SL g912 ( .A1(n_767), .A2(n_913), .B(n_914), .Y(n_912) );
INVx4_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND4xp25_ASAP7_75t_L g774 ( .A(n_775), .B(n_778), .C(n_779), .D(n_780), .Y(n_774) );
INVx1_ASAP7_75t_L g871 ( .A(n_783), .Y(n_871) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AO22x2_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_840), .B1(n_867), .B2(n_868), .Y(n_784) );
INVx1_ASAP7_75t_L g867 ( .A(n_785), .Y(n_867) );
XNOR2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_808), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B(n_805), .Y(n_786) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_797), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_789), .B(n_806), .C(n_807), .Y(n_805) );
AND4x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .C(n_795), .D(n_796), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_802), .Y(n_797) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_798), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NAND2x1_ASAP7_75t_L g808 ( .A(n_809), .B(n_833), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_815), .C(n_820), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B1(n_813), .B2(n_1218), .Y(n_810) );
INVx1_ASAP7_75t_L g838 ( .A(n_811), .Y(n_838) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_812), .B(n_816), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_812), .A2(n_821), .B1(n_822), .B2(n_1219), .Y(n_820) );
INVx1_ASAP7_75t_L g835 ( .A(n_813), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_816), .B(n_834), .C(n_837), .Y(n_833) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .Y(n_816) );
INVx1_ASAP7_75t_L g839 ( .A(n_821), .Y(n_839) );
INVx1_ASAP7_75t_L g836 ( .A(n_822), .Y(n_836) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_828), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g869 ( .A(n_841), .Y(n_869) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_860), .Y(n_844) );
NOR3xp33_ASAP7_75t_SL g845 ( .A(n_846), .B(n_851), .C(n_856), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B1(n_849), .B2(n_850), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B1(n_895), .B2(n_957), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
BUFx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
XNOR2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
NOR4xp75_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .C(n_886), .D(n_889), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
NAND2xp5_ASAP7_75t_SL g889 ( .A(n_890), .B(n_892), .Y(n_889) );
INVx2_ASAP7_75t_L g906 ( .A(n_891), .Y(n_906) );
INVx2_ASAP7_75t_SL g957 ( .A(n_895), .Y(n_957) );
OA22x2_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_920), .B1(n_921), .B2(n_956), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g956 ( .A(n_897), .Y(n_956) );
XNOR2x1_ASAP7_75t_L g897 ( .A(n_898), .B(n_919), .Y(n_897) );
NAND2x1_ASAP7_75t_L g898 ( .A(n_899), .B(n_904), .Y(n_898) );
AND4x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .C(n_902), .D(n_903), .Y(n_899) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .B(n_911), .Y(n_907) );
INVx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
AOI22x1_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_936), .B1(n_954), .B2(n_955), .Y(n_921) );
INVx2_ASAP7_75t_L g955 ( .A(n_922), .Y(n_955) );
INVx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
XNOR2x1_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
OR2x2_ASAP7_75t_L g925 ( .A(n_926), .B(n_931), .Y(n_925) );
NAND4xp25_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .C(n_929), .D(n_930), .Y(n_926) );
NAND4xp25_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .C(n_934), .D(n_935), .Y(n_931) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
BUFx2_ASAP7_75t_L g954 ( .A(n_937), .Y(n_954) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_940), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_939), .Y(n_938) );
NOR2x1_ASAP7_75t_L g940 ( .A(n_941), .B(n_947), .Y(n_940) );
NAND4xp25_ASAP7_75t_L g941 ( .A(n_942), .B(n_944), .C(n_945), .D(n_946), .Y(n_941) );
NAND4xp25_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .C(n_950), .D(n_951), .Y(n_947) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_1179), .B1(n_1181), .B2(n_1200), .C(n_1204), .Y(n_958) );
AOI211xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_1090), .B(n_1097), .C(n_1146), .Y(n_959) );
NAND5xp2_ASAP7_75t_L g960 ( .A(n_961), .B(n_1035), .C(n_1060), .D(n_1072), .E(n_1077), .Y(n_960) );
AOI211xp5_ASAP7_75t_SL g961 ( .A1(n_962), .A2(n_994), .B(n_998), .C(n_1027), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_977), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_963), .B(n_1026), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_963), .B(n_1034), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_963), .B(n_1079), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_963), .B(n_1131), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_963), .B(n_1164), .Y(n_1163) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx3_ASAP7_75t_L g1021 ( .A(n_964), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_964), .B(n_1042), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_964), .B(n_1000), .Y(n_1067) );
INVx2_ASAP7_75t_L g1100 ( .A(n_964), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_964), .B(n_1071), .Y(n_1109) );
NOR3xp33_ASAP7_75t_L g1156 ( .A(n_964), .B(n_1024), .C(n_1092), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g1178 ( .A(n_964), .B(n_1082), .Y(n_1178) );
AND2x2_ASAP7_75t_L g964 ( .A(n_965), .B(n_972), .Y(n_964) );
AND2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_969), .Y(n_966) );
AND2x4_ASAP7_75t_L g973 ( .A(n_967), .B(n_974), .Y(n_973) );
AND2x2_ASAP7_75t_L g990 ( .A(n_967), .B(n_969), .Y(n_990) );
AND2x4_ASAP7_75t_L g993 ( .A(n_967), .B(n_969), .Y(n_993) );
AND2x2_ASAP7_75t_L g970 ( .A(n_969), .B(n_971), .Y(n_970) );
AND2x2_ASAP7_75t_L g982 ( .A(n_969), .B(n_971), .Y(n_982) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_969), .B(n_971), .Y(n_1006) );
AND2x4_ASAP7_75t_L g976 ( .A(n_971), .B(n_974), .Y(n_976) );
AND2x4_ASAP7_75t_L g980 ( .A(n_971), .B(n_974), .Y(n_980) );
INVx3_ASAP7_75t_L g1095 ( .A(n_973), .Y(n_1095) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_976), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_977), .B(n_1032), .Y(n_1114) );
AND2x2_ASAP7_75t_L g977 ( .A(n_978), .B(n_983), .Y(n_977) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_978), .B(n_1020), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_978), .B(n_1023), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_978), .B(n_1037), .Y(n_1036) );
CKINVDCx6p67_ASAP7_75t_R g1042 ( .A(n_978), .Y(n_1042) );
AOI32xp33_ASAP7_75t_L g1077 ( .A1(n_978), .A2(n_1078), .A3(n_1080), .B1(n_1083), .B2(n_1087), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_978), .B(n_984), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_978), .B(n_1017), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_978), .B(n_1024), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_978), .B(n_985), .Y(n_1139) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_981), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_983), .B(n_1019), .Y(n_1063) );
INVx1_ASAP7_75t_L g1082 ( .A(n_983), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_983), .B(n_1042), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_983), .B(n_1059), .Y(n_1113) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_991), .Y(n_983) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_984), .A2(n_1032), .B1(n_1127), .B2(n_1152), .C(n_1153), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_984), .B(n_1042), .Y(n_1164) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_985), .B(n_991), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_985), .B(n_1024), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_985), .B(n_991), .Y(n_1038) );
AND2x2_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .Y(n_985) );
INVx1_ASAP7_75t_L g1024 ( .A(n_991), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_991), .B(n_1019), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_991), .B(n_1042), .Y(n_1136) );
INVxp67_ASAP7_75t_L g1007 ( .A(n_994), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_994), .B(n_1013), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_994), .B(n_1012), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_994), .B(n_1013), .Y(n_1071) );
INVx2_ASAP7_75t_L g1075 ( .A(n_994), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_994), .B(n_1000), .Y(n_1086) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_995), .B(n_1013), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_995), .B(n_1001), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
OAI21xp33_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1008), .B(n_1022), .Y(n_998) );
INVx1_ASAP7_75t_L g1134 ( .A(n_999), .Y(n_1134) );
AOI21xp33_ASAP7_75t_SL g1166 ( .A1(n_999), .A2(n_1149), .B(n_1167), .Y(n_1166) );
OR2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1007), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_1000), .B(n_1026), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1000), .B(n_1032), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1000), .B(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1000), .B(n_1075), .Y(n_1074) );
AOI32xp33_ASAP7_75t_L g1124 ( .A1(n_1000), .A2(n_1078), .A3(n_1125), .B1(n_1126), .B2(n_1128), .Y(n_1124) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1000), .Y(n_1150) );
INVx4_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1001), .B(n_1010), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1145 ( .A(n_1001), .B(n_1092), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1001), .B(n_1079), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_1001), .B(n_1052), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1001), .B(n_1032), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1005), .Y(n_1001) );
INVx2_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1007), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1016), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_1009), .B(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1011), .Y(n_1057) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1012), .Y(n_1032) );
INVx4_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1013), .B(n_1100), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1016), .B(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1019), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1017), .B(n_1042), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1017), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1069 ( .A(n_1018), .B(n_1020), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1019), .B(n_1038), .Y(n_1127) );
NOR2x1_ASAP7_75t_L g1061 ( .A(n_1020), .B(n_1051), .Y(n_1061) );
A2O1A1Ixp33_ASAP7_75t_L g1103 ( .A1(n_1020), .A2(n_1026), .B(n_1104), .C(n_1106), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g1110 ( .A1(n_1020), .A2(n_1086), .B1(n_1111), .B2(n_1116), .C(n_1121), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1020), .B(n_1046), .Y(n_1152) );
INVx3_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1021), .B(n_1038), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1021), .B(n_1089), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1021), .B(n_1046), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1025), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1023), .B(n_1042), .Y(n_1051) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1023), .Y(n_1081) );
O2A1O1Ixp33_ASAP7_75t_L g1066 ( .A1(n_1024), .A2(n_1067), .B(n_1068), .C(n_1070), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1024), .B(n_1042), .Y(n_1108) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1026), .Y(n_1154) );
AOI21xp33_ASAP7_75t_SL g1175 ( .A1(n_1026), .A2(n_1176), .B(n_1177), .Y(n_1175) );
AOI21xp33_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1030), .B(n_1033), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_1031), .A2(n_1050), .B1(n_1061), .B2(n_1159), .Y(n_1158) );
AOI32xp33_ASAP7_75t_L g1141 ( .A1(n_1032), .A2(n_1063), .A3(n_1104), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1032), .B(n_1163), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1033), .B(n_1104), .Y(n_1118) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
O2A1O1Ixp33_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1039), .B(n_1043), .C(n_1044), .Y(n_1035) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1038), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1038), .B(n_1059), .Y(n_1174) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1042), .B(n_1069), .Y(n_1068) );
A2O1A1Ixp33_ASAP7_75t_SL g1129 ( .A1(n_1043), .A2(n_1091), .B(n_1130), .C(n_1132), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1048), .B1(n_1049), .B2(n_1052), .C(n_1053), .Y(n_1044) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1050), .B(n_1071), .Y(n_1106) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1052), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_1052), .A2(n_1117), .B1(n_1119), .B2(n_1120), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1058), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1055), .B(n_1113), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1126 ( .A(n_1055), .B(n_1127), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1055), .Y(n_1172) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1056), .Y(n_1085) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_1057), .Y(n_1123) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1058), .Y(n_1176) );
O2A1O1Ixp33_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1062), .B(n_1064), .C(n_1066), .Y(n_1060) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1069), .Y(n_1142) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1076), .Y(n_1073) );
INVx3_ASAP7_75t_SL g1102 ( .A(n_1075), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1075), .B(n_1091), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1085), .Y(n_1144) );
INVxp33_ASAP7_75t_SL g1087 ( .A(n_1088), .Y(n_1087) );
OAI211xp5_ASAP7_75t_L g1097 ( .A1(n_1090), .A2(n_1098), .B(n_1110), .C(n_1137), .Y(n_1097) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1091), .B(n_1150), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_1092), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1096), .Y(n_1092) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1094), .Y(n_1180) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AOI211xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1102), .B(n_1103), .C(n_1107), .Y(n_1098) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1099), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_1099), .A2(n_1148), .B1(n_1151), .B2(n_1154), .Y(n_1147) );
OAI31xp33_ASAP7_75t_L g1155 ( .A1(n_1099), .A2(n_1105), .A3(n_1156), .B(n_1157), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1101), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1100), .B(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1101), .Y(n_1153) );
OAI211xp5_ASAP7_75t_SL g1121 ( .A1(n_1102), .A2(n_1122), .B(n_1124), .C(n_1129), .Y(n_1121) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1109), .Y(n_1107) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1108), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1114), .C(n_1115), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1160 ( .A1(n_1113), .A2(n_1148), .B1(n_1161), .B2(n_1165), .C(n_1166), .Y(n_1160) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_1133), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
A2O1A1Ixp33_ASAP7_75t_SL g1137 ( .A1(n_1138), .A2(n_1140), .B(n_1141), .C(n_1145), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1139), .B(n_1168), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NAND5xp2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1155), .C(n_1158), .D(n_1160), .E(n_1170), .Y(n_1146) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
A2O1A1Ixp33_ASAP7_75t_L g1170 ( .A1(n_1150), .A2(n_1171), .B(n_1173), .C(n_1175), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1186), .Y(n_1210) );
NOR2x1_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1194), .Y(n_1186) );
NAND4xp25_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .C(n_1191), .D(n_1193), .Y(n_1187) );
NAND4xp25_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .C(n_1197), .D(n_1198), .Y(n_1194) );
CKINVDCx16_ASAP7_75t_R g1200 ( .A(n_1201), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
endmodule