module real_aes_146_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_0), .A2(n_108), .B1(n_282), .B2(n_283), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_1), .B(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_2), .A2(n_72), .B1(n_292), .B2(n_316), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_3), .Y(n_655) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_4), .A2(n_157), .B1(n_246), .B2(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g588 ( .A(n_4), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_5), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_6), .A2(n_14), .B1(n_422), .B2(n_547), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_7), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_8), .A2(n_49), .B1(n_359), .B2(n_361), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_9), .A2(n_117), .B1(n_333), .B2(n_336), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g266 ( .A1(n_10), .A2(n_199), .B1(n_267), .B2(n_270), .Y(n_266) );
AOI22x1_ASAP7_75t_L g318 ( .A1(n_11), .A2(n_94), .B1(n_294), .B2(n_319), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_12), .A2(n_191), .B1(n_282), .B2(n_283), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_13), .B(n_457), .Y(n_456) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_15), .A2(n_46), .B1(n_246), .B2(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_15), .B(n_587), .Y(n_586) );
AO222x2_ASAP7_75t_L g562 ( .A1(n_16), .A2(n_45), .B1(n_176), .B2(n_242), .C1(n_270), .C2(n_311), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_17), .A2(n_177), .B1(n_282), .B2(n_283), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_18), .A2(n_114), .B1(n_311), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_19), .A2(n_153), .B1(n_345), .B2(n_499), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_20), .B(n_297), .Y(n_296) );
XNOR2xp5_ASAP7_75t_L g323 ( .A(n_20), .B(n_297), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_21), .A2(n_22), .B1(n_294), .B2(n_295), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_23), .A2(n_187), .B1(n_261), .B2(n_306), .Y(n_565) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_24), .A2(n_134), .B1(n_190), .B2(n_365), .C1(n_368), .C2(n_371), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_25), .A2(n_93), .B1(n_294), .B2(n_295), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_26), .A2(n_173), .B1(n_354), .B2(n_436), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g308 ( .A1(n_27), .A2(n_205), .B1(n_270), .B2(n_309), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_28), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_29), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g411 ( .A1(n_30), .A2(n_109), .B1(n_221), .B2(n_365), .C1(n_412), .C2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_31), .A2(n_36), .B1(n_333), .B2(n_385), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_32), .A2(n_97), .B1(n_401), .B2(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_33), .A2(n_63), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_34), .A2(n_83), .B1(n_267), .B2(n_273), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_35), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_37), .A2(n_214), .B1(n_354), .B2(n_356), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_38), .A2(n_215), .B1(n_607), .B2(n_609), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_39), .A2(n_207), .B1(n_371), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_169), .B1(n_306), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_41), .A2(n_119), .B1(n_336), .B2(n_496), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_42), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_43), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_44), .A2(n_138), .B1(n_341), .B2(n_345), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_47), .A2(n_77), .B1(n_273), .B2(n_311), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_48), .A2(n_104), .B1(n_328), .B2(n_331), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_50), .A2(n_106), .B1(n_390), .B2(n_391), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_51), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_52), .A2(n_209), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g281 ( .A1(n_53), .A2(n_189), .B1(n_282), .B2(n_283), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_54), .A2(n_140), .B1(n_286), .B2(n_294), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_55), .A2(n_110), .B1(n_390), .B2(n_391), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_56), .A2(n_194), .B1(n_288), .B2(n_292), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_57), .A2(n_141), .B1(n_422), .B2(n_447), .Y(n_666) );
INVx3_ASAP7_75t_L g246 ( .A(n_58), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_59), .A2(n_124), .B1(n_291), .B2(n_295), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_60), .A2(n_132), .B1(n_399), .B2(n_413), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_61), .A2(n_158), .B1(n_331), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_62), .A2(n_96), .B1(n_291), .B2(n_292), .Y(n_470) );
XOR2x2_ASAP7_75t_L g427 ( .A(n_64), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_65), .B(n_371), .Y(n_651) );
AO222x2_ASAP7_75t_L g241 ( .A1(n_66), .A2(n_115), .B1(n_137), .B2(n_242), .C1(n_258), .C2(n_261), .Y(n_241) );
INVx1_ASAP7_75t_L g373 ( .A(n_67), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_68), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_69), .A2(n_204), .B1(n_395), .B2(n_396), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_70), .A2(n_121), .B1(n_273), .B2(n_276), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_71), .Y(n_617) );
INVx1_ASAP7_75t_SL g247 ( .A(n_73), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_73), .B(n_102), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_74), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_75), .Y(n_302) );
INVx2_ASAP7_75t_L g228 ( .A(n_76), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_78), .A2(n_142), .B1(n_447), .B2(n_450), .Y(n_446) );
OA22x2_ASAP7_75t_L g378 ( .A1(n_79), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_79), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_80), .A2(n_120), .B1(n_331), .B2(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_81), .A2(n_200), .B1(n_291), .B2(n_292), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_82), .A2(n_186), .B1(n_418), .B2(n_420), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_84), .A2(n_91), .B1(n_356), .B2(n_401), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_85), .A2(n_216), .B1(n_390), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_86), .A2(n_155), .B1(n_347), .B2(n_350), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_87), .A2(n_156), .B1(n_341), .B2(n_522), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_88), .A2(n_116), .B1(n_601), .B2(n_603), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_89), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_90), .A2(n_112), .B1(n_401), .B2(n_402), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_92), .A2(n_179), .B1(n_319), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_95), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_98), .A2(n_113), .B1(n_328), .B2(n_418), .Y(n_439) );
XNOR2xp5_ASAP7_75t_SL g591 ( .A(n_99), .B(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_100), .A2(n_198), .B1(n_359), .B2(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_101), .A2(n_195), .B1(n_401), .B2(n_402), .Y(n_400) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_102), .A2(n_165), .B1(n_246), .B2(n_250), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_103), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_105), .A2(n_183), .B1(n_350), .B2(n_468), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_107), .A2(n_126), .B1(n_354), .B2(n_402), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_111), .A2(n_201), .B1(n_333), .B2(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_118), .A2(n_128), .B1(n_341), .B2(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g248 ( .A(n_122), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_123), .A2(n_151), .B1(n_333), .B2(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_125), .B(n_365), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_127), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_129), .A2(n_143), .B1(n_286), .B2(n_288), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_130), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g643 ( .A(n_131), .B(n_644), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_131), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_133), .A2(n_167), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_135), .A2(n_161), .B1(n_341), .B2(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_136), .A2(n_171), .B1(n_413), .B2(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g507 ( .A(n_139), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_144), .A2(n_159), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_145), .A2(n_152), .B1(n_384), .B2(n_385), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_146), .A2(n_208), .B1(n_413), .B2(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_147), .A2(n_206), .B1(n_333), .B2(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_148), .A2(n_184), .B1(n_319), .B2(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_149), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_150), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_154), .A2(n_172), .B1(n_270), .B2(n_309), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_160), .A2(n_178), .B1(n_286), .B2(n_295), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_162), .A2(n_218), .B1(n_387), .B2(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_163), .A2(n_559), .B1(n_560), .B2(n_573), .Y(n_558) );
INVx1_ASAP7_75t_L g573 ( .A(n_163), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_164), .A2(n_196), .B1(n_384), .B2(n_441), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_166), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_168), .A2(n_212), .B1(n_261), .B2(n_306), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_170), .A2(n_202), .B1(n_390), .B2(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g230 ( .A(n_174), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g584 ( .A(n_174), .Y(n_584) );
AO21x1_ASAP7_75t_L g675 ( .A1(n_174), .A2(n_226), .B(n_676), .Y(n_675) );
OA22x2_ASAP7_75t_L g406 ( .A1(n_175), .A2(n_407), .B1(n_408), .B2(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_175), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_180), .A2(n_223), .B(n_232), .C(n_590), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_181), .A2(n_213), .B1(n_361), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
AND2x2_ASAP7_75t_R g641 ( .A(n_182), .B(n_584), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_185), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_188), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_192), .A2(n_220), .B1(n_371), .B2(n_395), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_193), .A2(n_210), .B1(n_371), .B2(n_395), .Y(n_540) );
INVxp67_ASAP7_75t_L g227 ( .A(n_197), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_203), .A2(n_219), .B1(n_292), .B2(n_316), .Y(n_315) );
XNOR2x1_ASAP7_75t_L g534 ( .A(n_211), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_217), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVxp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_231), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g676 ( .A(n_231), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_477), .B1(n_579), .B2(n_580), .C(n_581), .Y(n_232) );
INVx1_ASAP7_75t_L g579 ( .A(n_233), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_374), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
XNOR2x1_ASAP7_75t_L g235 ( .A(n_236), .B(n_324), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_296), .B(n_322), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_237), .B(n_323), .Y(n_322) );
XNOR2x1_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_279), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_265), .Y(n_240) );
INVx2_ASAP7_75t_SL g301 ( .A(n_242), .Y(n_301) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_251), .Y(n_242) );
AND2x2_ASAP7_75t_L g270 ( .A(n_243), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g276 ( .A(n_243), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g311 ( .A(n_243), .B(n_277), .Y(n_311) );
AND2x4_ASAP7_75t_L g357 ( .A(n_243), .B(n_277), .Y(n_357) );
AND2x4_ASAP7_75t_L g363 ( .A(n_243), .B(n_271), .Y(n_363) );
AND2x2_ASAP7_75t_L g367 ( .A(n_243), .B(n_251), .Y(n_367) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_244), .Y(n_259) );
AND2x2_ASAP7_75t_L g263 ( .A(n_244), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g269 ( .A(n_244), .Y(n_269) );
OAI22x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g250 ( .A(n_246), .Y(n_250) );
INVx2_ASAP7_75t_L g254 ( .A(n_246), .Y(n_254) );
INVx1_ASAP7_75t_L g257 ( .A(n_246), .Y(n_257) );
INVx2_ASAP7_75t_L g264 ( .A(n_249), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_249), .B(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g284 ( .A(n_249), .Y(n_284) );
AND2x2_ASAP7_75t_L g286 ( .A(n_251), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g291 ( .A(n_251), .B(n_263), .Y(n_291) );
AND2x6_ASAP7_75t_L g294 ( .A(n_251), .B(n_268), .Y(n_294) );
AND2x2_ASAP7_75t_L g316 ( .A(n_251), .B(n_263), .Y(n_316) );
AND2x2_ASAP7_75t_L g330 ( .A(n_251), .B(n_268), .Y(n_330) );
AND2x4_ASAP7_75t_L g335 ( .A(n_251), .B(n_287), .Y(n_335) );
AND2x4_ASAP7_75t_L g349 ( .A(n_251), .B(n_263), .Y(n_349) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g260 ( .A(n_253), .B(n_256), .Y(n_260) );
AND2x4_ASAP7_75t_L g262 ( .A(n_253), .B(n_255), .Y(n_262) );
INVx1_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
INVxp67_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g274 ( .A(n_256), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_SL g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_259), .B(n_260), .Y(n_306) );
AND2x2_ASAP7_75t_L g372 ( .A(n_259), .B(n_260), .Y(n_372) );
AND2x4_ASAP7_75t_L g283 ( .A(n_260), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g292 ( .A(n_260), .B(n_287), .Y(n_292) );
AND2x4_ASAP7_75t_L g345 ( .A(n_260), .B(n_284), .Y(n_345) );
AND2x4_ASAP7_75t_L g351 ( .A(n_260), .B(n_287), .Y(n_351) );
INVx1_ASAP7_75t_SL g303 ( .A(n_261), .Y(n_303) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_L g267 ( .A(n_262), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g288 ( .A(n_262), .B(n_287), .Y(n_288) );
AND2x2_ASAP7_75t_L g309 ( .A(n_262), .B(n_268), .Y(n_309) );
AND2x4_ASAP7_75t_L g320 ( .A(n_262), .B(n_287), .Y(n_320) );
AND2x4_ASAP7_75t_L g360 ( .A(n_262), .B(n_268), .Y(n_360) );
AND2x2_ASAP7_75t_L g370 ( .A(n_262), .B(n_263), .Y(n_370) );
AND2x4_ASAP7_75t_L g273 ( .A(n_263), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g355 ( .A(n_263), .B(n_274), .Y(n_355) );
AND2x4_ASAP7_75t_L g287 ( .A(n_264), .B(n_269), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_272), .Y(n_265) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_268), .B(n_274), .Y(n_282) );
AND2x2_ASAP7_75t_L g342 ( .A(n_268), .B(n_274), .Y(n_342) );
AND2x6_ASAP7_75t_L g295 ( .A(n_274), .B(n_287), .Y(n_295) );
AND2x4_ASAP7_75t_L g338 ( .A(n_274), .B(n_287), .Y(n_338) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_275), .Y(n_278) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_289), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_298), .B(n_312), .Y(n_297) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_299), .B(n_307), .Y(n_298) );
OAI222xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_302), .B2(n_303), .C1(n_304), .C2(n_305), .Y(n_299) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_301), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_303), .Y(n_513) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx2_ASAP7_75t_L g618 ( .A(n_319), .Y(n_618) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
XOR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_373), .Y(n_324) );
NAND4xp75_ASAP7_75t_L g325 ( .A(n_326), .B(n_339), .C(n_352), .D(n_364), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_332), .Y(n_326) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g384 ( .A(n_329), .Y(n_384) );
INVx2_ASAP7_75t_SL g420 ( .A(n_329), .Y(n_420) );
INVx3_ASAP7_75t_L g496 ( .A(n_329), .Y(n_496) );
INVx2_ASAP7_75t_L g630 ( .A(n_329), .Y(n_630) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx3_ASAP7_75t_SL g468 ( .A(n_334), .Y(n_468) );
INVx2_ASAP7_75t_L g502 ( .A(n_334), .Y(n_502) );
INVx4_ASAP7_75t_L g555 ( .A(n_334), .Y(n_555) );
INVx2_ASAP7_75t_SL g623 ( .A(n_334), .Y(n_623) );
INVx8_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g385 ( .A(n_337), .Y(n_385) );
INVx2_ASAP7_75t_SL g418 ( .A(n_337), .Y(n_418) );
INVx2_ASAP7_75t_SL g497 ( .A(n_337), .Y(n_497) );
INVx2_ASAP7_75t_L g633 ( .A(n_337), .Y(n_633) );
INVx8_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g449 ( .A(n_342), .Y(n_449) );
BUFx3_ASAP7_75t_L g499 ( .A(n_342), .Y(n_499) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
OAI22xp33_ASAP7_75t_SL g635 ( .A1(n_344), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_635) );
INVx5_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g450 ( .A(n_345), .Y(n_450) );
BUFx2_ASAP7_75t_L g522 ( .A(n_345), .Y(n_522) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g390 ( .A(n_348), .Y(n_390) );
INVx3_ASAP7_75t_L g444 ( .A(n_348), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_348), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
INVx6_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g524 ( .A(n_349), .Y(n_524) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
BUFx2_ASAP7_75t_SL g552 ( .A(n_351), .Y(n_552) );
BUFx2_ASAP7_75t_SL g665 ( .A(n_351), .Y(n_665) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_358), .Y(n_352) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_355), .Y(n_401) );
INVx3_ASAP7_75t_L g462 ( .A(n_355), .Y(n_462) );
BUFx6f_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
BUFx4f_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
INVx2_ASAP7_75t_L g437 ( .A(n_357), .Y(n_437) );
BUFx3_ASAP7_75t_L g610 ( .A(n_357), .Y(n_610) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
BUFx2_ASAP7_75t_L g517 ( .A(n_360), .Y(n_517) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_360), .Y(n_613) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g399 ( .A(n_362), .Y(n_399) );
INVx2_ASAP7_75t_SL g412 ( .A(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
INVx2_ASAP7_75t_L g492 ( .A(n_362), .Y(n_492) );
INVx2_ASAP7_75t_L g518 ( .A(n_362), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_362), .A2(n_658), .B1(n_659), .B2(n_661), .Y(n_657) );
INVx6_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g538 ( .A(n_365), .Y(n_538) );
INVx4_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g431 ( .A(n_366), .Y(n_431) );
INVx4_ASAP7_75t_SL g457 ( .A(n_366), .Y(n_457) );
INVx3_ASAP7_75t_L g488 ( .A(n_366), .Y(n_488) );
INVx3_ASAP7_75t_SL g598 ( .A(n_366), .Y(n_598) );
INVx6_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g486 ( .A(n_369), .Y(n_486) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx5_ASAP7_75t_L g395 ( .A(n_370), .Y(n_395) );
BUFx3_ASAP7_75t_L g604 ( .A(n_370), .Y(n_604) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx3_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_424), .B2(n_476), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_378), .B1(n_404), .B2(n_405), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_393), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .C(n_388), .D(n_389), .Y(n_382) );
INVx1_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g445 ( .A(n_392), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .C(n_400), .D(n_403), .Y(n_393) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g602 ( .A(n_397), .Y(n_602) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .C(n_415), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .C(n_421), .D(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_451), .B1(n_473), .B2(n_475), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g428 ( .A(n_429), .B(n_438), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_430), .B(n_432), .C(n_434), .D(n_435), .Y(n_429) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g656 ( .A(n_437), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .C(n_443), .D(n_446), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g475 ( .A(n_451), .Y(n_475) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
XOR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_472), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_464), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .Y(n_459) );
INVx4_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g608 ( .A(n_462), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g580 ( .A(n_477), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_528), .B2(n_578), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OA22x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_505), .B2(n_506), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_504), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
XNOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_519), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
AOI22xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_556), .B1(n_574), .B2(n_575), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g577 ( .A(n_533), .Y(n_577) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_544), .Y(n_535) );
NOR2xp67_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_539), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g637 ( .A(n_548), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_557), .Y(n_574) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_566), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_583), .B(n_586), .Y(n_672) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OAI222xp33_ASAP7_75t_R g590 ( .A1(n_591), .A2(n_640), .B1(n_642), .B2(n_670), .C1(n_673), .C2(n_677), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND3x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_614), .C(n_626), .Y(n_593) );
NOR2xp67_ASAP7_75t_SL g594 ( .A(n_595), .B(n_605), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_599), .B(n_600), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g647 ( .A(n_598), .Y(n_647) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx6f_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g650 ( .A(n_604), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g654 ( .A(n_607), .Y(n_654) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx6f_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx4f_ASAP7_75t_SL g660 ( .A(n_613), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_624), .B2(n_625), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_635), .Y(n_626) );
OAI22xp33_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_631), .B1(n_632), .B2(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_662), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_652), .C(n_657), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_649), .B2(n_650), .C(n_651), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
CKINVDCx6p67_ASAP7_75t_R g671 ( .A(n_672), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_675), .Y(n_674) );
endmodule