module real_jpeg_17396_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_401),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_0),
.B(n_402),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.A3(n_28),
.B1(n_31),
.B2(n_37),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_1),
.A2(n_184),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_92),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_92),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_3),
.A2(n_92),
.B1(n_238),
.B2(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_5),
.A2(n_133),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_5),
.Y(n_281)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_6),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_7),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_7),
.A2(n_285),
.B1(n_304),
.B2(n_307),
.Y(n_303)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_9),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_10),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_10),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_10),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_13),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_374),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AO221x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_270),
.B1(n_272),
.B2(n_367),
.C(n_373),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_217),
.B(n_269),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_193),
.B(n_216),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_141),
.B(n_192),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_127),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_22),
.B(n_127),
.Y(n_192)
);

XOR2x2_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_64),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_23),
.B(n_96),
.C(n_125),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_24),
.B(n_43),
.Y(n_196)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_32),
.A2(n_281),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_34),
.Y(n_308)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_36),
.B(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_44),
.A2(n_131),
.B1(n_132),
.B2(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_45),
.B(n_53),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_98),
.B(n_101),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_48),
.A2(n_110),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_48),
.Y(n_173)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_48),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_52),
.B(n_282),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_56),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_60),
.A2(n_132),
.B(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_63),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_96),
.B1(n_125),
.B2(n_126),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_65),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_65),
.A2(n_125),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_65),
.B(n_275),
.C(n_276),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_65),
.A2(n_125),
.B1(n_275),
.B2(n_325),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_75),
.B1(n_81),
.B2(n_88),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_66),
.A2(n_75),
.B1(n_81),
.B2(n_88),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_66),
.A2(n_75),
.B(n_81),
.Y(n_338)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_66),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_74),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_74),
.Y(n_263)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_81),
.Y(n_389)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_95),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_96),
.A2(n_126),
.B1(n_144),
.B2(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_96),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_96),
.A2(n_126),
.B1(n_331),
.B2(n_359),
.Y(n_358)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_104),
.B1(n_114),
.B2(n_119),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_104),
.B1(n_114),
.B2(n_119),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_97),
.B(n_295),
.Y(n_313)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_145),
.A3(n_149),
.B1(n_151),
.B2(n_156),
.Y(n_144)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_104),
.Y(n_295)
);

NOR2x1p5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_108),
.Y(n_302)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_114),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_114),
.A2(n_295),
.B1(n_296),
.B2(n_303),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_116),
.Y(n_288)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_125),
.B(n_223),
.C(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.C(n_139),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_129),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_196),
.C(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_128),
.A2(n_129),
.B1(n_277),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_129),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_182),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_130),
.A2(n_163),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_131),
.A2(n_278),
.B1(n_282),
.B2(n_289),
.Y(n_277)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_140),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_388)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_166),
.B(n_191),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_162),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_163),
.B(n_254),
.Y(n_349)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_186),
.B(n_190),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_181),
.B(n_185),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_187),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_200),
.C(n_204),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_180),
.A2(n_278),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_184),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_215),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_215),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_214),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_213),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_200),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_200),
.A2(n_294),
.B(n_309),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_200),
.B(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_200),
.B(n_275),
.C(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_200),
.A2(n_213),
.B1(n_275),
.B2(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_229),
.B1(n_236),
.B2(n_246),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_237),
.B(n_242),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_229),
.B1(n_236),
.B2(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_206),
.B(n_236),
.Y(n_320)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_207),
.Y(n_394)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_207),
.Y(n_397)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_219),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_250),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_220),
.B(n_251),
.C(n_252),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_224),
.B(n_225),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_225),
.A2(n_297),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_227),
.A2(n_228),
.B1(n_337),
.B2(n_338),
.Y(n_344)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_228),
.Y(n_362)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_350),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_339),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_322),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_273),
.B(n_322),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_292),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_274),
.B(n_293),
.C(n_310),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_275),
.Y(n_325)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_310),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_298),
.A2(n_299),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_303),
.B(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_309),
.A2(n_381),
.B1(n_382),
.B2(n_398),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_311),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_315),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_321),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.C(n_329),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.C(n_337),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_342),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.C(n_348),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_346),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_349),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_363),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_353),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_358),
.C(n_360),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_362),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_370),
.Y(n_369)
);

NAND2x1_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_366),
.Y(n_368)
);

A2O1A1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B(n_371),
.C(n_372),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_399),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_377),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);


endmodule