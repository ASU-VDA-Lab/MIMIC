module real_jpeg_30343_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_0),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_0),
.Y(n_251)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_1),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_1),
.Y(n_78)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_78),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_1),
.B(n_106),
.Y(n_245)
);

OAI22x1_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_78),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_1),
.A2(n_272),
.A3(n_278),
.B1(n_282),
.B2(n_289),
.Y(n_271)
);

NAND2xp67_ASAP7_75t_SL g373 ( 
.A(n_1),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_1),
.B(n_161),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_4),
.B1(n_15),
.B2(n_18),
.Y(n_14)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_5),
.Y(n_257)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_5),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_6),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_7),
.A2(n_27),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_8),
.A2(n_44),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_8),
.A2(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_8),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_12),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_153),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_153),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_12),
.A2(n_153),
.B1(n_254),
.B2(n_258),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_13),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_234),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_232),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_209),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_21),
.B(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_116),
.C(n_172),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2x1_ASAP7_75t_L g421 ( 
.A(n_23),
.B(n_116),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_79),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_24),
.A2(n_80),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_25),
.Y(n_80)
);

XOR2x2_ASAP7_75t_L g430 ( 
.A(n_25),
.B(n_42),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_26),
.Y(n_208)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_31),
.Y(n_201)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_31),
.Y(n_204)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_31),
.Y(n_260)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_35),
.B(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_36),
.A2(n_198),
.B1(n_205),
.B2(n_208),
.Y(n_197)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_37),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_37),
.A2(n_253),
.B1(n_262),
.B2(n_319),
.Y(n_318)
);

NOR2x1_ASAP7_75t_R g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_53),
.B1(n_61),
.B2(n_73),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_43),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_52),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_64),
.B(n_69),
.Y(n_63)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_54),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_54),
.A2(n_63),
.B1(n_73),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_54),
.B(n_63),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_55),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_56),
.Y(n_376)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22x1_ASAP7_75t_L g335 ( 
.A1(n_62),
.A2(n_161),
.B1(n_327),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g364 ( 
.A1(n_64),
.A2(n_78),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_131),
.B1(n_134),
.B2(n_136),
.Y(n_130)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_65),
.Y(n_361)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_R g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_73),
.Y(n_327)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_85),
.B(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_78),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_78),
.B(n_130),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_78),
.B(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_113),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_81),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_83),
.A2(n_94),
.B1(n_112),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_83),
.A2(n_94),
.B1(n_112),
.B2(n_180),
.Y(n_429)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_84),
.B(n_95),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_88),
.A2(n_301),
.A3(n_304),
.B1(n_307),
.B2(n_310),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_88),
.A2(n_301),
.A3(n_304),
.B1(n_307),
.B2(n_310),
.Y(n_322)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_112),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_98),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_98),
.Y(n_313)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_107),
.Y(n_316)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_110),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_112),
.A2(n_180),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_171),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_157),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_118),
.A2(n_242),
.B1(n_243),
.B2(n_268),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_118),
.B(n_244),
.C(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_118),
.B(n_178),
.Y(n_407)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_158),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_128),
.B1(n_139),
.B2(n_149),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_120),
.A2(n_139),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_129),
.B1(n_140),
.B2(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_121),
.B(n_140),
.Y(n_226)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_128),
.A2(n_219),
.B(n_226),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_130),
.Y(n_403)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_146),
.Y(n_306)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_162),
.B(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx4f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_170),
.Y(n_293)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_172),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_173),
.B(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_187),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_174),
.A2(n_175),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_174),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_174),
.A2(n_175),
.B1(n_334),
.B2(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_174),
.B(n_228),
.C(n_326),
.Y(n_409)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g427 ( 
.A1(n_175),
.A2(n_176),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_177),
.B(n_268),
.C(n_394),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_186),
.Y(n_309)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g426 ( 
.A(n_188),
.B(n_427),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_240),
.C(n_269),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_189),
.A2(n_269),
.B1(n_270),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_189),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_189),
.B(n_317),
.C(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_189),
.A2(n_190),
.B1(n_350),
.B2(n_385),
.Y(n_384)
);

AO22x1_ASAP7_75t_L g396 ( 
.A1(n_189),
.A2(n_197),
.B1(n_340),
.B2(n_397),
.Y(n_396)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_191),
.Y(n_336)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_197),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_198),
.A2(n_205),
.B(n_261),
.Y(n_400)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx4f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_231),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_227),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_217),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_227),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_229),
.B(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_416),
.B(n_446),
.Y(n_235)
);

AOI211x1_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_341),
.B(n_389),
.C(n_415),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_329),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_295),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_239),
.B(n_295),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_241),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_267),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_246),
.B(n_372),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_252),
.B(n_261),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_251),
.Y(n_374)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_257),
.Y(n_369)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_267),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_267),
.B(n_355),
.Y(n_380)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_294),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_271),
.B(n_294),
.Y(n_337)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_323),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_297),
.B(n_323),
.C(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_298),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_317),
.B1(n_318),
.B2(n_322),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_300),
.B(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_R g377 ( 
.A(n_318),
.B(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_378),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_324),
.B(n_433),
.C(n_434),
.Y(n_432)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_338),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_338),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_337),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_334),
.A2(n_348),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_357),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_400),
.Y(n_399)
);

XOR2x2_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_400),
.Y(n_408)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_351),
.B(n_387),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_381),
.B(n_386),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_370),
.B(n_380),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_362),
.B(n_364),
.Y(n_357)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AOI21x1_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_377),
.B(n_379),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_382),
.B(n_383),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_410),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_418),
.Y(n_417)
);

NAND2x1_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_404),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_392),
.B(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_407),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_440),
.C(n_442),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_404),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.C(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_414),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_409),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_413),
.Y(n_418)
);

NAND4xp25_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.C(n_435),
.D(n_438),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_422),
.B(n_424),
.Y(n_419)
);

AND3x1_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_422),
.C(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_421),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.C(n_431),
.Y(n_424)
);

OAI22x1_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_426),
.B1(n_430),
.B2(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_443),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);


endmodule