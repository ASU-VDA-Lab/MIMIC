module real_jpeg_26374_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_352, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_352;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_89),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_30),
.C(n_44),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_1),
.B(n_72),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_1),
.A2(n_27),
.B1(n_169),
.B2(n_173),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_2),
.A2(n_49),
.B1(n_63),
.B2(n_66),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_2),
.A2(n_49),
.B1(n_78),
.B2(n_88),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_3),
.A2(n_38),
.B1(n_63),
.B2(n_66),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_3),
.A2(n_38),
.B1(n_81),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_59),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_59),
.B1(n_87),
.B2(n_88),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_63),
.B1(n_66),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_74),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_74),
.B1(n_78),
.B2(n_88),
.Y(n_233)
);

INVx8_ASAP7_75t_SL g85 ( 
.A(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_78),
.B1(n_88),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_9),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_9),
.A2(n_63),
.B1(n_66),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_92),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_10),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_10),
.A2(n_35),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_65),
.B1(n_78),
.B2(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_162)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_344),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_331),
.B(n_343),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_294),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_352),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_267),
.B(n_293),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_239),
.B(n_266),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_131),
.B(n_218),
.C(n_238),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_115),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_23),
.B(n_115),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_93),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_56),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_25),
.B(n_56),
.C(n_93),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_26),
.B(n_41),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_27),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_27),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_27),
.A2(n_36),
.B(n_151),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_27),
.A2(n_151),
.B(n_173),
.Y(n_245)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_28),
.A2(n_34),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_28),
.B(n_37),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_123),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_30),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_40),
.B(n_79),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_50),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_55),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_42),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_42),
.A2(n_52),
.B1(n_144),
.B2(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_42),
.B(n_79),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_42),
.A2(n_52),
.B(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_47),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_46),
.A2(n_70),
.B(n_184),
.C(n_186),
.Y(n_183)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_47),
.B(n_139),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g186 ( 
.A(n_47),
.B(n_66),
.C(n_69),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_50),
.B(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_58),
.B(n_60),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_51),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_51),
.A2(n_142),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_51),
.A2(n_142),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_52),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_52),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_75),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_58),
.B(n_142),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_61)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_66),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_80),
.B(n_84),
.C(n_113),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_63),
.B(n_79),
.CON(n_185),
.SN(n_185)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_77),
.C(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_67),
.A2(n_72),
.B1(n_129),
.B2(n_185),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_67),
.A2(n_104),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_67),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_67),
.A2(n_72),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_67),
.A2(n_235),
.B(n_274),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_67),
.A2(n_72),
.B(n_104),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_71),
.A2(n_102),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_71),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_71),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B(n_80),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_77),
.Y(n_286)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_78),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_82),
.A2(n_89),
.B1(n_99),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_82),
.B(n_285),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_82),
.A2(n_89),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_82),
.A2(n_319),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_83),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_89),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_89),
.B(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_105),
.B2(n_114),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_96),
.B(n_100),
.C(n_114),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_97),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_97),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_103),
.B(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_118),
.B(n_120),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_127),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_124),
.B(n_148),
.Y(n_224)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_127),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_217),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_212),
.B(n_216),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_196),
.B(n_211),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_179),
.B(n_195),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_158),
.B(n_178),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_140),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_153),
.C(n_156),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_165),
.B(n_177),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_164),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_171),
.B(n_176),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_190),
.C(n_191),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_206),
.C(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_229),
.C(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_265),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_250),
.B1(n_263),
.B2(n_264),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_264),
.C(n_265),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_245),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_244),
.A2(n_278),
.B(n_282),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_257),
.C(n_262),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_255),
.B(n_300),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_277),
.B1(n_288),
.B2(n_289),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_275),
.B(n_276),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_276),
.A2(n_296),
.B1(n_308),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_288),
.C(n_292),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_287),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_284),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_290),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_310),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_310),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_308),
.C(n_309),
.Y(n_295)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_298),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_303),
.C(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_313),
.C(n_323),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_304),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_315),
.C(n_317),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_323),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_333),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_341),
.B2(n_342),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_337),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_339),
.C(n_341),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_346),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_350),
.Y(n_349)
);


endmodule