module fake_jpeg_21603_n_328 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_52),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_33),
.Y(n_85)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_70),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_30),
.B1(n_39),
.B2(n_28),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_69),
.A2(n_93),
.B1(n_55),
.B2(n_28),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_74),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_25),
.B(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_77),
.B(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_30),
.B1(n_39),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_86),
.B1(n_89),
.B2(n_74),
.Y(n_122)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_82),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_36),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_36),
.B(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_42),
.B1(n_41),
.B2(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_42),
.B1(n_54),
.B2(n_53),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_60),
.B1(n_80),
.B2(n_67),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_24),
.B1(n_33),
.B2(n_37),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_112),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_53),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_108),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_49),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_49),
.B1(n_37),
.B2(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_127),
.B1(n_129),
.B2(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_117),
.Y(n_140)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_32),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_133),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_20),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_131),
.B(n_32),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_128),
.B1(n_4),
.B2(n_6),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_64),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_37),
.B1(n_28),
.B2(n_29),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_20),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_58),
.B(n_20),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_145),
.B1(n_159),
.B2(n_161),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_107),
.B(n_127),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_136),
.A2(n_137),
.B(n_141),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_107),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_60),
.B1(n_37),
.B2(n_73),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_2),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_104),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_3),
.B(n_37),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_111),
.B(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.Y(n_167)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_91),
.C(n_76),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_32),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_95),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_96),
.A2(n_27),
.B1(n_19),
.B2(n_7),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_27),
.B1(n_19),
.B2(n_7),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_109),
.B1(n_106),
.B2(n_111),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_27),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_109),
.B1(n_130),
.B2(n_115),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_105),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_187),
.Y(n_203)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_175),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_154),
.B1(n_160),
.B2(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_131),
.B1(n_121),
.B2(n_118),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_181),
.B1(n_164),
.B2(n_142),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_131),
.B1(n_121),
.B2(n_97),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_183),
.B(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_188),
.B1(n_191),
.B2(n_15),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_132),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_136),
.A2(n_115),
.B1(n_99),
.B2(n_120),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_8),
.B(n_9),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_116),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_140),
.A2(n_106),
.B1(n_9),
.B2(n_11),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_8),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_12),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_137),
.B(n_12),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_13),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_14),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_13),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_150),
.B1(n_162),
.B2(n_156),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_209),
.B1(n_213),
.B2(n_215),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_160),
.B1(n_158),
.B2(n_154),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_166),
.B1(n_141),
.B2(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_157),
.C(n_140),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_218),
.C(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_171),
.A2(n_148),
.B1(n_151),
.B2(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_143),
.C(n_15),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_191),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_16),
.B1(n_17),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_16),
.B1(n_17),
.B2(n_181),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_173),
.A2(n_17),
.B1(n_172),
.B2(n_193),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_229),
.B(n_233),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_168),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_199),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_242),
.C(n_218),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_225),
.B1(n_223),
.B2(n_212),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_210),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_168),
.C(n_174),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_208),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_185),
.B(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_177),
.B1(n_198),
.B2(n_188),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_221),
.B1(n_207),
.B2(n_183),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_260),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_262),
.B1(n_269),
.B2(n_271),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_206),
.B1(n_205),
.B2(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_266),
.Y(n_281)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_231),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_205),
.B1(n_213),
.B2(n_182),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_274),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_241),
.B1(n_222),
.B2(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_240),
.C(n_242),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_238),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_255),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_241),
.B1(n_225),
.B2(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_230),
.C(n_237),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_283),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

AO22x1_ASAP7_75t_SL g286 ( 
.A1(n_259),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_254),
.B1(n_263),
.B2(n_260),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_296),
.Y(n_302)
);

FAx1_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_267),
.CI(n_264),
.CON(n_290),
.SN(n_290)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_277),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_297),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_265),
.B(n_257),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_280),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_275),
.B(n_194),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_284),
.C(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_284),
.C(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_266),
.B1(n_243),
.B2(n_252),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_304),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_286),
.B(n_221),
.C(n_229),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_294),
.B1(n_295),
.B2(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_217),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_252),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_289),
.CI(n_296),
.CON(n_309),
.SN(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_300),
.B1(n_305),
.B2(n_291),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_305),
.C(n_207),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_286),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_312),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_308),
.B1(n_311),
.B2(n_310),
.Y(n_323)
);

OAI311xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_318),
.A3(n_322),
.B1(n_321),
.C1(n_309),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_309),
.B(n_246),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);

OAI221xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_246),
.B1(n_247),
.B2(n_195),
.C(n_219),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_247),
.Y(n_328)
);


endmodule