module real_jpeg_9568_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_17;
wire n_21;
wire n_29;
wire n_31;
wire n_24;
wire n_28;
wire n_23;
wire n_25;
wire n_22;
wire n_18;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_19),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_0),
.A2(n_29),
.B(n_32),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_14),
.C(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_SL g30 ( 
.A(n_4),
.B(n_6),
.C(n_15),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_SL g16 ( 
.A1(n_5),
.A2(n_17),
.A3(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_9),
.C(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND4xp25_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.D(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);


endmodule