module fake_jpeg_866_n_556 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_556);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_556;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_53),
.B(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_57),
.B(n_64),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_61),
.Y(n_162)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_18),
.C(n_1),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_32),
.B(n_48),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_18),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_88),
.B(n_1),
.Y(n_158)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_0),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_40),
.C(n_41),
.Y(n_120)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_24),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_103),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_120),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_106),
.B(n_121),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_26),
.B1(n_35),
.B2(n_46),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_109),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_51),
.B1(n_46),
.B2(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_111),
.A2(n_125),
.B1(n_135),
.B2(n_144),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_39),
.B(n_25),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_45),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_55),
.A2(n_34),
.B1(n_51),
.B2(n_46),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_134),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_34),
.B1(n_51),
.B2(n_46),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_147),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_34),
.B1(n_51),
.B2(n_38),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_26),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_26),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_35),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_158),
.B(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_79),
.B(n_35),
.Y(n_161)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_33),
.A3(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_170),
.B(n_179),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_38),
.B1(n_39),
.B2(n_33),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_171),
.B(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_173),
.B(n_176),
.Y(n_230)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_177),
.A2(n_192),
.B1(n_196),
.B2(n_201),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_178),
.B(n_187),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_104),
.C(n_101),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_184),
.A2(n_222),
.B(n_228),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_23),
.B1(n_25),
.B2(n_92),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_191),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_52),
.B1(n_74),
.B2(n_84),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_120),
.A2(n_111),
.B1(n_135),
.B2(n_144),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_97),
.C(n_90),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_221),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_83),
.B1(n_56),
.B2(n_78),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_59),
.B1(n_73),
.B2(n_69),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_215),
.B1(n_226),
.B2(n_146),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_23),
.B1(n_25),
.B2(n_80),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_122),
.A2(n_65),
.B1(n_50),
.B2(n_31),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

BUFx4f_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_118),
.A2(n_31),
.B1(n_19),
.B2(n_49),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_140),
.A2(n_31),
.B1(n_19),
.B2(n_47),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_217),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_123),
.B(n_19),
.Y(n_222)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_133),
.A2(n_138),
.B1(n_137),
.B2(n_143),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_133),
.A2(n_31),
.B1(n_19),
.B2(n_4),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_227),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

AND2x4_ASAP7_75t_SL g228 ( 
.A(n_132),
.B(n_19),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_231),
.A2(n_6),
.B(n_7),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_151),
.B1(n_137),
.B2(n_146),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_233),
.A2(n_280),
.B1(n_208),
.B2(n_194),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_236),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_130),
.B(n_122),
.C(n_166),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_246),
.A2(n_263),
.B(n_262),
.C(n_257),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_117),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_274),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_266),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_205),
.A2(n_130),
.B1(n_154),
.B2(n_138),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_277),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_222),
.A2(n_123),
.B(n_127),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_262),
.A2(n_6),
.B(n_7),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_129),
.B(n_31),
.C(n_19),
.Y(n_263)
);

NAND2x1_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_143),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_171),
.B(n_182),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_211),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_177),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_277),
.B1(n_227),
.B2(n_201),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_204),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_200),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_219),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_192),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_225),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_284),
.B(n_312),
.Y(n_363)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_175),
.B1(n_207),
.B2(n_210),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_286),
.A2(n_308),
.B1(n_313),
.B2(n_326),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_179),
.C(n_199),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_304),
.C(n_309),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_293),
.Y(n_362)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_231),
.A3(n_249),
.B1(n_242),
.B2(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_230),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_300),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_269),
.A2(n_170),
.B1(n_220),
.B2(n_213),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_297),
.A2(n_321),
.B1(n_281),
.B2(n_264),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_298),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_251),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_190),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_169),
.C(n_168),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_188),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_311),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_181),
.C(n_174),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_186),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_224),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_191),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_324),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_197),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_315),
.B(n_319),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_316),
.A2(n_317),
.B(n_281),
.Y(n_349)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_279),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_320),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_255),
.A2(n_218),
.B1(n_198),
.B2(n_189),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_221),
.C(n_214),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_257),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_216),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_257),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_325),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_268),
.A2(n_208),
.B1(n_216),
.B2(n_8),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_271),
.A2(n_259),
.B1(n_256),
.B2(n_243),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_327),
.A2(n_329),
.B1(n_278),
.B2(n_248),
.Y(n_359)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_250),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_259),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_246),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_365),
.C(n_373),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_337),
.A2(n_360),
.B1(n_370),
.B2(n_372),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_243),
.B(n_256),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_339),
.A2(n_346),
.B(n_347),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_358),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_263),
.B(n_260),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_291),
.A2(n_260),
.B(n_280),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_314),
.Y(n_383)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_295),
.B(n_248),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_359),
.A2(n_258),
.B1(n_10),
.B2(n_11),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_273),
.B1(n_253),
.B2(n_237),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_322),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_310),
.B1(n_313),
.B2(n_327),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_366),
.A2(n_369),
.B1(n_283),
.B2(n_285),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_278),
.B(n_267),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_330),
.B(n_282),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_310),
.A2(n_297),
.B1(n_303),
.B2(n_321),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_310),
.A2(n_273),
.B1(n_237),
.B2(n_267),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_309),
.A2(n_244),
.B1(n_241),
.B2(n_240),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_304),
.B(n_244),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_338),
.A2(n_296),
.B1(n_326),
.B2(n_293),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_391),
.B1(n_363),
.B2(n_361),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_376),
.B(n_380),
.Y(n_420)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_331),
.B(n_284),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_379),
.B(n_400),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_371),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_388),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_382),
.A2(n_383),
.B(n_384),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_288),
.B(n_290),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_385),
.A2(n_396),
.B1(n_399),
.B2(n_401),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_292),
.B(n_328),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_344),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_289),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_394),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_346),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_404),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_338),
.A2(n_324),
.B1(n_300),
.B2(n_329),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_336),
.B(n_299),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_318),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_402),
.C(n_390),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_302),
.B1(n_301),
.B2(n_294),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_294),
.B1(n_306),
.B2(n_307),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_241),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_337),
.A2(n_307),
.B1(n_240),
.B2(n_235),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_335),
.B(n_235),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_352),
.A2(n_347),
.B1(n_360),
.B2(n_349),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_403),
.A2(n_342),
.B1(n_359),
.B2(n_349),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_410),
.B1(n_370),
.B2(n_334),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_258),
.Y(n_407)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_9),
.B(n_11),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_408),
.Y(n_422)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_427),
.B1(n_382),
.B2(n_408),
.Y(n_449)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_373),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_418),
.C(n_439),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_345),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_423),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_421),
.B(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_342),
.Y(n_423)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_374),
.B(n_333),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_429),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_384),
.B(n_354),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_377),
.B(n_372),
.C(n_342),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_436),
.C(n_381),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_399),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_385),
.A2(n_388),
.B1(n_383),
.B2(n_398),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_435),
.A2(n_375),
.B1(n_391),
.B2(n_389),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_342),
.C(n_354),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_367),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_383),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_440),
.B(n_15),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_357),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_356),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_397),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_461),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_446),
.A2(n_459),
.B1(n_437),
.B2(n_422),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_375),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_460),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_392),
.B1(n_409),
.B2(n_405),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_448),
.A2(n_449),
.B1(n_450),
.B2(n_456),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_435),
.Y(n_451)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_461),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_407),
.C(n_357),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_458),
.C(n_466),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_410),
.B1(n_393),
.B2(n_378),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_348),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_343),
.C(n_350),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_343),
.B1(n_350),
.B2(n_406),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_356),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_12),
.Y(n_462)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_441),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_12),
.B(n_13),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_422),
.B(n_441),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_418),
.B(n_442),
.C(n_432),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_12),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_464),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_470),
.B(n_477),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_446),
.B1(n_450),
.B2(n_459),
.Y(n_497)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_473),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_444),
.B(n_423),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_476),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_454),
.B(n_439),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_467),
.Y(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_436),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_484),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_467),
.A2(n_416),
.B(n_433),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_480),
.A2(n_482),
.B(n_434),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_453),
.A2(n_433),
.B(n_438),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_454),
.B(n_443),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_413),
.C(n_424),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_490),
.C(n_492),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_413),
.C(n_424),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_492),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_466),
.B(n_431),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_457),
.Y(n_493)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_451),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_494),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_472),
.B(n_445),
.CI(n_455),
.CON(n_495),
.SN(n_495)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_503),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_497),
.A2(n_485),
.B1(n_486),
.B2(n_473),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_482),
.A2(n_469),
.B1(n_456),
.B2(n_465),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_502),
.A2(n_510),
.B1(n_477),
.B2(n_489),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_504),
.B(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_469),
.C(n_431),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_13),
.C(n_471),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_509),
.C(n_479),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_480),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_508),
.B(n_481),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_490),
.C(n_487),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_513),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_491),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_516),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_517),
.A2(n_523),
.B1(n_497),
.B2(n_495),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_504),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_521),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_484),
.C(n_475),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_499),
.C(n_498),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_505),
.Y(n_521)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_494),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_476),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_525),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_500),
.B(n_502),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_512),
.A2(n_496),
.B(n_493),
.C(n_501),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_526),
.B(n_533),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_520),
.A2(n_496),
.B(n_499),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_SL g539 ( 
.A(n_528),
.B(n_519),
.C(n_516),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_530),
.B(n_518),
.Y(n_538)
);

INVx11_ASAP7_75t_L g533 ( 
.A(n_522),
.Y(n_533)
);

OAI31xp67_ASAP7_75t_L g534 ( 
.A1(n_512),
.A2(n_510),
.A3(n_501),
.B(n_503),
.Y(n_534)
);

O2A1O1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_534),
.A2(n_514),
.B(n_495),
.C(n_517),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_535),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_537),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_538),
.B(n_541),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_539),
.A2(n_532),
.B1(n_534),
.B2(n_531),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_529),
.B(n_515),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_531),
.B(n_511),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_542),
.A2(n_536),
.B(n_527),
.Y(n_544)
);

AOI21xp33_ASAP7_75t_L g548 ( 
.A1(n_544),
.A2(n_543),
.B(n_540),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_526),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_548),
.A2(n_549),
.B(n_550),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_530),
.C(n_533),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_546),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_526),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_553),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_552),
.B(n_526),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_524),
.Y(n_556)
);


endmodule