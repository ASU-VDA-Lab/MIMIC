module fake_jpeg_11677_n_288 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_21),
.B1(n_36),
.B2(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_37),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_1),
.C(n_3),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_19),
.CON(n_56),
.SN(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_19),
.B1(n_37),
.B2(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_77),
.B1(n_20),
.B2(n_34),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_22),
.B1(n_44),
.B2(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_25),
.C(n_29),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_26),
.C(n_27),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_84),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_101),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_88),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_120),
.B1(n_68),
.B2(n_5),
.Y(n_134)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_28),
.A3(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_17),
.B(n_16),
.C(n_15),
.Y(n_131)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_113),
.C(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

OR2x4_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_4),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_117),
.B1(n_81),
.B2(n_62),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_57),
.B(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_67),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_66),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_83),
.B1(n_76),
.B2(n_74),
.Y(n_124)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_72),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_127),
.B1(n_109),
.B2(n_90),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_113),
.B(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_128),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_75),
.B1(n_80),
.B2(n_82),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_118),
.B(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_84),
.B1(n_75),
.B2(n_80),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_68),
.A3(n_62),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_12),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_68),
.C(n_7),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_102),
.C(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_10),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_103),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_162),
.C(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_158),
.B(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_116),
.B(n_110),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_175),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_97),
.B1(n_116),
.B2(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_126),
.B1(n_125),
.B2(n_163),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_104),
.B(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_91),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_86),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_107),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_143),
.B1(n_132),
.B2(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_90),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_94),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_104),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_11),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_12),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_13),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_189),
.B1(n_169),
.B2(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_137),
.B(n_141),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_183),
.B(n_156),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_137),
.B(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_171),
.C(n_158),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_125),
.B1(n_143),
.B2(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_125),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_150),
.B1(n_166),
.B2(n_165),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_132),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_154),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_146),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_155),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_13),
.B1(n_161),
.B2(n_163),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_168),
.B(n_178),
.C(n_164),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_220),
.B1(n_211),
.B2(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_212),
.B1(n_213),
.B2(n_225),
.Y(n_229)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_214),
.B1(n_216),
.B2(n_224),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_160),
.B(n_170),
.Y(n_211)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_226),
.B(n_184),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_179),
.B1(n_160),
.B2(n_169),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_179),
.B1(n_162),
.B2(n_151),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_162),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_217),
.C(n_201),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_195),
.B1(n_185),
.B2(n_181),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_152),
.B1(n_175),
.B2(n_172),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_205),
.B(n_183),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_198),
.B(n_188),
.C(n_192),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_237),
.B(n_238),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_235),
.B(n_242),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_184),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_210),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_197),
.C(n_199),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_206),
.B1(n_214),
.B2(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_247),
.B1(n_254),
.B2(n_255),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_236),
.B1(n_219),
.B2(n_233),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_243),
.B1(n_246),
.B2(n_249),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_213),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_222),
.B1(n_221),
.B2(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_228),
.C(n_197),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_265),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_237),
.B1(n_223),
.B2(n_241),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_245),
.B1(n_250),
.B2(n_252),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_192),
.B1(n_199),
.B2(n_203),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_207),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_258),
.B(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_267),
.B(n_269),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_266),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_203),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_256),
.C(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_265),
.C(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_200),
.B1(n_260),
.B2(n_196),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_268),
.C(n_196),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_269),
.B(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_273),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.Y(n_288)
);


endmodule