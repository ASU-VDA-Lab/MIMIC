module fake_jpeg_30711_n_365 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_67),
.B1(n_21),
.B2(n_24),
.Y(n_118)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_14),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_58),
.Y(n_96)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_11),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_64),
.C(n_76),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_15),
.B(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_17),
.A2(n_10),
.B1(n_9),
.B2(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_20),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_32),
.Y(n_111)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_22),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_37),
.B(n_16),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_SL g169 ( 
.A(n_83),
.B(n_100),
.C(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_84),
.B(n_105),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_101),
.B1(n_102),
.B2(n_118),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_2),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_95),
.B(n_111),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_36),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_26),
.B1(n_18),
.B2(n_23),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_47),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_36),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_18),
.B1(n_73),
.B2(n_57),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_35),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_60),
.A2(n_26),
.B1(n_77),
.B2(n_61),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_127),
.B1(n_45),
.B2(n_63),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_24),
.B1(n_80),
.B2(n_29),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_132),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_29),
.B(n_35),
.C(n_23),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_131),
.B(n_138),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_56),
.B(n_75),
.C(n_77),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_112),
.B(n_87),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_94),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_143),
.Y(n_176)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_151),
.B1(n_107),
.B2(n_92),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_142),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_55),
.B1(n_53),
.B2(n_49),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_94),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_165),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_149),
.Y(n_207)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_66),
.B1(n_61),
.B2(n_79),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_157),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_153),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_56),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_167),
.B1(n_135),
.B2(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_98),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_92),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_74),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_89),
.A2(n_2),
.B(n_5),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_7),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_5),
.B1(n_7),
.B2(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_172),
.Y(n_189)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_182),
.B(n_160),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_91),
.C(n_85),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_204),
.C(n_143),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_192),
.B1(n_173),
.B2(n_165),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_134),
.A2(n_103),
.B1(n_110),
.B2(n_93),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_130),
.B(n_97),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_97),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_132),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_110),
.B1(n_120),
.B2(n_122),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_211),
.B1(n_153),
.B2(n_156),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_120),
.C(n_81),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_149),
.A2(n_81),
.B(n_7),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_154),
.B(n_131),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_144),
.Y(n_206)
);

NAND2x1_ASAP7_75t_L g209 ( 
.A(n_133),
.B(n_135),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_150),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_138),
.B(n_170),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_143),
.B1(n_140),
.B2(n_139),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_228),
.B1(n_230),
.B2(n_192),
.Y(n_266)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_224),
.B(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_231),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_223),
.B(n_194),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_232),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_143),
.C(n_136),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_146),
.B1(n_137),
.B2(n_162),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_174),
.B(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_174),
.B(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_172),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_191),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_239),
.Y(n_249)
);

HAxp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_189),
.CON(n_236),
.SN(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_241),
.Y(n_255)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_188),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_177),
.B(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_188),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_183),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_176),
.C(n_207),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_261),
.C(n_208),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_220),
.B(n_229),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_184),
.B(n_182),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_176),
.Y(n_260)
);

AO22x1_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_209),
.B1(n_184),
.B2(n_205),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_264),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_221),
.B(n_185),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_230),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_223),
.B1(n_217),
.B2(n_228),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_194),
.B(n_183),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_225),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_294),
.B1(n_272),
.B2(n_249),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_262),
.B1(n_261),
.B2(n_268),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_260),
.B1(n_252),
.B2(n_256),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_277),
.Y(n_306)
);

AOI211xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_226),
.B(n_240),
.C(n_224),
.Y(n_280)
);

OAI321xp33_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_289),
.A3(n_250),
.B1(n_252),
.B2(n_267),
.C(n_251),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_214),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_283),
.C(n_247),
.Y(n_297)
);

OAI322xp33_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_234),
.A3(n_214),
.B1(n_233),
.B2(n_241),
.C1(n_213),
.C2(n_215),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_255),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_287),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_243),
.A3(n_186),
.B1(n_190),
.B2(n_232),
.C1(n_227),
.C2(n_198),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_200),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_208),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_200),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_262),
.A2(n_186),
.B1(n_237),
.B2(n_219),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_305),
.B1(n_312),
.B2(n_280),
.Y(n_320)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_297),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_271),
.B1(n_266),
.B2(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_257),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_285),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_275),
.A2(n_265),
.B1(n_250),
.B2(n_253),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_293),
.C(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_269),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_311),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_278),
.A2(n_265),
.B1(n_257),
.B2(n_251),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_316),
.B(n_321),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_320),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_278),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_246),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_273),
.B1(n_294),
.B2(n_286),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_286),
.B(n_258),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_325),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_298),
.A2(n_258),
.B(n_270),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_281),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_309),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_299),
.C(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.C(n_317),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_309),
.C(n_305),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_331),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_306),
.Y(n_331)
);

OAI211xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_297),
.B(n_307),
.C(n_311),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_239),
.B(n_187),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_312),
.B1(n_259),
.B2(n_276),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_254),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_270),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_347),
.C(n_329),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_336),
.A2(n_319),
.B(n_318),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_344),
.B(n_342),
.Y(n_349)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_337),
.B(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

AOI31xp67_ASAP7_75t_SL g343 ( 
.A1(n_332),
.A2(n_322),
.A3(n_316),
.B(n_259),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_343),
.A2(n_346),
.B1(n_203),
.B2(n_187),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_254),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_354),
.C(n_339),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_349),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g355 ( 
.A(n_350),
.B(n_351),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_337),
.B(n_254),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_181),
.B(n_203),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_347),
.A2(n_181),
.B1(n_203),
.B2(n_345),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_358),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_356),
.B(n_353),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_359),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_355),
.A2(n_350),
.B(n_203),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_360),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_361),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_363),
.Y(n_365)
);


endmodule