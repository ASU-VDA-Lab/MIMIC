module fake_jpeg_13519_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_72),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_1),
.C(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_57),
.Y(n_77)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_60),
.B1(n_59),
.B2(n_45),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_76),
.B1(n_48),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_59),
.B1(n_49),
.B2(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_54),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_85),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_61),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_62),
.B1(n_48),
.B2(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_63),
.C(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_51),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_55),
.B(n_57),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_67),
.B1(n_49),
.B2(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_24),
.B1(n_39),
.B2(n_11),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_30),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_7),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_40),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_29),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_99),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_121),
.B1(n_125),
.B2(n_115),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_35),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_124),
.C(n_103),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_37),
.C(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_127),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_100),
.CI(n_107),
.CON(n_131),
.SN(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_130),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_141),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_128),
.C(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_142),
.B(n_133),
.Y(n_144)
);

OAI31xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_131),
.A3(n_141),
.B(n_109),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_118),
.A3(n_127),
.B1(n_116),
.B2(n_121),
.C1(n_111),
.C2(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_136),
.C(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_134),
.C(n_115),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_148),
.Y(n_149)
);


endmodule