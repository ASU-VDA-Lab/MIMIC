module real_jpeg_4094_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_1),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_1),
.A2(n_198),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_1),
.A2(n_30),
.B1(n_174),
.B2(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_96),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_96),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_85),
.B1(n_96),
.B2(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_6),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_12),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_7),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_89),
.B1(n_126),
.B2(n_131),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_49),
.B1(n_89),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_89),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_12),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_12),
.A2(n_56),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_12),
.A2(n_56),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_12),
.A2(n_56),
.B1(n_185),
.B2(n_230),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_12),
.A2(n_140),
.B(n_266),
.C(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_12),
.B(n_61),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_12),
.B(n_300),
.C(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_12),
.B(n_124),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_12),
.B(n_119),
.C(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_12),
.B(n_32),
.Y(n_337)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_413),
.B(n_417),
.Y(n_19)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_147),
.B(n_412),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_144),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_22),
.B(n_144),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_133),
.C(n_142),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_23),
.B(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_58),
.C(n_91),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_24),
.A2(n_195),
.B1(n_206),
.B2(n_207),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_24),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_24),
.B(n_154),
.C(n_207),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_24),
.B(n_245),
.C(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_24),
.A2(n_206),
.B1(n_245),
.B2(n_338),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_24),
.A2(n_206),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_54),
.B2(n_57),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_25),
.A2(n_31),
.B1(n_54),
.B2(n_57),
.Y(n_232)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_28),
.Y(n_138)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_29),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_31),
.B(n_54),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_31),
.A2(n_57),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_31),
.A2(n_54),
.B(n_57),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_31),
.B(n_57),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_44),
.Y(n_31)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_34),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_35),
.Y(n_266)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_40),
.Y(n_132)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_56),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_57),
.A2(n_134),
.B(n_141),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_58),
.A2(n_91),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_58),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_58),
.B(n_232),
.C(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_58),
.A2(n_387),
.B1(n_389),
.B2(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_87),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_60),
.A2(n_73),
.B1(n_158),
.B2(n_163),
.Y(n_157)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_60),
.A2(n_73),
.B1(n_158),
.B2(n_163),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_60),
.A2(n_73),
.B(n_163),
.Y(n_349)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_71),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_73),
.B(n_163),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_80),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_87),
.A2(n_211),
.B1(n_213),
.B2(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_90),
.Y(n_212)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_91),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_99),
.B1(n_124),
.B2(n_125),
.Y(n_91)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_92),
.Y(n_390)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_98),
.Y(n_270)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_99),
.A2(n_124),
.B1(n_196),
.B2(n_201),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_99),
.B(n_196),
.Y(n_391)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_101),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_100),
.A2(n_101),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_101),
.A2(n_390),
.B(n_391),
.Y(n_389)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_109),
.B2(n_112),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_118),
.Y(n_320)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_133),
.B(n_142),
.Y(n_409)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_143),
.B(n_196),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_144),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_144),
.B(n_414),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_145),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_407),
.B(n_411),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_378),
.B(n_404),
.Y(n_148)
);

OAI211xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_277),
.B(n_373),
.C(n_377),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_252),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_151),
.A2(n_252),
.B(n_374),
.C(n_376),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_233),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_152),
.B(n_233),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_208),
.C(n_220),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_153),
.B(n_208),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_194),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_169),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_155),
.A2(n_169),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_155),
.A2(n_262),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_156),
.A2(n_157),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_176),
.B1(n_183),
.B2(n_190),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_170),
.A2(n_225),
.B(n_228),
.Y(n_224)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_173),
.Y(n_303)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_176),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_177),
.A2(n_229),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_177),
.A2(n_229),
.B1(n_273),
.B2(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_182),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_195),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_195),
.A2(n_207),
.B1(n_222),
.B2(n_223),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_195),
.B(n_222),
.C(n_317),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_195),
.A2(n_207),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_195),
.B(n_258),
.C(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

INVx6_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_219),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_215),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.B(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_219),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_215),
.A2(n_239),
.B(n_240),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_216),
.B(n_229),
.Y(n_323)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.C(n_232),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_222),
.A2(n_223),
.B1(n_296),
.B2(n_304),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_304),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_224),
.Y(n_365)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_232),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_232),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_232),
.A2(n_258),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_232),
.A2(n_258),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_232),
.A2(n_258),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_232),
.B(n_383),
.C(n_388),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_250),
.B2(n_251),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_241),
.B1(n_242),
.B2(n_249),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_241),
.B(n_249),
.C(n_251),
.Y(n_403)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_245),
.B(n_248),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_245),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_248),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_248),
.A2(n_393),
.B1(n_397),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_253),
.B(n_255),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.C(n_263),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_256),
.B(n_260),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_272),
.C(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_330),
.C(n_332),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_263),
.B(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_264),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_265),
.A2(n_271),
.B1(n_272),
.B2(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_265),
.Y(n_355)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_272),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_291),
.Y(n_292)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_357),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_342),
.B(n_356),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_327),
.B(n_341),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_314),
.B(n_326),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_306),
.B(n_313),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_293),
.B(n_305),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_290),
.B(n_292),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_294),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_336),
.C(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_324),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_340),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_332),
.B1(n_333),
.B2(n_339),
.Y(n_328)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_344),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_352),
.C(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_360),
.B(n_368),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_360),
.C(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_366),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_364),
.A2(n_366),
.B1(n_367),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_370),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_399),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_392),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_392),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.C(n_398),
.Y(n_392)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_403),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_410),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_418),
.Y(n_417)
);


endmodule