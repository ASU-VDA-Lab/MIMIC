module fake_jpeg_29862_n_57 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_17),
.A3(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_23),
.C(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_5),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_22),
.B(n_4),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_36),
.C(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_39),
.C(n_7),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_8),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_45),
.B(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_53),
.B(n_51),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_47),
.C(n_48),
.Y(n_57)
);


endmodule