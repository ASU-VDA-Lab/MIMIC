module fake_aes_7053_n_10 (n_1, n_0, n_10);
input n_1;
input n_0;
output n_10;
wire n_2;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
BUFx2_ASAP7_75t_L g2 ( .A(n_1), .Y(n_2) );
NAND2xp5_ASAP7_75t_L g3 ( .A(n_2), .B(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_3), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_6), .B(n_5), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_7), .Y(n_8) );
INVx2_ASAP7_75t_SL g9 ( .A(n_8), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
endmodule