module fake_jpeg_27916_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_33),
.B1(n_28),
.B2(n_24),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_86)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_40),
.B1(n_28),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_75),
.B1(n_81),
.B2(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_84),
.Y(n_108)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_74),
.B1(n_89),
.B2(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_41),
.B1(n_25),
.B2(n_19),
.Y(n_75)
);

AND2x4_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_43),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_39),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_30),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_41),
.B1(n_25),
.B2(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_25),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_92),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_88),
.B1(n_96),
.B2(n_39),
.Y(n_112)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_23),
.B1(n_21),
.B2(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_56),
.B1(n_60),
.B2(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_14),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_43),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_16),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_23),
.B1(n_21),
.B2(n_17),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_115),
.B1(n_107),
.B2(n_102),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_55),
.B1(n_58),
.B2(n_54),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_105),
.B1(n_125),
.B2(n_75),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_45),
.B1(n_17),
.B2(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_76),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_37),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_90),
.B(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_65),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_72),
.B1(n_91),
.B2(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_129),
.A2(n_1),
.B(n_3),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_94),
.B1(n_68),
.B2(n_85),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_87),
.B1(n_63),
.B2(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_63),
.B1(n_93),
.B2(n_73),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_135),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_121),
.B1(n_125),
.B2(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_156),
.B1(n_157),
.B2(n_115),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_104),
.B(n_107),
.C(n_18),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_80),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_71),
.C(n_77),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_106),
.C(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_113),
.B1(n_111),
.B2(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_151),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_90),
.B1(n_66),
.B2(n_20),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_66),
.B1(n_77),
.B2(n_13),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_107),
.B1(n_102),
.B2(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_15),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_15),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_20),
.B1(n_77),
.B2(n_26),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_16),
.B1(n_26),
.B2(n_18),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_16),
.B1(n_26),
.B2(n_18),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_120),
.C(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_173),
.C(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_168),
.B1(n_171),
.B2(n_184),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_102),
.B1(n_124),
.B2(n_103),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_27),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_123),
.C(n_27),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_123),
.C(n_27),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_123),
.C(n_27),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_186),
.C(n_157),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_1),
.B(n_3),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_183),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_191),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_14),
.C(n_13),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_133),
.B1(n_144),
.B2(n_136),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_147),
.B1(n_141),
.B2(n_7),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_190),
.B1(n_155),
.B2(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_142),
.B1(n_138),
.B2(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_216),
.B1(n_189),
.B2(n_168),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_154),
.C(n_137),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_203),
.B(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_206),
.A2(n_207),
.B(n_211),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_140),
.B(n_156),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_158),
.A2(n_141),
.B1(n_6),
.B2(n_7),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_165),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_5),
.C(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_188),
.C(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_219),
.A2(n_201),
.B1(n_199),
.B2(n_212),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_226),
.B1(n_240),
.B2(n_243),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_210),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_224),
.B1(n_231),
.B2(n_228),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_166),
.B1(n_179),
.B2(n_165),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_173),
.C(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_165),
.C(n_167),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_165),
.C(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_5),
.C(n_7),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_236),
.C(n_218),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_8),
.C(n_9),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_192),
.A2(n_8),
.B(n_9),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_202),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_205),
.B1(n_192),
.B2(n_197),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_250),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_214),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_248),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_197),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_196),
.B1(n_215),
.B2(n_204),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_254),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_209),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_216),
.B1(n_196),
.B2(n_194),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_206),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_262),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_223),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_217),
.B1(n_198),
.B2(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_227),
.C(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_275),
.C(n_253),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_227),
.B1(n_225),
.B2(n_195),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_279),
.B1(n_200),
.B2(n_237),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_220),
.C(n_236),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_220),
.B1(n_249),
.B2(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_235),
.C(n_222),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_243),
.B1(n_195),
.B2(n_207),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_247),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_287),
.Y(n_301)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_258),
.B(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2x1_ASAP7_75t_R g286 ( 
.A(n_271),
.B(n_251),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_265),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_254),
.C(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_268),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_10),
.C(n_11),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_11),
.C(n_12),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_277),
.B(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_291),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_266),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_283),
.C(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_309),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_268),
.C(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_285),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_286),
.B(n_11),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_298),
.B(n_300),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_299),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_302),
.B1(n_308),
.B2(n_303),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_296),
.Y(n_323)
);


endmodule