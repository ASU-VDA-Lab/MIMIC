module fake_jpeg_30483_n_256 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_17),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_53),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_21),
.B(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_59),
.Y(n_84)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_0),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_76),
.B1(n_40),
.B2(n_33),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_41),
.B(n_11),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_97),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_46),
.B1(n_61),
.B2(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_26),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_19),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_111),
.B1(n_116),
.B2(n_120),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_64),
.B(n_25),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_47),
.B1(n_58),
.B2(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_119),
.B1(n_66),
.B2(n_67),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_123),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_45),
.B1(n_33),
.B2(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_50),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_78),
.B(n_88),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_124),
.B1(n_76),
.B2(n_98),
.Y(n_139)
);

NAND2x1_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_30),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_67),
.B(n_87),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_68),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_2),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_8),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_150),
.B1(n_153),
.B2(n_115),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_156),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_78),
.B(n_73),
.C(n_72),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_140),
.B(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_9),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_122),
.B(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_95),
.B1(n_73),
.B2(n_87),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_117),
.B1(n_130),
.B2(n_107),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_91),
.B1(n_66),
.B2(n_9),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_91),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_120),
.B(n_103),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_165),
.B(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_144),
.B1(n_132),
.B2(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_144),
.B1(n_146),
.B2(n_132),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_153),
.B1(n_134),
.B2(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_126),
.B1(n_138),
.B2(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_110),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_170),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_113),
.A3(n_123),
.B1(n_129),
.B2(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

XOR2x2_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_118),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_141),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_115),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_146),
.C(n_144),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_118),
.B(n_130),
.Y(n_180)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_199),
.Y(n_208)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_195),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_200),
.B1(n_161),
.B2(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_180),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_159),
.B(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_213),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

OA21x2_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_172),
.B(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_168),
.B1(n_166),
.B2(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_195),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_193),
.C(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_176),
.Y(n_213)
);

AO221x1_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_171),
.B1(n_178),
.B2(n_173),
.C(n_174),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_224),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_182),
.C(n_141),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_210),
.B(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_197),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_194),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_208),
.C(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_232),
.C(n_225),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_203),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_201),
.C(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_220),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_240),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_232),
.A2(n_223),
.B1(n_189),
.B2(n_191),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_206),
.B1(n_184),
.B2(n_198),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_188),
.B1(n_206),
.B2(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_228),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_245),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_188),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_242),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_126),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_237),
.B(n_241),
.C(n_238),
.D(n_198),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_127),
.B(n_128),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_253),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_249),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_128),
.Y(n_256)
);


endmodule