module fake_jpeg_11939_n_521 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_521);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_521;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_0),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_2),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_70),
.Y(n_109)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_2),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_81),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_80),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_3),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_87),
.Y(n_123)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_24),
.B(n_3),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_101),
.B(n_50),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_104),
.B(n_116),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_29),
.B1(n_31),
.B2(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_59),
.A2(n_23),
.B1(n_45),
.B2(n_49),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_110),
.A2(n_49),
.B1(n_47),
.B2(n_30),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_56),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_49),
.B1(n_23),
.B2(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_33),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_131),
.B(n_143),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_42),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_27),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_45),
.B1(n_23),
.B2(n_49),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_62),
.A2(n_31),
.B1(n_22),
.B2(n_47),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_155),
.A2(n_43),
.B1(n_52),
.B2(n_80),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_19),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_60),
.B(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_43),
.Y(n_172)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_134),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_167),
.B(n_183),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_168),
.B(n_172),
.Y(n_251)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_98),
.B1(n_94),
.B2(n_93),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_170),
.A2(n_207),
.B1(n_150),
.B2(n_115),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_171),
.Y(n_275)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_91),
.B1(n_90),
.B2(n_82),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_190),
.B1(n_209),
.B2(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_106),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_176),
.B(n_178),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_177),
.B(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_179),
.A2(n_141),
.B1(n_121),
.B2(n_113),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_109),
.B(n_42),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_199),
.Y(n_226)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_41),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_192),
.C(n_196),
.Y(n_237)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_47),
.B1(n_83),
.B2(n_41),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_102),
.B(n_38),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_105),
.B(n_38),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_122),
.B(n_37),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_129),
.C(n_151),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_37),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_127),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_203),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_36),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_30),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_204),
.Y(n_262)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_206),
.B(n_210),
.Y(n_276)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_108),
.A2(n_30),
.B1(n_19),
.B2(n_80),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_118),
.B(n_3),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_118),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_212),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_107),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_156),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_123),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_218),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_224),
.B1(n_14),
.B2(n_15),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_128),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_219),
.B1(n_213),
.B2(n_195),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_132),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_179),
.A2(n_140),
.B1(n_160),
.B2(n_137),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_243),
.B1(n_249),
.B2(n_253),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_144),
.B1(n_150),
.B2(n_115),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_190),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_141),
.C(n_121),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_262),
.C(n_272),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_176),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_265),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_258),
.B1(n_259),
.B2(n_191),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_140),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_172),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_167),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_254),
.A2(n_267),
.B1(n_270),
.B2(n_253),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_SL g255 ( 
.A1(n_192),
.A2(n_11),
.B(n_12),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_255),
.A2(n_184),
.B1(n_181),
.B2(n_186),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_166),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_175),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_178),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_220),
.A2(n_16),
.B1(n_17),
.B2(n_210),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_196),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_183),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_211),
.A2(n_187),
.B1(n_180),
.B2(n_209),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_278),
.A2(n_285),
.B(n_289),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_242),
.B(n_165),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_281),
.B(n_290),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_237),
.B(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_307),
.C(n_313),
.Y(n_352)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_215),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_204),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_286),
.A2(n_293),
.B(n_306),
.Y(n_342)
);

NOR2x1p5_ASAP7_75t_SL g287 ( 
.A(n_225),
.B(n_174),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_295),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_227),
.A2(n_219),
.B1(n_169),
.B2(n_197),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_288),
.A2(n_302),
.B1(n_323),
.B2(n_241),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_204),
.B(n_188),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_230),
.B(n_173),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_292),
.A2(n_298),
.B1(n_303),
.B2(n_268),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_256),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_198),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_205),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_237),
.B(n_208),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_225),
.A2(n_217),
.B1(n_189),
.B2(n_182),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_240),
.A2(n_221),
.B1(n_275),
.B2(n_263),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_259),
.A2(n_276),
.B1(n_246),
.B2(n_252),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_235),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_236),
.C(n_270),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_226),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_315),
.Y(n_328)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_235),
.A2(n_243),
.B(n_228),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_317),
.B1(n_277),
.B2(n_271),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_233),
.A2(n_247),
.B(n_266),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_314),
.B(n_316),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_240),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_314),
.B(n_293),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_247),
.C(n_267),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_229),
.A2(n_263),
.B(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_254),
.A2(n_230),
.B(n_238),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_249),
.A2(n_258),
.B1(n_239),
.B2(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_231),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_275),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_324),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_238),
.A2(n_261),
.B1(n_244),
.B2(n_277),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_325),
.A2(n_332),
.B1(n_338),
.B2(n_340),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_261),
.B1(n_241),
.B2(n_244),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_327),
.A2(n_335),
.B(n_337),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_279),
.A2(n_248),
.B1(n_268),
.B2(n_250),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_334),
.A2(n_337),
.B1(n_347),
.B2(n_353),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_278),
.A2(n_264),
.B(n_271),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_248),
.B1(n_264),
.B2(n_234),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_279),
.A2(n_234),
.B1(n_248),
.B2(n_310),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_280),
.B1(n_317),
.B2(n_304),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_296),
.B1(n_295),
.B2(n_287),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_341),
.A2(n_358),
.B1(n_340),
.B2(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_297),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_345),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_312),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_298),
.B1(n_278),
.B2(n_306),
.Y(n_347)
);

XNOR2x2_ASAP7_75t_SL g348 ( 
.A(n_289),
.B(n_316),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_342),
.Y(n_375)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_349),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_310),
.A2(n_287),
.B1(n_285),
.B2(n_312),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_286),
.B(n_300),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_361),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_305),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_359),
.C(n_336),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_307),
.A2(n_301),
.B1(n_299),
.B2(n_313),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_299),
.B(n_301),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_360),
.A2(n_322),
.B(n_324),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_320),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_309),
.A2(n_294),
.B1(n_311),
.B2(n_315),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_362),
.A2(n_347),
.B1(n_350),
.B2(n_339),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_283),
.Y(n_363)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_291),
.B(n_321),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_361),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_384),
.Y(n_401)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_372),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_351),
.A2(n_362),
.B(n_353),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_374),
.A2(n_393),
.B1(n_396),
.B2(n_394),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_335),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_350),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_377),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_344),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_389),
.C(n_355),
.Y(n_399)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_380),
.Y(n_405)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_350),
.A2(n_348),
.B(n_326),
.C(n_330),
.Y(n_381)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_352),
.B(n_336),
.CI(n_354),
.CON(n_382),
.SN(n_382)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_391),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_328),
.B(n_364),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_383),
.B(n_395),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_331),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_388),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_387),
.A2(n_389),
.B1(n_373),
.B2(n_371),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_348),
.B(n_326),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_345),
.B(n_349),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_390),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_343),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_356),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_392),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_330),
.A2(n_327),
.B(n_334),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_355),
.B(n_364),
.CI(n_325),
.CON(n_395),
.SN(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_327),
.A2(n_329),
.B1(n_335),
.B2(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_410),
.C(n_392),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_383),
.B(n_343),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_407),
.B(n_427),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_333),
.C(n_346),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_377),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_387),
.A2(n_335),
.B1(n_332),
.B2(n_333),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_419),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_368),
.A2(n_366),
.B1(n_390),
.B2(n_371),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_356),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_422),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_346),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_398),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_423),
.B(n_398),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_424),
.A2(n_425),
.B1(n_426),
.B2(n_417),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_388),
.B1(n_377),
.B2(n_396),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_388),
.B1(n_377),
.B2(n_381),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_385),
.B(n_380),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_408),
.Y(n_428)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_373),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_444),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_434),
.A2(n_440),
.B1(n_448),
.B2(n_449),
.Y(n_459)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_403),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_450),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_424),
.A2(n_368),
.B1(n_379),
.B2(n_384),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_372),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_445),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_445),
.B(n_411),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_365),
.C(n_382),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_447),
.C(n_409),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_382),
.C(n_376),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_425),
.A2(n_379),
.B1(n_376),
.B2(n_395),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_415),
.A2(n_395),
.B1(n_369),
.B2(n_370),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_451),
.B(n_420),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_454),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_422),
.C(n_406),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_415),
.B(n_417),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_458),
.A2(n_465),
.B(n_400),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_443),
.A2(n_426),
.B1(n_412),
.B2(n_413),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_434),
.B1(n_428),
.B2(n_430),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_464),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_441),
.A2(n_413),
.B(n_406),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_419),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_454),
.C(n_453),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_414),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_432),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_440),
.A2(n_418),
.B1(n_420),
.B2(n_412),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_471),
.A2(n_443),
.B1(n_442),
.B2(n_400),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_474),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_435),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_477),
.B1(n_484),
.B2(n_460),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_402),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_483),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_459),
.A2(n_423),
.B1(n_446),
.B2(n_447),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_464),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_461),
.Y(n_497)
);

OAI221xp5_ASAP7_75t_L g480 ( 
.A1(n_468),
.A2(n_451),
.B1(n_439),
.B2(n_448),
.C(n_397),
.Y(n_480)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_481),
.A2(n_465),
.B1(n_458),
.B2(n_470),
.Y(n_487)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_469),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_459),
.A2(n_367),
.B1(n_438),
.B2(n_471),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_463),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_486),
.B(n_455),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_495),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_490),
.Y(n_500)
);

INVx11_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_492),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_484),
.A2(n_455),
.B1(n_467),
.B2(n_462),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_475),
.B1(n_486),
.B2(n_481),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_497),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_463),
.C(n_466),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_478),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_479),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_502),
.B(n_491),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_482),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_506),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_482),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_509),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_500),
.A2(n_489),
.B(n_498),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_497),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_510),
.B(n_511),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_508),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_499),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_515),
.A2(n_516),
.B(n_493),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_512),
.B(n_507),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_499),
.C(n_506),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_513),
.B(n_505),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_519),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_495),
.Y(n_521)
);


endmodule