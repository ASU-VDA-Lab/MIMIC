module fake_aes_1349_n_1622 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_381, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1622);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_381;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1622;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_899;
wire n_716;
wire n_568;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_1611;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_852;
wire n_484;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1432;
wire n_1315;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_659;
wire n_432;
wire n_386;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_1607;
wire n_906;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_16), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_212), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_126), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_12), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_78), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_192), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_33), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_296), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_200), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_141), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_182), .Y(n_393) );
INVxp33_ASAP7_75t_SL g394 ( .A(n_259), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_91), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_249), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_106), .Y(n_397) );
INVxp33_ASAP7_75t_L g398 ( .A(n_41), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_311), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_153), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_202), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_173), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_101), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_66), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_1), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_186), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_109), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_217), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_345), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_11), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_222), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_136), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_171), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_109), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_147), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_243), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_11), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_215), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_82), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_195), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_265), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_245), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_24), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_198), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_62), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_121), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_218), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_157), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_339), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_239), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_350), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_123), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_137), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_84), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_89), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_162), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_145), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_122), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_302), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_310), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_24), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_115), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_348), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_312), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_36), .Y(n_451) );
INVxp33_ASAP7_75t_L g452 ( .A(n_366), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_154), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_85), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_27), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_278), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_264), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_187), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_204), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_352), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_10), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_126), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_163), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_43), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_288), .B(n_103), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_180), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_240), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_137), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_368), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_191), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_263), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_39), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_156), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_233), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_32), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_306), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_129), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_20), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_8), .Y(n_479) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_48), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_50), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_377), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_327), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_357), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_79), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_376), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_83), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_87), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_115), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_274), .Y(n_490) );
INVxp33_ASAP7_75t_L g491 ( .A(n_307), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_78), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_62), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_169), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_193), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_52), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_225), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_279), .Y(n_498) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_111), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_253), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_131), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_362), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_326), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_155), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_328), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_82), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_309), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_149), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_305), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_131), .Y(n_510) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_100), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_68), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_176), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_174), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_5), .Y(n_515) );
INVxp33_ASAP7_75t_L g516 ( .A(n_49), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_48), .B(n_371), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_223), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_111), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_30), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_39), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_207), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_178), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_59), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_161), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_267), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_79), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_28), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_51), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_64), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_224), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_370), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_81), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_160), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_49), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_375), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_167), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_331), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_12), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_63), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_44), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_100), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_0), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_175), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_323), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_221), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_359), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_276), .Y(n_548) );
INVxp33_ASAP7_75t_SL g549 ( .A(n_344), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_281), .Y(n_550) );
BUFx8_ASAP7_75t_SL g551 ( .A(n_1), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_236), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_148), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_363), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_325), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_68), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_333), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_144), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_102), .Y(n_559) );
INVxp33_ASAP7_75t_SL g560 ( .A(n_38), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_297), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_107), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_283), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_354), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_108), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_321), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_361), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_165), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_43), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_103), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_286), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_105), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_216), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_145), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_413), .B(n_0), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_413), .Y(n_576) );
BUFx2_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_452), .B(n_2), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_398), .B(n_2), .Y(n_579) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_413), .B(n_3), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_390), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_426), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_480), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_390), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_390), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_390), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_426), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_400), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_400), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_429), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_390), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_429), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_401), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_428), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_401), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_398), .B(n_3), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_423), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_428), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_432), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_432), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_446), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_452), .B(n_4), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_464), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_516), .B(n_491), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_428), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_446), .B(n_4), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_528), .B(n_5), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_538), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_428), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_516), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_428), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_459), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_464), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_510), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_458), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_604), .B(n_491), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_597), .B(n_459), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_597), .B(n_507), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_576), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_581), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_577), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_610), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_576), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_576), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_581), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_581), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_588), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_604), .B(n_528), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_588), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_608), .B(n_466), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_588), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_597), .B(n_423), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_577), .B(n_604), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_577), .B(n_462), .Y(n_640) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_604), .B(n_507), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_579), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_582), .B(n_508), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_606), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_606), .B(n_462), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_606), .B(n_510), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_582), .B(n_508), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_582), .B(n_537), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_589), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_581), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_608), .B(n_503), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_583), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_645), .A2(n_590), .B(n_592), .C(n_587), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_657), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_624), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
AND3x1_ASAP7_75t_L g662 ( .A(n_617), .B(n_596), .C(n_579), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_639), .B(n_624), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_627), .A2(n_608), .B1(n_488), .B2(n_468), .Y(n_664) );
BUFx3_ASAP7_75t_L g665 ( .A(n_616), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_644), .A2(n_596), .B1(n_579), .B2(n_606), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_621), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_616), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_644), .A2(n_596), .B1(n_579), .B2(n_606), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_616), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_625), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_625), .Y(n_672) );
OAI22xp5_ASAP7_75t_SL g673 ( .A1(n_627), .A2(n_448), .B1(n_421), .B2(n_560), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_647), .Y(n_674) );
AND2x6_ASAP7_75t_L g675 ( .A(n_647), .B(n_596), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_639), .B(n_606), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_626), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_639), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_626), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_623), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_639), .A2(n_602), .B1(n_590), .B2(n_592), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_628), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_636), .B(n_602), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_628), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_639), .B(n_578), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_656), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_655), .B(n_587), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_631), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_631), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_647), .A2(n_590), .B1(n_592), .B2(n_587), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_633), .B(n_649), .Y(n_691) );
BUFx3_ASAP7_75t_L g692 ( .A(n_649), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_645), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_617), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_645), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_645), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_617), .Y(n_697) );
BUFx3_ASAP7_75t_L g698 ( .A(n_649), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_648), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_643), .B(n_599), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_632), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_638), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
CKINVDCx11_ASAP7_75t_R g704 ( .A(n_640), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_632), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_643), .B(n_599), .Y(n_706) );
AND3x1_ASAP7_75t_L g707 ( .A(n_619), .B(n_607), .C(n_575), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_634), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_640), .B(n_408), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_638), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_634), .Y(n_711) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_640), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_649), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_635), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_648), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_638), .B(n_599), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_635), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_637), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_638), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_638), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_649), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_637), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_642), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_648), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_642), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_651), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_651), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_648), .A2(n_600), .B1(n_580), .B2(n_607), .Y(n_728) );
BUFx2_ASAP7_75t_SL g729 ( .A(n_648), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_653), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_633), .B(n_394), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_633), .B(n_394), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g733 ( .A(n_653), .B(n_580), .Y(n_733) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_618), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_715), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_700), .A2(n_646), .B(n_652), .C(n_650), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_676), .A2(n_600), .B1(n_620), .B2(n_619), .Y(n_737) );
BUFx2_ASAP7_75t_L g738 ( .A(n_680), .Y(n_738) );
OAI21x1_ASAP7_75t_L g739 ( .A1(n_661), .A2(n_650), .B(n_646), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_715), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_660), .B(n_620), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_696), .Y(n_742) );
BUFx12f_ASAP7_75t_L g743 ( .A(n_704), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_707), .B(n_652), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_687), .A2(n_706), .B(n_695), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_694), .A2(n_448), .B1(n_421), .B2(n_445), .Y(n_746) );
AND2x6_ASAP7_75t_L g747 ( .A(n_676), .B(n_517), .Y(n_747) );
INVx8_ASAP7_75t_L g748 ( .A(n_675), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_696), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_707), .B(n_575), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_673), .B(n_575), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_715), .Y(n_752) );
INVx4_ASAP7_75t_L g753 ( .A(n_675), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_697), .B(n_489), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_686), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_693), .A2(n_654), .B(n_629), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_662), .B(n_506), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_693), .A2(n_629), .B(n_622), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_675), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g760 ( .A1(n_664), .A2(n_663), .B(n_658), .C(n_716), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_715), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_671), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_665), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_671), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_724), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_675), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_672), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_685), .B(n_560), .Y(n_768) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_678), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_662), .A2(n_445), .B1(n_536), .B2(n_457), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_724), .Y(n_771) );
NAND2x1p5_ASAP7_75t_L g772 ( .A(n_699), .B(n_678), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_675), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_692), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_675), .A2(n_536), .B1(n_552), .B2(n_457), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_676), .A2(n_593), .B1(n_595), .B2(n_589), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_724), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_676), .A2(n_593), .B1(n_595), .B2(n_589), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_724), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_675), .Y(n_780) );
BUFx3_ASAP7_75t_L g781 ( .A(n_692), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_659), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g783 ( .A1(n_731), .A2(n_580), .B(n_549), .Y(n_783) );
NOR2xp67_ASAP7_75t_SL g784 ( .A(n_729), .B(n_456), .Y(n_784) );
NAND2xp33_ASAP7_75t_L g785 ( .A(n_670), .B(n_552), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_691), .B(n_383), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_692), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_672), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_698), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_679), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_698), .Y(n_791) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_670), .Y(n_792) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_699), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_683), .A2(n_541), .B(n_562), .C(n_527), .Y(n_794) );
BUFx3_ASAP7_75t_L g795 ( .A(n_698), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_679), .Y(n_796) );
INVx5_ASAP7_75t_L g797 ( .A(n_699), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_691), .Y(n_798) );
BUFx3_ASAP7_75t_L g799 ( .A(n_670), .Y(n_799) );
BUFx8_ASAP7_75t_SL g800 ( .A(n_685), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_682), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_691), .A2(n_589), .B1(n_595), .B2(n_593), .Y(n_802) );
BUFx2_ASAP7_75t_L g803 ( .A(n_699), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_673), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_729), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_682), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_666), .A2(n_463), .B1(n_514), .B2(n_483), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_701), .Y(n_808) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_670), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_669), .B(n_518), .Y(n_810) );
OR2x6_ASAP7_75t_SL g811 ( .A(n_712), .B(n_385), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_681), .B(n_545), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_719), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_685), .A2(n_496), .B1(n_406), .B2(n_554), .Y(n_814) );
INVx5_ASAP7_75t_L g815 ( .A(n_713), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_691), .A2(n_496), .B1(n_406), .B2(n_511), .C(n_499), .Y(n_816) );
OR2x6_ASAP7_75t_L g817 ( .A(n_702), .B(n_427), .Y(n_817) );
INVx4_ASAP7_75t_L g818 ( .A(n_713), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_674), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_719), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_701), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_685), .B(n_549), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_714), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_709), .B(n_386), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_L g825 ( .A1(n_703), .A2(n_387), .B(n_392), .C(n_389), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_714), .Y(n_826) );
BUFx12f_ASAP7_75t_L g827 ( .A(n_733), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_713), .Y(n_828) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_670), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_702), .B(n_603), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_718), .Y(n_831) );
INVxp67_ASAP7_75t_L g832 ( .A(n_728), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_681), .B(n_417), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_665), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_732), .A2(n_473), .B1(n_435), .B2(n_388), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_713), .A2(n_593), .B1(n_595), .B2(n_589), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_728), .B(n_388), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_713), .A2(n_593), .B1(n_595), .B2(n_589), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g839 ( .A1(n_710), .A2(n_430), .B1(n_427), .B2(n_397), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_695), .A2(n_629), .B(n_622), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_718), .Y(n_841) );
INVx5_ASAP7_75t_L g842 ( .A(n_713), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_722), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_721), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_690), .A2(n_473), .B1(n_435), .B2(n_391), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_733), .B(n_721), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_721), .Y(n_847) );
INVx3_ASAP7_75t_L g848 ( .A(n_665), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_721), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_710), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_720), .B(n_721), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_741), .B(n_733), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_743), .Y(n_853) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_738), .B(n_721), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_775), .A2(n_720), .B1(n_674), .B2(n_667), .Y(n_855) );
INVx6_ASAP7_75t_L g856 ( .A(n_797), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_833), .B(n_722), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_746), .B(n_726), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_751), .B(n_726), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_753), .B(n_674), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_762), .Y(n_861) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_783), .A2(n_614), .B1(n_613), .B2(n_603), .C(n_405), .Y(n_862) );
AO31x2_ASAP7_75t_L g863 ( .A1(n_736), .A2(n_615), .A3(n_586), .B(n_591), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_832), .A2(n_430), .B1(n_530), .B2(n_404), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_747), .A2(n_667), .B1(n_677), .B2(n_661), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_760), .A2(n_708), .B(n_705), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_827), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_768), .A2(n_614), .B1(n_613), .B2(n_603), .C(n_415), .Y(n_868) );
BUFx4f_ASAP7_75t_L g869 ( .A(n_827), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_762), .Y(n_870) );
INVx2_ASAP7_75t_SL g871 ( .A(n_743), .Y(n_871) );
AOI221xp5_ASAP7_75t_SL g872 ( .A1(n_794), .A2(n_711), .B1(n_717), .B2(n_708), .C(n_705), .Y(n_872) );
INVx4_ASAP7_75t_L g873 ( .A(n_748), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_753), .B(n_677), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_768), .A2(n_614), .B1(n_613), .B2(n_437), .C(n_438), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_764), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_747), .A2(n_757), .B1(n_744), .B2(n_750), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_739), .A2(n_717), .B(n_711), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_817), .A2(n_593), .B1(n_601), .B2(n_595), .Y(n_879) );
INVx6_ASAP7_75t_L g880 ( .A(n_797), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_846), .Y(n_881) );
OR2x6_ASAP7_75t_L g882 ( .A(n_748), .B(n_753), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_804), .A2(n_409), .B1(n_439), .B2(n_395), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_817), .Y(n_884) );
NAND2xp5_ASAP7_75t_SL g885 ( .A(n_805), .B(n_670), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_770), .A2(n_684), .B1(n_689), .B2(n_688), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_747), .A2(n_725), .B1(n_727), .B2(n_723), .Y(n_887) );
BUFx2_ASAP7_75t_L g888 ( .A(n_755), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_830), .Y(n_889) );
AOI221x1_ASAP7_75t_SL g890 ( .A1(n_807), .A2(n_443), .B1(n_447), .B2(n_442), .C(n_440), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_755), .B(n_723), .Y(n_891) );
OAI222xp33_ASAP7_75t_L g892 ( .A1(n_804), .A2(n_461), .B1(n_454), .B2(n_472), .C1(n_455), .C2(n_451), .Y(n_892) );
BUFx12f_ASAP7_75t_L g893 ( .A(n_782), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_737), .B(n_745), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_830), .Y(n_895) );
AND2x4_ASAP7_75t_L g896 ( .A(n_797), .B(n_684), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_850), .A2(n_688), .B1(n_689), .B2(n_725), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_747), .A2(n_730), .B1(n_727), .B2(n_493), .Y(n_898) );
INVx1_ASAP7_75t_SL g899 ( .A(n_811), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_737), .B(n_730), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_817), .A2(n_601), .B1(n_612), .B2(n_530), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_830), .Y(n_902) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_748), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_813), .Y(n_904) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_785), .A2(n_475), .B1(n_478), .B2(n_477), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_786), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_764), .Y(n_907) );
AOI21x1_ASAP7_75t_L g908 ( .A1(n_739), .A2(n_557), .B(n_537), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_747), .A2(n_551), .B1(n_668), .B2(n_517), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_822), .A2(n_493), .B1(n_431), .B2(n_601), .Y(n_910) );
INVx1_ASAP7_75t_SL g911 ( .A(n_850), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_798), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_736), .A2(n_668), .B(n_734), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_825), .A2(n_481), .B1(n_487), .B2(n_485), .C(n_479), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_754), .B(n_492), .Y(n_915) );
OAI222xp33_ASAP7_75t_L g916 ( .A1(n_817), .A2(n_519), .B1(n_512), .B2(n_520), .C1(n_515), .C2(n_501), .Y(n_916) );
INVx3_ASAP7_75t_L g917 ( .A(n_797), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_800), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_780), .B(n_521), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_735), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_767), .Y(n_921) );
INVxp67_ASAP7_75t_L g922 ( .A(n_820), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_824), .A2(n_524), .B1(n_535), .B2(n_533), .C(n_529), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_767), .A2(n_612), .B1(n_601), .B2(n_540), .Y(n_924) );
BUFx6f_ASAP7_75t_L g925 ( .A(n_748), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_740), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_752), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_756), .A2(n_557), .B(n_601), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_788), .Y(n_929) );
INVx2_ASAP7_75t_SL g930 ( .A(n_815), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_788), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g932 ( .A1(n_814), .A2(n_539), .B(n_543), .C(n_542), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_790), .Y(n_933) );
OAI21xp5_ASAP7_75t_SL g934 ( .A1(n_812), .A2(n_551), .B(n_556), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_790), .Y(n_935) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_785), .A2(n_559), .B1(n_565), .B2(n_558), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_796), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_816), .B(n_569), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_796), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_822), .A2(n_572), .B1(n_574), .B2(n_570), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_810), .B(n_601), .Y(n_941) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_792), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_824), .A2(n_612), .B(n_393), .C(n_396), .Y(n_943) );
OR2x6_ASAP7_75t_L g944 ( .A(n_759), .B(n_431), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_761), .Y(n_945) );
AOI22xp33_ASAP7_75t_SL g946 ( .A1(n_773), .A2(n_493), .B1(n_431), .B2(n_612), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_837), .B(n_612), .Y(n_947) );
O2A1O1Ixp33_ASAP7_75t_SL g948 ( .A1(n_801), .A2(n_808), .B(n_821), .C(n_806), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_801), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_776), .B(n_612), .Y(n_950) );
O2A1O1Ixp33_ASAP7_75t_SL g951 ( .A1(n_806), .A2(n_465), .B(n_407), .C(n_410), .Y(n_951) );
NOR2xp33_ASAP7_75t_SL g952 ( .A(n_784), .B(n_391), .Y(n_952) );
BUFx3_ASAP7_75t_L g953 ( .A(n_815), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_780), .Y(n_954) );
BUFx3_ASAP7_75t_L g955 ( .A(n_815), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_808), .A2(n_493), .B1(n_431), .B2(n_416), .Y(n_956) );
INVx4_ASAP7_75t_L g957 ( .A(n_842), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_765), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g959 ( .A1(n_766), .A2(n_493), .B1(n_431), .B2(n_534), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_821), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g961 ( .A(n_800), .B(n_548), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_845), .A2(n_573), .B1(n_534), .B2(n_399), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_776), .B(n_399), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_774), .B(n_403), .Y(n_964) );
OR2x6_ASAP7_75t_L g965 ( .A(n_772), .B(n_384), .Y(n_965) );
CKINVDCx11_ASAP7_75t_R g966 ( .A(n_774), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_823), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_758), .A2(n_630), .B(n_622), .Y(n_968) );
OAI21x1_ASAP7_75t_L g969 ( .A1(n_840), .A2(n_826), .B(n_823), .Y(n_969) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_839), .A2(n_419), .B1(n_424), .B2(n_420), .C(n_418), .Y(n_970) );
AND2x4_ASAP7_75t_L g971 ( .A(n_781), .B(n_434), .Y(n_971) );
OAI21x1_ASAP7_75t_L g972 ( .A1(n_826), .A2(n_654), .B(n_630), .Y(n_972) );
INVx3_ASAP7_75t_L g973 ( .A(n_772), .Y(n_973) );
BUFx3_ASAP7_75t_L g974 ( .A(n_815), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_778), .B(n_402), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g976 ( .A1(n_831), .A2(n_573), .B1(n_412), .B2(n_414), .Y(n_976) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_792), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_778), .B(n_402), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_771), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_777), .Y(n_980) );
O2A1O1Ixp33_ASAP7_75t_L g981 ( .A1(n_851), .A2(n_425), .B(n_436), .C(n_433), .Y(n_981) );
INVxp67_ASAP7_75t_L g982 ( .A(n_803), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_802), .B(n_412), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_781), .B(n_467), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_802), .B(n_414), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_831), .A2(n_449), .B1(n_450), .B2(n_444), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_795), .A2(n_470), .B1(n_476), .B2(n_453), .Y(n_987) );
NOR2x1_ASAP7_75t_SL g988 ( .A(n_842), .B(n_482), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_911), .B(n_836), .Y(n_989) );
NOR2xp67_ASAP7_75t_L g990 ( .A(n_867), .B(n_842), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g991 ( .A1(n_890), .A2(n_791), .B1(n_789), .B2(n_787), .C(n_836), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_864), .A2(n_838), .B1(n_779), .B2(n_793), .C(n_835), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_899), .A2(n_842), .B1(n_818), .B2(n_769), .Y(n_993) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_942), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_913), .A2(n_843), .B(n_841), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_904), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_913), .A2(n_843), .B(n_841), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_881), .Y(n_998) );
INVx1_ASAP7_75t_SL g999 ( .A(n_965), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_906), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_877), .A2(n_818), .B1(n_842), .B2(n_819), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_877), .A2(n_819), .B1(n_844), .B2(n_828), .Y(n_1002) );
OAI211xp5_ASAP7_75t_SL g1003 ( .A1(n_934), .A2(n_571), .B(n_564), .C(n_838), .Y(n_1003) );
OAI21xp5_ASAP7_75t_L g1004 ( .A1(n_894), .A2(n_866), .B(n_878), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_852), .B(n_742), .Y(n_1005) );
OAI211xp5_ASAP7_75t_L g1006 ( .A1(n_909), .A2(n_522), .B(n_566), .C(n_497), .Y(n_1006) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_869), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_869), .A2(n_834), .B1(n_848), .B2(n_763), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_973), .B(n_847), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_891), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_857), .Y(n_1011) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_853), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_914), .A2(n_849), .B1(n_834), .B2(n_848), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_965), .A2(n_749), .B1(n_742), .B2(n_848), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_858), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_884), .A2(n_834), .B1(n_763), .B2(n_799), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_864), .A2(n_749), .B1(n_490), .B2(n_494), .C(n_486), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_888), .B(n_763), .Y(n_1018) );
BUFx8_ASAP7_75t_L g1019 ( .A(n_871), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_861), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_914), .A2(n_799), .B1(n_809), .B2(n_792), .Y(n_1021) );
OA21x2_ASAP7_75t_L g1022 ( .A1(n_908), .A2(n_615), .B(n_586), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_884), .A2(n_422), .B1(n_469), .B2(n_441), .Y(n_1023) );
NAND2xp33_ASAP7_75t_R g1024 ( .A(n_965), .B(n_422), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_883), .A2(n_484), .B1(n_505), .B2(n_498), .C(n_495), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_905), .A2(n_809), .B1(n_829), .B2(n_792), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_859), .B(n_809), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_897), .A2(n_829), .B1(n_809), .B2(n_441), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_893), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_883), .A2(n_525), .B1(n_526), .B2(n_513), .C(n_509), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_905), .A2(n_829), .B1(n_532), .B2(n_544), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_901), .A2(n_829), .B1(n_500), .B2(n_502), .Y(n_1032) );
AOI21xp5_ASAP7_75t_L g1033 ( .A1(n_866), .A2(n_734), .B(n_654), .Y(n_1033) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_940), .A2(n_550), .B1(n_561), .B2(n_547), .C(n_531), .Y(n_1034) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_973), .B(n_563), .Y(n_1035) );
NOR2x1_ASAP7_75t_SL g1036 ( .A(n_882), .B(n_567), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_912), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_938), .B(n_469), .Y(n_1038) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_873), .B(n_568), .Y(n_1039) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_932), .A2(n_502), .B(n_504), .C(n_500), .Y(n_1040) );
AND2x4_ASAP7_75t_SL g1041 ( .A(n_918), .B(n_458), .Y(n_1041) );
BUFx4f_ASAP7_75t_L g1042 ( .A(n_856), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_870), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_936), .A2(n_546), .B1(n_553), .B2(n_504), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_936), .A2(n_553), .B1(n_555), .B2(n_546), .Y(n_1045) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_948), .A2(n_734), .B(n_630), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_920), .Y(n_1047) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_892), .A2(n_460), .B1(n_523), .B2(n_471), .C(n_411), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_901), .A2(n_555), .B1(n_615), .B2(n_586), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_922), .B(n_6), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_915), .A2(n_474), .B1(n_458), .B2(n_615), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_887), .A2(n_615), .B1(n_586), .B2(n_591), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_887), .A2(n_591), .B1(n_594), .B2(n_585), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_922), .B(n_6), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_876), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_926), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_963), .B(n_7), .Y(n_1057) );
INVx5_ASAP7_75t_SL g1058 ( .A(n_882), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_894), .A2(n_734), .B(n_591), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_927), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_952), .A2(n_474), .B1(n_458), .B2(n_9), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_923), .A2(n_474), .B1(n_458), .B2(n_594), .C(n_585), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_945), .Y(n_1063) );
A2O1A1Ixp33_ASAP7_75t_L g1064 ( .A1(n_981), .A2(n_879), .B(n_886), .C(n_872), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_975), .B(n_7), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_862), .B(n_474), .C(n_585), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_932), .A2(n_474), .B1(n_584), .B2(n_581), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_953), .Y(n_1068) );
AOI21xp33_ASAP7_75t_L g1069 ( .A1(n_981), .A2(n_594), .B(n_585), .Y(n_1069) );
OAI21xp5_ASAP7_75t_L g1070 ( .A1(n_900), .A2(n_598), .B(n_594), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_879), .A2(n_605), .B1(n_609), .B2(n_598), .Y(n_1071) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_900), .A2(n_605), .B1(n_609), .B2(n_598), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_907), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_875), .B(n_8), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1075 ( .A1(n_875), .A2(n_605), .B(n_609), .C(n_598), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_955), .Y(n_1076) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_988), .A2(n_961), .B1(n_978), .B2(n_944), .Y(n_1077) );
OAI211xp5_ASAP7_75t_L g1078 ( .A1(n_868), .A2(n_609), .B(n_605), .C(n_584), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_923), .A2(n_611), .B1(n_584), .B2(n_581), .C(n_734), .Y(n_1079) );
INVx11_ASAP7_75t_L g1080 ( .A(n_966), .Y(n_1080) );
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_892), .A2(n_611), .B1(n_584), .B2(n_581), .C(n_734), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_898), .A2(n_584), .B1(n_611), .B2(n_581), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_921), .Y(n_1083) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_862), .B(n_611), .C(n_584), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_983), .B(n_9), .Y(n_1085) );
AOI221xp5_ASAP7_75t_SL g1086 ( .A1(n_910), .A2(n_611), .B1(n_584), .B2(n_641), .C(n_618), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_985), .A2(n_14), .B1(n_10), .B2(n_13), .Y(n_1087) );
AOI222xp33_ASAP7_75t_L g1088 ( .A1(n_868), .A2(n_13), .B1(n_14), .B2(n_15), .C1(n_16), .C2(n_17), .Y(n_1088) );
A2O1A1Ixp33_ASAP7_75t_L g1089 ( .A1(n_898), .A2(n_910), .B(n_943), .C(n_941), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_929), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_982), .B(n_15), .Y(n_1091) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_916), .A2(n_17), .B1(n_18), .B2(n_19), .C1(n_20), .C2(n_21), .Y(n_1092) );
BUFx2_ASAP7_75t_L g1093 ( .A(n_974), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_976), .A2(n_611), .B1(n_584), .B2(n_618), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_982), .B(n_18), .Y(n_1095) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_930), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_944), .A2(n_22), .B1(n_19), .B2(n_21), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_958), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_916), .A2(n_611), .B1(n_584), .B2(n_641), .C(n_618), .Y(n_1099) );
INVx2_ASAP7_75t_SL g1100 ( .A(n_856), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g1101 ( .A1(n_944), .A2(n_611), .B1(n_584), .B2(n_25), .Y(n_1101) );
INVx1_ASAP7_75t_SL g1102 ( .A(n_896), .Y(n_1102) );
AND2x4_ASAP7_75t_SL g1103 ( .A(n_957), .B(n_611), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_856), .A2(n_611), .B1(n_25), .B2(n_22), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_979), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_970), .A2(n_641), .B1(n_618), .B2(n_27), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_986), .B(n_23), .Y(n_1107) );
INVx3_ASAP7_75t_L g1108 ( .A(n_957), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_970), .A2(n_641), .B1(n_618), .B2(n_28), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_865), .A2(n_29), .B1(n_23), .B2(n_26), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_986), .A2(n_641), .B1(n_618), .B2(n_30), .C(n_31), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_931), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_933), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_919), .A2(n_641), .B1(n_31), .B2(n_26), .Y(n_1114) );
AND2x6_ASAP7_75t_L g1115 ( .A(n_903), .B(n_29), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_935), .Y(n_1116) );
AOI22xp33_ASAP7_75t_SL g1117 ( .A1(n_880), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_937), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_946), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_855), .A2(n_38), .B1(n_35), .B2(n_37), .Y(n_1120) );
OAI222xp33_ASAP7_75t_L g1121 ( .A1(n_962), .A2(n_37), .B1(n_40), .B2(n_41), .C1(n_42), .C2(n_44), .Y(n_1121) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_964), .B(n_40), .Y(n_1122) );
OAI21x1_ASAP7_75t_L g1123 ( .A1(n_968), .A2(n_641), .B(n_150), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_919), .A2(n_46), .B1(n_42), .B2(n_45), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_924), .A2(n_45), .B1(n_46), .B2(n_47), .C(n_50), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_882), .A2(n_52), .B1(n_47), .B2(n_51), .Y(n_1126) );
AO31x2_ASAP7_75t_L g1127 ( .A1(n_956), .A2(n_55), .A3(n_53), .B(n_54), .Y(n_1127) );
A2O1A1Ixp33_ASAP7_75t_L g1128 ( .A1(n_889), .A2(n_55), .B(n_53), .C(n_54), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_1024), .A2(n_976), .B1(n_962), .B2(n_946), .C(n_959), .Y(n_1129) );
NOR2xp33_ASAP7_75t_R g1130 ( .A(n_1029), .B(n_917), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1131 ( .A(n_1005), .B(n_896), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_999), .B(n_939), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_996), .Y(n_1133) );
INVx4_ASAP7_75t_SL g1134 ( .A(n_1115), .Y(n_1134) );
OAI31xp33_ASAP7_75t_SL g1135 ( .A1(n_999), .A2(n_854), .A3(n_959), .B(n_956), .Y(n_1135) );
NAND2x1p5_ASAP7_75t_L g1136 ( .A(n_1042), .B(n_873), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1020), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1010), .B(n_964), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1043), .Y(n_1139) );
OAI211xp5_ASAP7_75t_L g1140 ( .A1(n_1092), .A2(n_987), .B(n_951), .C(n_950), .Y(n_1140) );
OAI21xp33_ASAP7_75t_L g1141 ( .A1(n_1048), .A2(n_984), .B(n_971), .Y(n_1141) );
OAI21xp5_ASAP7_75t_SL g1142 ( .A1(n_1041), .A2(n_924), .B(n_917), .Y(n_1142) );
AO21x2_ASAP7_75t_L g1143 ( .A1(n_1004), .A2(n_928), .B(n_885), .Y(n_1143) );
AOI21xp5_ASAP7_75t_L g1144 ( .A1(n_1014), .A2(n_1033), .B(n_995), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_1011), .A2(n_895), .B1(n_902), .B2(n_947), .C(n_980), .Y(n_1145) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_1019), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_990), .Y(n_1147) );
INVx3_ASAP7_75t_L g1148 ( .A(n_1058), .Y(n_1148) );
NAND2xp5_ASAP7_75t_SL g1149 ( .A(n_1077), .B(n_1032), .Y(n_1149) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_1092), .A2(n_960), .B(n_967), .C(n_949), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_998), .Y(n_1151) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1058), .Y(n_1152) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_1036), .A2(n_880), .B1(n_874), .B2(n_971), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_1003), .A2(n_874), .B1(n_984), .B2(n_880), .Y(n_1154) );
OAI221xp5_ASAP7_75t_SL g1155 ( .A1(n_1107), .A2(n_1088), .B1(n_1025), .B2(n_1030), .C(n_1085), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_1057), .A2(n_860), .B1(n_954), .B2(n_925), .Y(n_1156) );
OAI221xp5_ASAP7_75t_L g1157 ( .A1(n_1064), .A2(n_954), .B1(n_925), .B2(n_903), .C(n_977), .Y(n_1157) );
AND2x4_ASAP7_75t_SL g1158 ( .A(n_1007), .B(n_903), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1065), .A2(n_860), .B1(n_925), .B2(n_969), .Y(n_1159) );
OR2x6_ASAP7_75t_L g1160 ( .A(n_1076), .B(n_942), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1047), .Y(n_1161) );
NAND4xp25_ASAP7_75t_L g1162 ( .A(n_1088), .B(n_58), .C(n_56), .D(n_57), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1091), .B(n_1095), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_1044), .A2(n_977), .B1(n_942), .B2(n_863), .C(n_59), .Y(n_1164) );
OA21x2_ASAP7_75t_L g1165 ( .A1(n_1004), .A2(n_972), .B(n_863), .Y(n_1165) );
AND2x2_ASAP7_75t_SL g1166 ( .A(n_1042), .B(n_977), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1015), .B(n_863), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1168 ( .A(n_1050), .Y(n_1168) );
BUFx6f_ASAP7_75t_L g1169 ( .A(n_994), .Y(n_1169) );
OAI33xp33_ASAP7_75t_L g1170 ( .A1(n_1087), .A2(n_56), .A3(n_57), .B1(n_58), .B2(n_60), .B3(n_61), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1074), .A2(n_63), .B1(n_60), .B2(n_61), .Y(n_1171) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_1019), .Y(n_1172) );
OAI33xp33_ASAP7_75t_L g1173 ( .A1(n_1110), .A2(n_64), .A3(n_65), .B1(n_66), .B2(n_67), .B3(n_69), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_1122), .A2(n_69), .B1(n_65), .B2(n_67), .Y(n_1174) );
NAND3xp33_ASAP7_75t_L g1175 ( .A(n_1104), .B(n_70), .C(n_71), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1055), .Y(n_1176) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_1032), .A2(n_1040), .B1(n_1013), .B2(n_1045), .Y(n_1177) );
INVx2_ASAP7_75t_SL g1178 ( .A(n_1080), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1056), .Y(n_1179) );
OAI22xp5_ASAP7_75t_SL g1180 ( .A1(n_1117), .A2(n_72), .B1(n_70), .B2(n_71), .Y(n_1180) );
OAI31xp33_ASAP7_75t_L g1181 ( .A1(n_1006), .A2(n_74), .A3(n_72), .B(n_73), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1060), .Y(n_1182) );
AO21x2_ASAP7_75t_L g1183 ( .A1(n_997), .A2(n_73), .B(n_74), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1031), .A2(n_77), .B1(n_75), .B2(n_76), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1054), .B(n_75), .Y(n_1185) );
OA21x2_ASAP7_75t_L g1186 ( .A1(n_1086), .A2(n_151), .B(n_146), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1037), .B(n_76), .Y(n_1187) );
NAND4xp25_ASAP7_75t_SL g1188 ( .A(n_1125), .B(n_77), .C(n_80), .D(n_81), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g1189 ( .A1(n_1119), .A2(n_80), .B1(n_83), .B2(n_84), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_1121), .A2(n_85), .B1(n_86), .B2(n_87), .C(n_88), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1035), .B(n_86), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1192 ( .A(n_1108), .B(n_88), .Y(n_1192) );
NOR3xp33_ASAP7_75t_L g1193 ( .A(n_1034), .B(n_89), .C(n_90), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1073), .Y(n_1194) );
BUFx3_ASAP7_75t_L g1195 ( .A(n_1093), .Y(n_1195) );
OA21x2_ASAP7_75t_L g1196 ( .A1(n_1086), .A2(n_158), .B(n_152), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1197 ( .A1(n_1059), .A2(n_164), .B(n_159), .Y(n_1197) );
INVx3_ASAP7_75t_L g1198 ( .A(n_1058), .Y(n_1198) );
NOR2x1_ASAP7_75t_L g1199 ( .A(n_1119), .B(n_90), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_989), .B(n_91), .Y(n_1200) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_1000), .A2(n_92), .B1(n_93), .B2(n_94), .C(n_95), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1068), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1063), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1083), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1035), .B(n_92), .Y(n_1205) );
OAI211xp5_ASAP7_75t_L g1206 ( .A1(n_1023), .A2(n_93), .B(n_94), .C(n_95), .Y(n_1206) );
OR2x6_ASAP7_75t_L g1207 ( .A(n_1108), .B(n_96), .Y(n_1207) );
OAI31xp33_ASAP7_75t_L g1208 ( .A1(n_1126), .A2(n_96), .A3(n_97), .B(n_98), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1090), .Y(n_1209) );
OAI21xp5_ASAP7_75t_L g1210 ( .A1(n_1089), .A2(n_97), .B(n_98), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1096), .B(n_99), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1021), .A2(n_99), .B1(n_101), .B2(n_102), .Y(n_1212) );
OAI31xp33_ASAP7_75t_SL g1213 ( .A1(n_1110), .A2(n_104), .A3(n_105), .B(n_106), .Y(n_1213) );
OAI31xp33_ASAP7_75t_L g1214 ( .A1(n_1120), .A2(n_104), .A3(n_107), .B(n_108), .Y(n_1214) );
BUFx3_ASAP7_75t_L g1215 ( .A(n_1012), .Y(n_1215) );
OAI33xp33_ASAP7_75t_L g1216 ( .A1(n_1097), .A2(n_110), .A3(n_112), .B1(n_113), .B2(n_114), .B3(n_116), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1112), .Y(n_1217) );
OAI33xp33_ASAP7_75t_L g1218 ( .A1(n_1061), .A2(n_110), .A3(n_112), .B1(n_113), .B2(n_114), .B3(n_116), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1018), .B(n_117), .Y(n_1219) );
OAI33xp33_ASAP7_75t_L g1220 ( .A1(n_1098), .A2(n_117), .A3(n_118), .B1(n_119), .B2(n_120), .B3(n_121), .Y(n_1220) );
NAND3xp33_ASAP7_75t_L g1221 ( .A(n_1128), .B(n_118), .C(n_119), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1105), .B(n_120), .Y(n_1222) );
INVx4_ASAP7_75t_L g1223 ( .A(n_1115), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_1106), .A2(n_122), .B1(n_123), .B2(n_124), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1113), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1116), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1038), .B(n_124), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_992), .A2(n_125), .B1(n_127), .B2(n_128), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1118), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1102), .B(n_125), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_1102), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1232 ( .A(n_1039), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1002), .B(n_127), .Y(n_1233) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_1017), .A2(n_128), .B1(n_129), .B2(n_130), .C(n_132), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g1235 ( .A1(n_991), .A2(n_130), .B1(n_132), .B2(n_133), .C(n_134), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_1111), .A2(n_133), .B1(n_134), .B2(n_135), .C(n_136), .Y(n_1236) );
BUFx3_ASAP7_75t_L g1237 ( .A(n_1100), .Y(n_1237) );
OAI211xp5_ASAP7_75t_L g1238 ( .A1(n_1124), .A2(n_135), .B(n_138), .C(n_139), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1039), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_1109), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_1240) );
AOI222xp33_ASAP7_75t_L g1241 ( .A1(n_1115), .A2(n_140), .B1(n_141), .B2(n_142), .C1(n_143), .C2(n_144), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_997), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1127), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1127), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_1115), .A2(n_143), .B1(n_166), .B2(n_168), .Y(n_1245) );
AOI21xp5_ASAP7_75t_L g1246 ( .A1(n_1046), .A2(n_381), .B(n_172), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1001), .A2(n_170), .B1(n_177), .B2(n_179), .Y(n_1247) );
OAI211xp5_ASAP7_75t_L g1248 ( .A1(n_1067), .A2(n_181), .B(n_183), .C(n_184), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_1081), .A2(n_185), .B1(n_188), .B2(n_189), .Y(n_1249) );
AO21x2_ASAP7_75t_L g1250 ( .A1(n_1070), .A2(n_1123), .B(n_1084), .Y(n_1250) );
BUFx3_ASAP7_75t_L g1251 ( .A(n_1103), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1027), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1127), .Y(n_1253) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1009), .Y(n_1254) );
NAND2xp5_ASAP7_75t_SL g1255 ( .A(n_993), .B(n_1008), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1009), .Y(n_1256) );
AND2x6_ASAP7_75t_L g1257 ( .A(n_994), .B(n_190), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_1062), .A2(n_194), .B1(n_196), .B2(n_197), .C(n_199), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1151), .Y(n_1259) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_1242), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1202), .B(n_1132), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1262 ( .A(n_1172), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1133), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1231), .Y(n_1264) );
NAND3xp33_ASAP7_75t_L g1265 ( .A(n_1241), .B(n_1051), .C(n_1114), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1161), .B(n_1026), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_1129), .A2(n_1155), .B1(n_1207), .B2(n_1153), .Y(n_1267) );
INVx4_ASAP7_75t_L g1268 ( .A(n_1134), .Y(n_1268) );
INVx3_ASAP7_75t_L g1269 ( .A(n_1223), .Y(n_1269) );
INVxp67_ASAP7_75t_SL g1270 ( .A(n_1252), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1179), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1191), .B(n_1049), .Y(n_1272) );
INVx2_ASAP7_75t_SL g1273 ( .A(n_1146), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1205), .B(n_1028), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1138), .B(n_1101), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1200), .B(n_1070), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1131), .B(n_1016), .Y(n_1277) );
AOI33xp33_ASAP7_75t_L g1278 ( .A1(n_1182), .A2(n_1094), .A3(n_1099), .B1(n_1075), .B2(n_1069), .B3(n_1078), .Y(n_1278) );
NAND3xp33_ASAP7_75t_L g1279 ( .A(n_1213), .B(n_1052), .C(n_1053), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1203), .Y(n_1280) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1165), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1131), .B(n_1071), .Y(n_1282) );
AOI22xp33_ASAP7_75t_SL g1283 ( .A1(n_1129), .A2(n_1082), .B1(n_1079), .B2(n_1071), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1225), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1226), .Y(n_1285) );
INVx2_ASAP7_75t_SL g1286 ( .A(n_1130), .Y(n_1286) );
BUFx2_ASAP7_75t_SL g1287 ( .A(n_1215), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1134), .B(n_994), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1289 ( .A(n_1162), .B(n_1052), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_1155), .A2(n_1053), .B1(n_1072), .B2(n_1066), .C(n_1082), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1211), .B(n_1072), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1229), .Y(n_1292) );
NAND4xp25_ASAP7_75t_L g1293 ( .A(n_1174), .B(n_201), .C(n_203), .D(n_205), .Y(n_1293) );
BUFx3_ASAP7_75t_L g1294 ( .A(n_1251), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1185), .B(n_1022), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1137), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1139), .Y(n_1297) );
OAI221xp5_ASAP7_75t_L g1298 ( .A1(n_1141), .A2(n_1022), .B1(n_208), .B2(n_209), .C(n_210), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1168), .B(n_206), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1176), .Y(n_1300) );
AOI22xp33_ASAP7_75t_SL g1301 ( .A1(n_1223), .A2(n_211), .B1(n_213), .B2(n_214), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1167), .Y(n_1302) );
AOI22xp5_ASAP7_75t_L g1303 ( .A1(n_1140), .A2(n_219), .B1(n_220), .B2(n_226), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1195), .B(n_227), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1232), .B(n_380), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1239), .B(n_228), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1194), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1204), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1163), .B(n_1145), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1145), .B(n_379), .Y(n_1310) );
AND2x4_ASAP7_75t_L g1311 ( .A(n_1134), .B(n_229), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1209), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1217), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1187), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1315 ( .A(n_1160), .B(n_230), .Y(n_1315) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1165), .Y(n_1316) );
NAND3xp33_ASAP7_75t_SL g1317 ( .A(n_1142), .B(n_231), .C(n_232), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_1207), .A2(n_234), .B1(n_235), .B2(n_237), .Y(n_1318) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1243), .Y(n_1319) );
AO21x2_ASAP7_75t_L g1320 ( .A1(n_1144), .A2(n_238), .B(n_241), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_1188), .A2(n_242), .B1(n_244), .B2(n_246), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1187), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1222), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1207), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1244), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1192), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1230), .B(n_247), .Y(n_1327) );
OA21x2_ASAP7_75t_L g1328 ( .A1(n_1144), .A2(n_248), .B(n_250), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1219), .B(n_378), .Y(n_1329) );
OAI22xp5_ASAP7_75t_SL g1330 ( .A1(n_1178), .A2(n_251), .B1(n_252), .B2(n_254), .Y(n_1330) );
AND2x4_ASAP7_75t_L g1331 ( .A(n_1160), .B(n_255), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1332 ( .A(n_1167), .B(n_256), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_1188), .A2(n_257), .B1(n_258), .B2(n_260), .Y(n_1333) );
INVx1_ASAP7_75t_SL g1334 ( .A(n_1237), .Y(n_1334) );
NAND2xp5_ASAP7_75t_SL g1335 ( .A(n_1135), .B(n_261), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1254), .B(n_373), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1192), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1147), .Y(n_1338) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1253), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_1190), .B(n_262), .C(n_266), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1233), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1227), .B(n_268), .Y(n_1342) );
AOI211xp5_ASAP7_75t_L g1343 ( .A1(n_1180), .A2(n_269), .B(n_270), .C(n_271), .Y(n_1343) );
AOI31xp33_ASAP7_75t_L g1344 ( .A1(n_1190), .A2(n_272), .A3(n_273), .B(n_275), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1256), .B(n_277), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1233), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1143), .Y(n_1347) );
OAI211xp5_ASAP7_75t_L g1348 ( .A1(n_1201), .A2(n_280), .B(n_282), .C(n_284), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1166), .B(n_285), .Y(n_1349) );
AND2x4_ASAP7_75t_L g1350 ( .A(n_1169), .B(n_1160), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_1199), .A2(n_287), .B1(n_289), .B2(n_290), .Y(n_1351) );
INVx3_ASAP7_75t_L g1352 ( .A(n_1136), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1183), .Y(n_1353) );
AOI221xp5_ASAP7_75t_L g1354 ( .A1(n_1189), .A2(n_291), .B1(n_292), .B2(n_293), .C(n_294), .Y(n_1354) );
OAI31xp33_ASAP7_75t_L g1355 ( .A1(n_1140), .A2(n_295), .A3(n_298), .B(n_300), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1201), .B(n_301), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_1193), .A2(n_303), .B1(n_304), .B2(n_308), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1235), .B(n_313), .Y(n_1358) );
AOI221xp5_ASAP7_75t_L g1359 ( .A1(n_1234), .A2(n_314), .B1(n_315), .B2(n_316), .C(n_317), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1183), .Y(n_1360) );
OAI31xp33_ASAP7_75t_L g1361 ( .A1(n_1206), .A2(n_318), .A3(n_319), .B(n_320), .Y(n_1361) );
NAND3xp33_ASAP7_75t_L g1362 ( .A(n_1181), .B(n_322), .C(n_324), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1149), .B(n_372), .Y(n_1363) );
NOR3xp33_ASAP7_75t_L g1364 ( .A(n_1206), .B(n_1234), .C(n_1238), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1148), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1148), .Y(n_1366) );
AND2x4_ASAP7_75t_L g1367 ( .A(n_1152), .B(n_329), .Y(n_1367) );
BUFx2_ASAP7_75t_L g1368 ( .A(n_1152), .Y(n_1368) );
INVx2_ASAP7_75t_L g1369 ( .A(n_1143), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1284), .B(n_1235), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1259), .Y(n_1371) );
OAI31xp33_ASAP7_75t_L g1372 ( .A1(n_1267), .A2(n_1238), .A3(n_1208), .B(n_1136), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1285), .B(n_1210), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1292), .B(n_1228), .Y(n_1374) );
O2A1O1Ixp33_ASAP7_75t_L g1375 ( .A1(n_1335), .A2(n_1184), .B(n_1240), .C(n_1224), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1261), .B(n_1270), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1309), .B(n_1171), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1263), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1302), .B(n_1159), .Y(n_1379) );
OAI21xp5_ASAP7_75t_L g1380 ( .A1(n_1344), .A2(n_1335), .B(n_1340), .Y(n_1380) );
AOI221x1_ASAP7_75t_L g1381 ( .A1(n_1317), .A2(n_1197), .B1(n_1246), .B2(n_1221), .C(n_1198), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1302), .B(n_1250), .Y(n_1382) );
NOR3xp33_ASAP7_75t_L g1383 ( .A(n_1317), .B(n_1220), .C(n_1216), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1319), .B(n_1250), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1319), .B(n_1169), .Y(n_1385) );
INVx2_ASAP7_75t_L g1386 ( .A(n_1339), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1339), .B(n_1169), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1271), .Y(n_1388) );
OAI31xp33_ASAP7_75t_L g1389 ( .A1(n_1324), .A2(n_1214), .A3(n_1157), .B(n_1175), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1280), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1338), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1270), .Y(n_1392) );
OR2x6_ASAP7_75t_L g1393 ( .A(n_1268), .B(n_1255), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1264), .B(n_1156), .Y(n_1394) );
INVx1_ASAP7_75t_SL g1395 ( .A(n_1287), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1264), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1323), .B(n_1198), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1296), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1326), .B(n_1216), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1314), .B(n_1236), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1297), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1300), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1353), .B(n_1360), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1307), .B(n_1150), .Y(n_1404) );
NAND3xp33_ASAP7_75t_L g1405 ( .A(n_1364), .B(n_1236), .C(n_1245), .Y(n_1405) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1281), .Y(n_1406) );
INVxp33_ASAP7_75t_L g1407 ( .A(n_1350), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1325), .B(n_1186), .Y(n_1408) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_1260), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1308), .Y(n_1410) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_1294), .Y(n_1411) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1281), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1312), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1313), .B(n_1150), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1334), .B(n_1164), .Y(n_1415) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_1350), .Y(n_1416) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1316), .Y(n_1417) );
INVx2_ASAP7_75t_L g1418 ( .A(n_1316), .Y(n_1418) );
OAI21xp33_ASAP7_75t_L g1419 ( .A1(n_1364), .A2(n_1157), .B(n_1164), .Y(n_1419) );
BUFx2_ASAP7_75t_L g1420 ( .A(n_1294), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1322), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1337), .Y(n_1422) );
AOI21xp5_ASAP7_75t_L g1423 ( .A1(n_1355), .A2(n_1196), .B(n_1186), .Y(n_1423) );
INVx1_ASAP7_75t_SL g1424 ( .A(n_1262), .Y(n_1424) );
AOI22xp5_ASAP7_75t_L g1425 ( .A1(n_1289), .A2(n_1154), .B1(n_1177), .B2(n_1212), .Y(n_1425) );
AOI21xp33_ASAP7_75t_L g1426 ( .A1(n_1289), .A2(n_1248), .B(n_1247), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1325), .B(n_1196), .Y(n_1427) );
AOI21xp5_ASAP7_75t_SL g1428 ( .A1(n_1311), .A2(n_1258), .B(n_1257), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1275), .B(n_1170), .Y(n_1429) );
NAND4xp25_ASAP7_75t_L g1430 ( .A(n_1265), .B(n_1258), .C(n_1197), .D(n_1249), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1295), .B(n_1257), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1266), .Y(n_1432) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1347), .Y(n_1433) );
NAND5xp2_ASAP7_75t_L g1434 ( .A(n_1343), .B(n_1248), .C(n_1246), .D(n_1170), .E(n_1173), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1276), .B(n_1158), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_1341), .B(n_1220), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1260), .B(n_1257), .Y(n_1437) );
NAND2xp5_ASAP7_75t_SL g1438 ( .A(n_1269), .B(n_1257), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1332), .B(n_1257), .Y(n_1439) );
INVx3_ASAP7_75t_L g1440 ( .A(n_1268), .Y(n_1440) );
OAI31xp33_ASAP7_75t_L g1441 ( .A1(n_1293), .A2(n_1173), .A3(n_1218), .B(n_334), .Y(n_1441) );
BUFx2_ASAP7_75t_SL g1442 ( .A(n_1286), .Y(n_1442) );
NAND4xp25_ASAP7_75t_L g1443 ( .A(n_1321), .B(n_1218), .C(n_332), .D(n_335), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1346), .B(n_330), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1272), .B(n_336), .Y(n_1445) );
NAND4xp25_ASAP7_75t_L g1446 ( .A(n_1321), .B(n_337), .C(n_338), .D(n_340), .Y(n_1446) );
INVx2_ASAP7_75t_L g1447 ( .A(n_1369), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1282), .B(n_341), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1291), .B(n_342), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1274), .B(n_343), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1365), .Y(n_1451) );
OAI31xp33_ASAP7_75t_L g1452 ( .A1(n_1299), .A2(n_346), .A3(n_347), .B(n_349), .Y(n_1452) );
AOI31xp67_ASAP7_75t_SL g1453 ( .A1(n_1310), .A2(n_351), .A3(n_355), .B(n_356), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1273), .B(n_358), .Y(n_1454) );
AND2x4_ASAP7_75t_L g1455 ( .A(n_1269), .B(n_360), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1392), .Y(n_1456) );
NAND3xp33_ASAP7_75t_L g1457 ( .A(n_1429), .B(n_1366), .C(n_1333), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1391), .B(n_1376), .Y(n_1458) );
INVxp67_ASAP7_75t_L g1459 ( .A(n_1409), .Y(n_1459) );
AND3x2_ASAP7_75t_L g1460 ( .A(n_1428), .B(n_1311), .C(n_1368), .Y(n_1460) );
AOI22xp5_ASAP7_75t_L g1461 ( .A1(n_1429), .A2(n_1277), .B1(n_1299), .B2(n_1356), .Y(n_1461) );
OAI21xp33_ASAP7_75t_SL g1462 ( .A1(n_1438), .A2(n_1333), .B(n_1304), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1411), .B(n_1350), .Y(n_1463) );
AOI21xp33_ASAP7_75t_L g1464 ( .A1(n_1399), .A2(n_1363), .B(n_1305), .Y(n_1464) );
O2A1O1Ixp33_ASAP7_75t_L g1465 ( .A1(n_1372), .A2(n_1377), .B(n_1397), .C(n_1400), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1432), .B(n_1332), .Y(n_1466) );
INVxp67_ASAP7_75t_L g1467 ( .A(n_1409), .Y(n_1467) );
HB1xp67_ASAP7_75t_L g1468 ( .A(n_1403), .Y(n_1468) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_1405), .A2(n_1279), .B1(n_1283), .B2(n_1362), .Y(n_1469) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_1428), .A2(n_1361), .B(n_1298), .Y(n_1470) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1406), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1396), .B(n_1332), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1371), .B(n_1262), .Y(n_1473) );
NAND2x1_ASAP7_75t_SL g1474 ( .A(n_1440), .B(n_1352), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1378), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1420), .B(n_1327), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1388), .Y(n_1477) );
OAI21xp33_ASAP7_75t_L g1478 ( .A1(n_1419), .A2(n_1303), .B(n_1283), .Y(n_1478) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1390), .B(n_1306), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_1421), .B(n_1352), .Y(n_1480) );
NOR3xp33_ASAP7_75t_L g1481 ( .A(n_1443), .B(n_1348), .C(n_1330), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1422), .B(n_1342), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1416), .B(n_1288), .Y(n_1483) );
OR2x2_ASAP7_75t_L g1484 ( .A(n_1398), .B(n_1331), .Y(n_1484) );
CKINVDCx16_ASAP7_75t_R g1485 ( .A(n_1442), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1401), .Y(n_1486) );
AOI32xp33_ASAP7_75t_L g1487 ( .A1(n_1395), .A2(n_1349), .A3(n_1301), .B1(n_1367), .B2(n_1331), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1416), .B(n_1288), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1402), .Y(n_1489) );
INVx1_ASAP7_75t_SL g1490 ( .A(n_1424), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1410), .B(n_1315), .Y(n_1491) );
NOR2xp33_ASAP7_75t_L g1492 ( .A(n_1415), .B(n_1329), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1413), .Y(n_1493) );
INVx1_ASAP7_75t_SL g1494 ( .A(n_1454), .Y(n_1494) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1394), .B(n_1315), .Y(n_1495) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_1403), .Y(n_1496) );
INVx2_ASAP7_75t_L g1497 ( .A(n_1406), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1399), .B(n_1290), .Y(n_1498) );
INVx2_ASAP7_75t_SL g1499 ( .A(n_1440), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1451), .B(n_1358), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1386), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1386), .Y(n_1502) );
NOR3xp33_ASAP7_75t_L g1503 ( .A(n_1446), .B(n_1318), .C(n_1359), .Y(n_1503) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1379), .B(n_1336), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1407), .B(n_1367), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1404), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1379), .B(n_1320), .Y(n_1507) );
XNOR2xp5_ASAP7_75t_L g1508 ( .A(n_1425), .B(n_1301), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1407), .B(n_1345), .Y(n_1509) );
OR2x2_ASAP7_75t_L g1510 ( .A(n_1414), .B(n_1320), .Y(n_1510) );
INVxp67_ASAP7_75t_L g1511 ( .A(n_1382), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1373), .B(n_1351), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_1468), .B(n_1418), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1475), .Y(n_1514) );
AND2x4_ASAP7_75t_L g1515 ( .A(n_1468), .B(n_1437), .Y(n_1515) );
AOI21xp5_ASAP7_75t_L g1516 ( .A1(n_1470), .A2(n_1438), .B(n_1380), .Y(n_1516) );
NAND2xp33_ASAP7_75t_L g1517 ( .A(n_1487), .B(n_1439), .Y(n_1517) );
INVxp67_ASAP7_75t_L g1518 ( .A(n_1506), .Y(n_1518) );
OAI21xp33_ASAP7_75t_SL g1519 ( .A1(n_1474), .A2(n_1439), .B(n_1393), .Y(n_1519) );
INVx2_ASAP7_75t_L g1520 ( .A(n_1471), .Y(n_1520) );
O2A1O1Ixp33_ASAP7_75t_L g1521 ( .A1(n_1498), .A2(n_1389), .B(n_1383), .C(n_1375), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1477), .Y(n_1522) );
NOR2xp33_ASAP7_75t_L g1523 ( .A(n_1508), .B(n_1436), .Y(n_1523) );
XNOR2xp5_ASAP7_75t_L g1524 ( .A(n_1490), .B(n_1393), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1486), .Y(n_1525) );
INVx1_ASAP7_75t_SL g1526 ( .A(n_1485), .Y(n_1526) );
INVx2_ASAP7_75t_L g1527 ( .A(n_1471), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1489), .Y(n_1528) );
XNOR2xp5_ASAP7_75t_L g1529 ( .A(n_1476), .B(n_1393), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1463), .B(n_1431), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_1496), .B(n_1382), .Y(n_1531) );
INVx1_ASAP7_75t_SL g1532 ( .A(n_1473), .Y(n_1532) );
INVx1_ASAP7_75t_SL g1533 ( .A(n_1458), .Y(n_1533) );
INVx1_ASAP7_75t_SL g1534 ( .A(n_1496), .Y(n_1534) );
XNOR2x2_ASAP7_75t_L g1535 ( .A(n_1494), .B(n_1437), .Y(n_1535) );
NOR2xp33_ASAP7_75t_L g1536 ( .A(n_1465), .B(n_1370), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1456), .B(n_1384), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1493), .Y(n_1538) );
INVxp33_ASAP7_75t_L g1539 ( .A(n_1481), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1459), .Y(n_1540) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1459), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1511), .B(n_1384), .Y(n_1542) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_1461), .A2(n_1453), .B1(n_1440), .B2(n_1435), .Y(n_1543) );
OAI22xp33_ASAP7_75t_L g1544 ( .A1(n_1484), .A2(n_1444), .B1(n_1430), .B2(n_1381), .Y(n_1544) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1497), .Y(n_1545) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1467), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_1511), .B(n_1387), .Y(n_1547) );
OR2x2_ASAP7_75t_L g1548 ( .A(n_1495), .B(n_1418), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1501), .Y(n_1549) );
INVxp67_ASAP7_75t_L g1550 ( .A(n_1492), .Y(n_1550) );
XNOR2xp5_ASAP7_75t_L g1551 ( .A(n_1460), .B(n_1448), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1502), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1504), .B(n_1417), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1480), .Y(n_1554) );
INVxp67_ASAP7_75t_L g1555 ( .A(n_1492), .Y(n_1555) );
AOI221xp5_ASAP7_75t_L g1556 ( .A1(n_1469), .A2(n_1374), .B1(n_1434), .B2(n_1441), .C(n_1426), .Y(n_1556) );
O2A1O1Ixp33_ASAP7_75t_L g1557 ( .A1(n_1478), .A2(n_1450), .B(n_1445), .C(n_1449), .Y(n_1557) );
OAI21xp5_ASAP7_75t_L g1558 ( .A1(n_1481), .A2(n_1455), .B(n_1351), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1472), .B(n_1412), .Y(n_1559) );
XOR2x2_ASAP7_75t_L g1560 ( .A(n_1460), .B(n_1455), .Y(n_1560) );
O2A1O1Ixp5_ASAP7_75t_L g1561 ( .A1(n_1457), .A2(n_1455), .B(n_1423), .C(n_1431), .Y(n_1561) );
OAI21xp33_ASAP7_75t_L g1562 ( .A1(n_1469), .A2(n_1385), .B(n_1357), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1497), .Y(n_1563) );
OA22x2_ASAP7_75t_L g1564 ( .A1(n_1499), .A2(n_1505), .B1(n_1488), .B2(n_1483), .Y(n_1564) );
INVxp67_ASAP7_75t_L g1565 ( .A(n_1510), .Y(n_1565) );
AOI211xp5_ASAP7_75t_SL g1566 ( .A1(n_1464), .A2(n_1453), .B(n_1408), .C(n_1427), .Y(n_1566) );
AND3x1_ASAP7_75t_L g1567 ( .A(n_1503), .B(n_1452), .C(n_1357), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1509), .B(n_1412), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1491), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g1570 ( .A1(n_1466), .A2(n_1417), .B1(n_1328), .B2(n_1354), .Y(n_1570) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1500), .Y(n_1571) );
AOI22xp5_ASAP7_75t_L g1572 ( .A1(n_1517), .A2(n_1539), .B1(n_1536), .B2(n_1567), .Y(n_1572) );
NAND3xp33_ASAP7_75t_L g1573 ( .A(n_1521), .B(n_1539), .C(n_1556), .Y(n_1573) );
O2A1O1Ixp33_ASAP7_75t_L g1574 ( .A1(n_1536), .A2(n_1517), .B(n_1516), .C(n_1523), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1540), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1541), .Y(n_1576) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1513), .Y(n_1577) );
OAI21xp5_ASAP7_75t_L g1578 ( .A1(n_1561), .A2(n_1523), .B(n_1558), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g1579 ( .A1(n_1544), .A2(n_1557), .B(n_1562), .Y(n_1579) );
AOI22xp33_ASAP7_75t_L g1580 ( .A1(n_1564), .A2(n_1543), .B1(n_1544), .B2(n_1550), .Y(n_1580) );
A2O1A1Ixp33_ASAP7_75t_L g1581 ( .A1(n_1519), .A2(n_1526), .B(n_1561), .C(n_1566), .Y(n_1581) );
AOI22xp5_ASAP7_75t_L g1582 ( .A1(n_1564), .A2(n_1550), .B1(n_1555), .B2(n_1515), .Y(n_1582) );
AOI22xp5_ASAP7_75t_L g1583 ( .A1(n_1555), .A2(n_1515), .B1(n_1569), .B2(n_1518), .Y(n_1583) );
AOI221xp5_ASAP7_75t_L g1584 ( .A1(n_1571), .A2(n_1565), .B1(n_1534), .B2(n_1533), .C(n_1554), .Y(n_1584) );
NOR2x1_ASAP7_75t_SL g1585 ( .A(n_1547), .B(n_1560), .Y(n_1585) );
INVxp67_ASAP7_75t_L g1586 ( .A(n_1524), .Y(n_1586) );
AOI22xp33_ASAP7_75t_SL g1587 ( .A1(n_1535), .A2(n_1462), .B1(n_1515), .B2(n_1532), .Y(n_1587) );
XNOR2x1_ASAP7_75t_L g1588 ( .A(n_1529), .B(n_1551), .Y(n_1588) );
BUFx6f_ASAP7_75t_L g1589 ( .A(n_1573), .Y(n_1589) );
INVxp67_ASAP7_75t_SL g1590 ( .A(n_1574), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g1591 ( .A(n_1575), .Y(n_1591) );
AOI221xp5_ASAP7_75t_L g1592 ( .A1(n_1579), .A2(n_1565), .B1(n_1525), .B2(n_1538), .C(n_1522), .Y(n_1592) );
OAI21xp5_ASAP7_75t_L g1593 ( .A1(n_1572), .A2(n_1570), .B(n_1503), .Y(n_1593) );
A2O1A1Ixp33_ASAP7_75t_L g1594 ( .A1(n_1581), .A2(n_1531), .B(n_1528), .C(n_1514), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1578), .B(n_1546), .Y(n_1595) );
OAI21xp33_ASAP7_75t_L g1596 ( .A1(n_1580), .A2(n_1542), .B(n_1553), .Y(n_1596) );
AOI22xp5_ASAP7_75t_L g1597 ( .A1(n_1587), .A2(n_1568), .B1(n_1512), .B2(n_1530), .Y(n_1597) );
NAND4xp25_ASAP7_75t_L g1598 ( .A(n_1582), .B(n_1507), .C(n_1482), .D(n_1479), .Y(n_1598) );
AOI22xp5_ASAP7_75t_L g1599 ( .A1(n_1586), .A2(n_1552), .B1(n_1549), .B2(n_1537), .Y(n_1599) );
AOI31xp33_ASAP7_75t_L g1600 ( .A1(n_1590), .A2(n_1588), .A3(n_1584), .B(n_1585), .Y(n_1600) );
AND4x1_ASAP7_75t_L g1601 ( .A(n_1593), .B(n_1583), .C(n_1576), .D(n_1535), .Y(n_1601) );
OAI22xp33_ASAP7_75t_SL g1602 ( .A1(n_1597), .A2(n_1577), .B1(n_1563), .B2(n_1559), .Y(n_1602) );
AO22x2_ASAP7_75t_L g1603 ( .A1(n_1595), .A2(n_1545), .B1(n_1527), .B2(n_1520), .Y(n_1603) );
NAND5xp2_ASAP7_75t_L g1604 ( .A(n_1594), .B(n_1427), .C(n_1408), .D(n_1328), .E(n_1278), .Y(n_1604) );
BUFx2_ASAP7_75t_L g1605 ( .A(n_1591), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1606 ( .A(n_1592), .B(n_1548), .Y(n_1606) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1599), .Y(n_1607) );
XNOR2xp5_ASAP7_75t_L g1608 ( .A(n_1601), .B(n_1598), .Y(n_1608) );
NAND2xp5_ASAP7_75t_SL g1609 ( .A(n_1600), .B(n_1589), .Y(n_1609) );
INVxp67_ASAP7_75t_L g1610 ( .A(n_1605), .Y(n_1610) );
NOR4xp75_ASAP7_75t_L g1611 ( .A(n_1606), .B(n_1596), .C(n_1328), .D(n_365), .Y(n_1611) );
AOI22xp5_ASAP7_75t_SL g1612 ( .A1(n_1602), .A2(n_1545), .B1(n_1527), .B2(n_1520), .Y(n_1612) );
XNOR2xp5_ASAP7_75t_L g1613 ( .A(n_1609), .B(n_1607), .Y(n_1613) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_1608), .A2(n_1603), .B1(n_1602), .B2(n_1604), .Y(n_1614) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1610), .Y(n_1615) );
INVx2_ASAP7_75t_L g1616 ( .A(n_1612), .Y(n_1616) );
AND3x2_ASAP7_75t_L g1617 ( .A(n_1615), .B(n_1611), .C(n_1603), .Y(n_1617) );
OR3x1_ASAP7_75t_L g1618 ( .A(n_1613), .B(n_1278), .C(n_364), .Y(n_1618) );
AOI22xp5_ASAP7_75t_L g1619 ( .A1(n_1618), .A2(n_1614), .B1(n_1616), .B2(n_1433), .Y(n_1619) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1617), .Y(n_1620) );
BUFx2_ASAP7_75t_L g1621 ( .A(n_1620), .Y(n_1621) );
AOI21xp5_ASAP7_75t_L g1622 ( .A1(n_1621), .A2(n_1619), .B(n_1447), .Y(n_1622) );
endmodule