module real_jpeg_33035_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_1),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_4),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_5),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_5),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_5),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_6),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_6),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_7),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_78),
.Y(n_77)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_8),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_8),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

NAND2x2_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_10),
.B(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_85),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_12),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_12),
.B(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_15),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_15),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_15),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_15),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_15),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_171),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_170),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2x1_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

NAND2x1p5_ASAP7_75t_L g170 ( 
.A(n_20),
.B(n_127),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_66),
.C(n_104),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_22),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.C(n_49),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_23),
.B(n_274),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_24),
.B(n_28),
.C(n_31),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_30),
.Y(n_136)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_30),
.Y(n_183)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_30),
.Y(n_253)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_37),
.A2(n_38),
.B1(n_49),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_40),
.B(n_46),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_43),
.Y(n_186)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_47),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_47),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_47),
.Y(n_242)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_49),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_60),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_50),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_264)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_55),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_59),
.Y(n_205)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_67),
.B(n_105),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_82),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_68),
.B(n_83),
.C(n_90),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.C(n_77),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_69),
.B(n_280),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g239 ( 
.A1(n_70),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_70),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_70),
.B(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_72),
.B(n_77),
.Y(n_280)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_89),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_87),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_95),
.C(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_103),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_123),
.C(n_125),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_115),
.C(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_111),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_154),
.Y(n_127)
);

XOR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_153),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

HB1xp67_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_161),
.A2(n_162),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_283),
.B(n_288),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_271),
.B(n_282),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_246),
.B(n_269),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_221),
.B(n_245),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_198),
.B(n_220),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_193),
.B(n_197),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_192),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_212),
.B2(n_213),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_206),
.C(n_212),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_216),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_223),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_236),
.C(n_239),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_265),
.C(n_268),
.Y(n_246)
);

O2A1O1Ixp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_248),
.B(n_268),
.C(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_254),
.C(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_262),
.C(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_281),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_277),
.C(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_286),
.Y(n_288)
);


endmodule