module fake_netlist_6_1728_n_73 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_73);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_73;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_24;
wire n_18;
wire n_21;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_72;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_48;
wire n_47;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_3),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_0),
.B1(n_12),
.B2(n_14),
.Y(n_31)
);

AND2x6_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_2),
.Y(n_32)
);

NAND2x1p5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_23),
.Y(n_38)
);

O2A1O1Ixp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_20),
.B(n_29),
.C(n_24),
.Y(n_39)
);

NAND2x1p5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_23),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_20),
.B(n_29),
.C(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_31),
.B1(n_20),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_25),
.B1(n_19),
.B2(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_18),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_30),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_25),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_45),
.B(n_48),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_52),
.B1(n_53),
.B2(n_51),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_53),
.B(n_47),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_53),
.B(n_47),
.Y(n_64)
);

OAI321xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_25),
.A3(n_21),
.B1(n_5),
.B2(n_22),
.C(n_26),
.Y(n_65)
);

AOI221xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.C(n_21),
.Y(n_66)
);

NOR2x1p5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_64),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_26),
.B(n_27),
.C(n_65),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

XNOR2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_26),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_R g71 ( 
.A(n_70),
.B(n_27),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_69),
.B(n_27),
.Y(n_72)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_27),
.Y(n_73)
);


endmodule