module fake_jpeg_19563_n_145 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_74),
.Y(n_84)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_70),
.B1(n_59),
.B2(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_67),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_69),
.B1(n_63),
.B2(n_57),
.Y(n_86)
);

OAI211xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_89),
.B(n_48),
.C(n_61),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_53),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_53),
.CON(n_88),
.SN(n_88)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_60),
.B1(n_50),
.B2(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_96),
.Y(n_105)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_99),
.B1(n_100),
.B2(n_84),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_95),
.B(n_64),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_48),
.B1(n_58),
.B2(n_3),
.Y(n_108)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_1),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_106),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_20),
.B(n_44),
.C(n_43),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_18),
.C(n_40),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_12),
.C(n_33),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_2),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_17),
.A3(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_45),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_120),
.Y(n_128)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_126),
.B1(n_21),
.B2(n_24),
.C(n_27),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_125),
.B1(n_105),
.B2(n_111),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_111),
.B1(n_112),
.B2(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_133),
.C(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_128),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_126),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_118),
.C(n_130),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_28),
.B(n_6),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_6),
.Y(n_145)
);


endmodule