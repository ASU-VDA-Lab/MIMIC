module fake_jpeg_6715_n_81 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_53),
.B1(n_42),
.B2(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_44),
.B1(n_50),
.B2(n_49),
.Y(n_59)
);

XNOR2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_38),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_58),
.B1(n_61),
.B2(n_57),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.C(n_8),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_6),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_9),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_10),
.C(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_13),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_19),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.C1(n_26),
.C2(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_28),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_29),
.C(n_31),
.Y(n_81)
);


endmodule