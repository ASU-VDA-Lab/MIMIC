module fake_netlist_6_3507_n_1984 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1984);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1984;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_95),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_65),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_35),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

INVxp67_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_64),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_80),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_135),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_13),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_61),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_66),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_109),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_19),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_57),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_12),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_130),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_36),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_101),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_49),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_22),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_133),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_152),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_81),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_97),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_51),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_157),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_102),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_153),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_127),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_13),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_96),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_117),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_86),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_100),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_68),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_9),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_55),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_34),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_119),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_142),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_57),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_17),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_129),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_49),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_113),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_105),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_29),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_18),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_160),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_118),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_171),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_134),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_108),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_141),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_59),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_166),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_65),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_190),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_31),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_79),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_187),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_77),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_56),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_174),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_89),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_186),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_70),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_73),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_136),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_83),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_45),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_54),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_98),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_45),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_17),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_106),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_110),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_155),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_116),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_188),
.Y(n_323)
);

BUFx8_ASAP7_75t_SL g324 ( 
.A(n_84),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_33),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_56),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_131),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_147),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_144),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_90),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_145),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_21),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_183),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_40),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_143),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_3),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_162),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_39),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_18),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_128),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_0),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_61),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_1),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_62),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_104),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_46),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_121),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_37),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_112),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_26),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_149),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_194),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_185),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_126),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_164),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_66),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_25),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_115),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_54),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_189),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_58),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_5),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_103),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_12),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_36),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_123),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_122),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_11),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_44),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_167),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_92),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_85),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_43),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_24),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_156),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_50),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_41),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_78),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_27),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_38),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_111),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_151),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_52),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_175),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_16),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_93),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_51),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_39),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_168),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_74),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_62),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_30),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_225),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_294),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_215),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_294),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_226),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_228),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_237),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_294),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_393),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_230),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_205),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_294),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_294),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_231),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_236),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g412 ( 
.A(n_200),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_294),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_294),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_238),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_239),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_244),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_247),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_252),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_218),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_200),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_359),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_265),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_270),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_324),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_227),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_271),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_272),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_232),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_233),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_255),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_202),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_343),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_243),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_343),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_248),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_202),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_343),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_343),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_354),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_251),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_279),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_280),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_284),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_253),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_208),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_240),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_257),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_220),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_246),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_262),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_259),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_260),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_274),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_276),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_285),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_220),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_278),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_264),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_220),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_286),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_300),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_304),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_281),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_298),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_299),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_315),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_220),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_208),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_267),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_336),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_341),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_316),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_346),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_349),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_210),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_273),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_367),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_220),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_367),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_305),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_351),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_366),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_487),
.A2(n_222),
.B1(n_394),
.B2(n_210),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_403),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_440),
.B(n_201),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_451),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_417),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_R g516 ( 
.A(n_396),
.B(n_340),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_456),
.B(n_201),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_405),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_433),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_436),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_203),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_412),
.A2(n_249),
.B1(n_379),
.B2(n_325),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_203),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_401),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_438),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_400),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_206),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_443),
.B(n_206),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_423),
.B(n_235),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_450),
.B(n_280),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_404),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_408),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_409),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_413),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_446),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_429),
.B(n_235),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_414),
.B(n_245),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_437),
.B(n_214),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_401),
.B(n_292),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_402),
.B(n_212),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_496),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_496),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_492),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_459),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g560 ( 
.A(n_463),
.B(n_214),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_448),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_462),
.B(n_296),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_465),
.B(n_296),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_454),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_471),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_474),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_402),
.B(n_245),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_406),
.B(n_292),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_309),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_468),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_552),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_372),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_406),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_552),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_560),
.A2(n_309),
.B1(n_326),
.B2(n_317),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_562),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_522),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_539),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_573),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_524),
.Y(n_593)
);

OAI22x1_ASAP7_75t_L g594 ( 
.A1(n_519),
.A2(n_399),
.B1(n_490),
.B2(n_483),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_573),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_542),
.B(n_410),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_553),
.B(n_372),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_571),
.B(n_410),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_517),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_576),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_576),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_548),
.B(n_458),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_533),
.B(n_411),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_411),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_567),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_R g608 ( 
.A(n_533),
.B(n_415),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_568),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_568),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_560),
.A2(n_309),
.B1(n_326),
.B2(n_317),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_545),
.B(n_425),
.C(n_407),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_529),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_512),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_529),
.Y(n_618)
);

CKINVDCx6p67_ASAP7_75t_R g619 ( 
.A(n_523),
.Y(n_619)
);

INVxp33_ASAP7_75t_L g620 ( 
.A(n_531),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_530),
.B(n_415),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_539),
.B(n_217),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_513),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_549),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_549),
.A2(n_362),
.B1(n_490),
.B2(n_483),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_514),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_549),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_572),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_567),
.Y(n_636)
);

BUFx6f_ASAP7_75t_SL g637 ( 
.A(n_505),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_520),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_572),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_572),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_527),
.B(n_418),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_527),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_535),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_540),
.B(n_418),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_460),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_574),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_536),
.B(n_420),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_540),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_574),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_541),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_502),
.B(n_420),
.Y(n_657)
);

BUFx16f_ASAP7_75t_R g658 ( 
.A(n_503),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_516),
.A2(n_219),
.B1(n_224),
.B2(n_212),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_534),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_545),
.B(n_480),
.C(n_427),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_574),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_505),
.B(n_421),
.Y(n_664)
);

INVx4_ASAP7_75t_SL g665 ( 
.A(n_574),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_546),
.A2(n_234),
.B(n_217),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_526),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_546),
.A2(n_362),
.B1(n_386),
.B2(n_382),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_521),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_499),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_521),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_505),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_564),
.B(n_421),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_505),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_500),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_504),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

BUFx6f_ASAP7_75t_SL g679 ( 
.A(n_538),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_507),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_268),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_424),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_507),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_575),
.B(n_497),
.C(n_498),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_509),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_534),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_575),
.B(n_478),
.C(n_472),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_510),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_510),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_554),
.B(n_466),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_504),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_537),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_538),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_504),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_526),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_526),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_526),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_547),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_543),
.Y(n_705)
);

AND3x2_ASAP7_75t_L g706 ( 
.A(n_564),
.B(n_269),
.C(n_268),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_543),
.B(n_424),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_538),
.B(n_479),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_504),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_543),
.B(n_430),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_575),
.A2(n_385),
.B1(n_361),
.B2(n_269),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_538),
.B(n_485),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_543),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_565),
.B(n_430),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_431),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_506),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_556),
.A2(n_486),
.B1(n_489),
.B2(n_488),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_544),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_558),
.B(n_481),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_547),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_506),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_544),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_559),
.A2(n_361),
.B1(n_312),
.B2(n_385),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_561),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_566),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_506),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_544),
.B(n_431),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_506),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_579),
.B(n_434),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_581),
.B(n_544),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_435),
.C(n_434),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_544),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_590),
.B(n_650),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_591),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_719),
.B(n_435),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_582),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_590),
.A2(n_484),
.B1(n_473),
.B2(n_467),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_589),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_637),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_592),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_650),
.B(n_491),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_719),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_586),
.B(n_551),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_657),
.A2(n_312),
.B1(n_293),
.B2(n_307),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_591),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_627),
.B(n_551),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_591),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_583),
.A2(n_557),
.B(n_556),
.C(n_580),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_595),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_616),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_672),
.B(n_555),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_695),
.B(n_566),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_672),
.B(n_555),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_674),
.B(n_698),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_645),
.B(n_455),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_708),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_605),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_627),
.B(n_555),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_634),
.Y(n_762)
);

NOR3xp33_ASAP7_75t_L g763 ( 
.A(n_604),
.B(n_470),
.C(n_457),
.Y(n_763)
);

INVx6_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_605),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_605),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_621),
.B(n_246),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_621),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_674),
.B(n_457),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_634),
.B(n_246),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_SL g772 ( 
.A(n_620),
.B(n_432),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_698),
.B(n_470),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_724),
.B(n_475),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_588),
.A2(n_246),
.B1(n_263),
.B2(n_355),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_603),
.B(n_475),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_697),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_648),
.B(n_476),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_697),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_609),
.B(n_476),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_684),
.B(n_477),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_609),
.B(n_477),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_628),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_708),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_598),
.B(n_596),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_595),
.Y(n_787)
);

O2A1O1Ixp5_ASAP7_75t_L g788 ( 
.A1(n_624),
.A2(n_501),
.B(n_511),
.C(n_199),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_624),
.B(n_246),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_707),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_617),
.B(n_495),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_666),
.A2(n_557),
.B(n_580),
.C(n_577),
.Y(n_792)
);

INVx8_ASAP7_75t_L g793 ( 
.A(n_637),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_617),
.B(n_495),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_593),
.B(n_615),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_501),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_712),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_712),
.B(n_563),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_729),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_600),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_623),
.B(n_501),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_710),
.B(n_196),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_624),
.B(n_263),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_600),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_652),
.B(n_321),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_625),
.B(n_511),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_628),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_625),
.B(n_511),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_585),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_350),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_602),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_673),
.A2(n_352),
.B1(n_392),
.B2(n_310),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_664),
.B(n_318),
.C(n_313),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_660),
.B(n_219),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_727),
.B(n_196),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_626),
.B(n_204),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_630),
.B(n_558),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_631),
.B(n_250),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_632),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_624),
.B(n_263),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_660),
.B(n_224),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_602),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_671),
.B(n_263),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_632),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_599),
.B(n_569),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_633),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_671),
.B(n_263),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_638),
.B(n_254),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_638),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_L g831 ( 
.A(n_683),
.B(n_220),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_692),
.B(n_578),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_639),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_628),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_599),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_671),
.B(n_355),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_636),
.A2(n_508),
.B(n_506),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_622),
.B(n_197),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_639),
.B(n_256),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_599),
.B(n_569),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_643),
.B(n_355),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_643),
.B(n_355),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_R g843 ( 
.A(n_593),
.B(n_615),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_644),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_613),
.A2(n_333),
.B1(n_287),
.B2(n_283),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_601),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_646),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_646),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_597),
.B(n_197),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_687),
.B(n_198),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_653),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_687),
.B(n_198),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_655),
.B(n_355),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_655),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_659),
.B(n_220),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_628),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_670),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_715),
.A2(n_320),
.B1(n_319),
.B2(n_275),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_692),
.B(n_578),
.Y(n_859)
);

AO22x2_ASAP7_75t_L g860 ( 
.A1(n_689),
.A2(n_266),
.B1(n_290),
.B2(n_258),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_614),
.B(n_207),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_584),
.B(n_207),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_670),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_601),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_675),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_675),
.B(n_577),
.Y(n_866)
);

INVx8_ASAP7_75t_L g867 ( 
.A(n_637),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_676),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_669),
.B(n_211),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_661),
.B(n_332),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_683),
.A2(n_220),
.B1(n_306),
.B2(n_314),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_661),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_669),
.B(n_211),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_680),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_678),
.B(n_291),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_678),
.B(n_302),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_681),
.B(n_327),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_614),
.B(n_334),
.C(n_339),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_720),
.B(n_347),
.C(n_370),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_618),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_680),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_682),
.B(n_353),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_681),
.B(n_364),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_685),
.B(n_369),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_685),
.B(n_508),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_706),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_720),
.B(n_371),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_825),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_825),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_733),
.B(n_790),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_760),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_820),
.B(n_658),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_827),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_872),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_830),
.Y(n_895)
);

BUFx4f_ASAP7_75t_L g896 ( 
.A(n_741),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_736),
.B(n_704),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_SL g898 ( 
.A(n_743),
.B(n_376),
.C(n_375),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_775),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_843),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_843),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_830),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_798),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_757),
.B(n_682),
.Y(n_904)
);

AOI221xp5_ASAP7_75t_SL g905 ( 
.A1(n_845),
.A2(n_594),
.B1(n_668),
.B2(n_711),
.C(n_723),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_SL g906 ( 
.A(n_835),
.B(n_799),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_760),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_786),
.A2(n_679),
.B1(n_683),
.B2(n_705),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_833),
.Y(n_909)
);

OR2x2_ASAP7_75t_SL g910 ( 
.A(n_814),
.B(n_662),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_759),
.B(n_662),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_815),
.B(n_686),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_SL g913 ( 
.A(n_743),
.B(n_376),
.C(n_375),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_815),
.B(n_686),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_819),
.B(n_688),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_826),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_833),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_760),
.B(n_702),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_760),
.B(n_702),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_748),
.A2(n_679),
.B1(n_718),
.B2(n_690),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_880),
.B(n_618),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_744),
.B(n_619),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_741),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_762),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_844),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_777),
.B(n_704),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_784),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_770),
.B(n_702),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_844),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_847),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_770),
.B(n_651),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_738),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_772),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_SL g934 ( 
.A(n_878),
.B(n_388),
.C(n_378),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_741),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_784),
.Y(n_936)
);

NOR2x1p5_ASAP7_75t_L g937 ( 
.A(n_822),
.B(n_619),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_848),
.B(n_693),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_886),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_847),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_778),
.B(n_780),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_785),
.B(n_797),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_784),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_851),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_758),
.B(n_694),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_770),
.B(n_651),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_810),
.A2(n_725),
.B1(n_594),
.B2(n_378),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_793),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_762),
.B(n_770),
.Y(n_949)
);

NOR2x1p5_ASAP7_75t_L g950 ( 
.A(n_887),
.B(n_725),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_851),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_795),
.B(n_704),
.Y(n_952)
);

BUFx2_ASAP7_75t_SL g953 ( 
.A(n_755),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_776),
.A2(n_747),
.B1(n_854),
.B2(n_805),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_854),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_863),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_735),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_793),
.B(n_717),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_863),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_732),
.A2(n_718),
.B(n_663),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_758),
.B(n_647),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_771),
.A2(n_767),
.B(n_803),
.C(n_789),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_784),
.B(n_654),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_793),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_781),
.B(n_388),
.Y(n_965)
);

BUFx8_ASAP7_75t_SL g966 ( 
.A(n_870),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_779),
.B(n_647),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_748),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_807),
.B(n_654),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_874),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_783),
.A2(n_794),
.B(n_791),
.C(n_805),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_768),
.Y(n_972)
);

NOR2x2_ASAP7_75t_L g973 ( 
.A(n_747),
.B(n_704),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_840),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_779),
.A2(n_683),
.B1(n_701),
.B2(n_722),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_735),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_832),
.B(n_649),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_810),
.A2(n_683),
.B1(n_701),
.B2(n_722),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_832),
.B(n_649),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_817),
.B(n_717),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_731),
.B(n_700),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_769),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_881),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_776),
.A2(n_683),
.B1(n_717),
.B2(n_394),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_737),
.Y(n_985)
);

INVx3_ASAP7_75t_SL g986 ( 
.A(n_867),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_807),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_734),
.A2(n_700),
.B1(n_703),
.B2(n_705),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_867),
.B(n_667),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_859),
.B(n_656),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_773),
.B(n_703),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_866),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_866),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_768),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_859),
.B(n_713),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_807),
.B(n_656),
.Y(n_996)
);

AND3x1_ASAP7_75t_L g997 ( 
.A(n_879),
.B(n_390),
.C(n_395),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_867),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_750),
.B(n_713),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_SL g1000 ( 
.A1(n_753),
.A2(n_838),
.B1(n_764),
.B2(n_395),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_747),
.A2(n_860),
.B1(n_871),
.B2(n_730),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_765),
.B(n_585),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_737),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_764),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_746),
.A2(n_667),
.B(n_691),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_865),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_764),
.B(n_213),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_860),
.A2(n_390),
.B1(n_241),
.B2(n_261),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_739),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_868),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_766),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_869),
.B(n_585),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_869),
.B(n_587),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_834),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_774),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_782),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_873),
.B(n_587),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_846),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_834),
.B(n_667),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_763),
.B(n_861),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_739),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_873),
.B(n_587),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_882),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_856),
.B(n_667),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_838),
.A2(n_587),
.B1(n_607),
.B2(n_691),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_SL g1027 ( 
.A(n_812),
.B(n_342),
.C(n_360),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_730),
.B(n_607),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_740),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_740),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_742),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_862),
.B(n_607),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_862),
.A2(n_607),
.B1(n_691),
.B2(n_721),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_742),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_882),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_745),
.Y(n_1037)
);

OAI21xp33_ASAP7_75t_SL g1038 ( 
.A1(n_789),
.A2(n_691),
.B(n_610),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_871),
.A2(n_241),
.B1(n_242),
.B2(n_261),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_813),
.B(n_850),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_745),
.A2(n_241),
.B1(n_242),
.B2(n_261),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_752),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_752),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_846),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_852),
.B(n_665),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_849),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_802),
.B(n_610),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_787),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_787),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_856),
.B(n_665),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_751),
.B(n_635),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_864),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_816),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_864),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_796),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_818),
.B(n_611),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_754),
.A2(n_612),
.B(n_642),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_831),
.B(n_213),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_800),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_829),
.B(n_611),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_839),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_800),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_756),
.B(n_216),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_876),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_917),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_927),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_921),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_971),
.B(n_858),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_917),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_R g1070 ( 
.A(n_901),
.B(n_801),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_926),
.B(n_792),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_945),
.B(n_804),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_SL g1073 ( 
.A1(n_945),
.A2(n_884),
.B(n_877),
.C(n_875),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1004),
.B(n_809),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_897),
.B(n_855),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_890),
.B(n_855),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_927),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_899),
.B(n_767),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_980),
.B(n_804),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_954),
.A2(n_821),
.B1(n_803),
.B2(n_771),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_965),
.A2(n_1027),
.B(n_1021),
.C(n_961),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_927),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_929),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_954),
.A2(n_821),
.B1(n_811),
.B2(n_823),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_894),
.B(n_749),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1032),
.A2(n_761),
.B(n_612),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_921),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_SL g1088 ( 
.A1(n_932),
.A2(n_947),
.B1(n_910),
.B2(n_900),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_903),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1005),
.A2(n_885),
.B(n_788),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_927),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_929),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_916),
.B(n_876),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_974),
.B(n_811),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_967),
.A2(n_883),
.B(n_853),
.C(n_842),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_962),
.A2(n_823),
.B(n_883),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_982),
.A2(n_806),
.B1(n_808),
.B2(n_277),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_853),
.B(n_842),
.C(n_841),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_984),
.A2(n_841),
.B1(n_836),
.B2(n_828),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_888),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1020),
.A2(n_612),
.B(n_837),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_1051),
.A2(n_836),
.B(n_828),
.C(n_824),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1040),
.A2(n_329),
.B1(n_345),
.B2(n_337),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_952),
.B(n_216),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_984),
.A2(n_1001),
.B1(n_1039),
.B2(n_1009),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_889),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_963),
.A2(n_824),
.B(n_728),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_912),
.B(n_629),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_914),
.B(n_629),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_977),
.B(n_640),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_933),
.B(n_365),
.C(n_363),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_957),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_991),
.A2(n_728),
.B(n_726),
.C(n_721),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_957),
.Y(n_1114)
);

CKINVDCx8_ASAP7_75t_R g1115 ( 
.A(n_953),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_941),
.A2(n_640),
.B(n_641),
.C(n_635),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1057),
.A2(n_726),
.B(n_716),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1064),
.A2(n_716),
.B(n_709),
.C(n_699),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1053),
.B(n_1017),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_958),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_979),
.A2(n_635),
.B(n_699),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_902),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1025),
.A2(n_612),
.B(n_642),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1025),
.A2(n_612),
.B(n_642),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_960),
.A2(n_642),
.B(n_508),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_911),
.B(n_1024),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_987),
.B(n_677),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_952),
.B(n_223),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_985),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_909),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1061),
.B(n_677),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_925),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1001),
.A2(n_357),
.B1(n_358),
.B2(n_344),
.Y(n_1133)
);

NAND2x1_ASAP7_75t_L g1134 ( 
.A(n_987),
.B(n_677),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_995),
.B(n_696),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_990),
.B(n_696),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1013),
.A2(n_508),
.B(n_696),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_940),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1014),
.A2(n_696),
.B(n_665),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_944),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1018),
.A2(n_665),
.B(n_209),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1022),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1046),
.B(n_223),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_951),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1023),
.A2(n_330),
.B(n_288),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1000),
.B(n_373),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_389),
.B1(n_387),
.B2(n_384),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_981),
.A2(n_389),
.B(n_387),
.C(n_384),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1022),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_892),
.B(n_373),
.Y(n_1150)
);

CKINVDCx8_ASAP7_75t_R g1151 ( 
.A(n_948),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1029),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1038),
.A2(n_1051),
.B(n_1028),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_936),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_936),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1029),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_990),
.B(n_374),
.Y(n_1158)
);

AO21x2_ASAP7_75t_L g1159 ( 
.A1(n_920),
.A2(n_242),
.B(n_348),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_955),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1035),
.A2(n_383),
.B1(n_380),
.B2(n_377),
.Y(n_1161)
);

INVx6_ASAP7_75t_L g1162 ( 
.A(n_939),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_1036),
.B1(n_1024),
.B2(n_993),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_942),
.B(n_374),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_904),
.A2(n_311),
.B(n_368),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1034),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1041),
.A2(n_1036),
.B1(n_992),
.B2(n_908),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_981),
.A2(n_377),
.B(n_356),
.C(n_308),
.Y(n_1168)
);

INVx3_ASAP7_75t_SL g1169 ( 
.A(n_964),
.Y(n_1169)
);

AND2x2_ASAP7_75t_SL g1170 ( 
.A(n_896),
.B(n_348),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_958),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_936),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1012),
.B(n_282),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1012),
.B(n_289),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_936),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_942),
.B(n_295),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1040),
.A2(n_323),
.B1(n_335),
.B2(n_331),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_915),
.A2(n_348),
.B(n_3),
.C(n_4),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_998),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_943),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_968),
.A2(n_328),
.B1(n_322),
.B2(n_303),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_893),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1033),
.A2(n_301),
.B(n_297),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1060),
.A2(n_193),
.B(n_180),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1056),
.A2(n_161),
.B(n_159),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_SL g1186 ( 
.A1(n_892),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_L g1187 ( 
.A1(n_969),
.A2(n_146),
.B(n_138),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_895),
.B(n_137),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_997),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.C(n_11),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1034),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_968),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_972),
.A2(n_15),
.B1(n_16),
.B2(n_22),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_924),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_949),
.B(n_132),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_950),
.B(n_23),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_972),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_943),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_937),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1047),
.A2(n_28),
.B(n_31),
.C(n_32),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_930),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_922),
.B(n_28),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_996),
.A2(n_120),
.B(n_114),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_938),
.A2(n_32),
.B(n_34),
.C(n_37),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_943),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_922),
.B(n_40),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_SL g1206 ( 
.A(n_906),
.B(n_41),
.C(n_42),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1006),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_943),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1055),
.B(n_46),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1049),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1004),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_L g1212 ( 
.A(n_905),
.B(n_48),
.C(n_52),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_956),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1081),
.A2(n_1047),
.B(n_1016),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1153),
.A2(n_1026),
.B(n_978),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1090),
.A2(n_928),
.B(n_918),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1098),
.A2(n_1056),
.A3(n_959),
.B(n_983),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1213),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1100),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1150),
.B(n_966),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1126),
.B(n_934),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1193),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_1153),
.A2(n_975),
.B(n_999),
.Y(n_1223)
);

AND2x6_ASAP7_75t_SL g1224 ( 
.A(n_1146),
.B(n_989),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1119),
.B(n_1008),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1066),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1089),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1065),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1211),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1076),
.B(n_949),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_1066),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1107),
.A2(n_919),
.B(n_931),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1069),
.Y(n_1233)
);

NAND2x1_ASAP7_75t_L g1234 ( 
.A(n_1180),
.B(n_1015),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1102),
.A2(n_999),
.B(n_970),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1106),
.Y(n_1236)
);

INVxp33_ASAP7_75t_SL g1237 ( 
.A(n_1088),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1083),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1078),
.B(n_1055),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1105),
.A2(n_913),
.B(n_898),
.C(n_1016),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1096),
.A2(n_1113),
.B(n_1121),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1066),
.Y(n_1242)
);

OAI21xp33_ASAP7_75t_L g1243 ( 
.A1(n_1105),
.A2(n_898),
.B(n_1008),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1143),
.B(n_986),
.Y(n_1244)
);

NOR4xp25_ASAP7_75t_L g1245 ( 
.A(n_1199),
.B(n_1007),
.C(n_1011),
.D(n_1002),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1180),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1068),
.A2(n_1050),
.B(n_946),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1075),
.B(n_1079),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1185),
.A2(n_988),
.B(n_1045),
.C(n_994),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1158),
.B(n_986),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1139),
.A2(n_931),
.B(n_1062),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1173),
.B(n_935),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1120),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1071),
.A2(n_1031),
.B(n_1030),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1197),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1079),
.B(n_994),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1154),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1085),
.B(n_1063),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1067),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1212),
.B(n_1037),
.C(n_1042),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1171),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1072),
.A2(n_1019),
.B(n_1044),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1201),
.B(n_923),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1122),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1211),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1096),
.A2(n_1048),
.B(n_1043),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1095),
.A2(n_1010),
.B(n_1059),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1125),
.A2(n_976),
.B(n_1003),
.Y(n_1268)
);

AND2x6_ASAP7_75t_SL g1269 ( 
.A(n_1195),
.B(n_989),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1080),
.A2(n_891),
.B1(n_907),
.B2(n_989),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1115),
.B(n_1063),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1093),
.B(n_1108),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1108),
.B(n_1058),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1169),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1109),
.B(n_1058),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1080),
.A2(n_1045),
.B(n_1052),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1109),
.B(n_1044),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1163),
.B(n_1054),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1211),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1185),
.A2(n_973),
.B(n_1054),
.C(n_58),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1130),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1137),
.A2(n_1054),
.B(n_75),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1148),
.A2(n_48),
.B(n_53),
.C(n_59),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1073),
.A2(n_1054),
.B(n_76),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1174),
.B(n_1087),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1170),
.B(n_53),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1167),
.A2(n_60),
.B(n_63),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1205),
.B(n_60),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1164),
.B(n_63),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1163),
.B(n_67),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_R g1291 ( 
.A(n_1151),
.B(n_71),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1209),
.B(n_82),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1133),
.A2(n_87),
.B(n_88),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1123),
.A2(n_1124),
.B(n_1101),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1099),
.A2(n_1086),
.B(n_1084),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1110),
.A2(n_1084),
.B(n_1141),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1188),
.A2(n_1116),
.B(n_1187),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1198),
.B(n_1074),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1132),
.Y(n_1300)
);

OAI22x1_ASAP7_75t_L g1301 ( 
.A1(n_1103),
.A2(n_1177),
.B1(n_1176),
.B2(n_1194),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1074),
.B(n_1110),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1138),
.A2(n_1160),
.B1(n_1140),
.B2(n_1144),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1162),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1092),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1182),
.B(n_1200),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1094),
.B(n_1197),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1114),
.Y(n_1308)
);

AOI211x1_ASAP7_75t_L g1309 ( 
.A1(n_1191),
.A2(n_1192),
.B(n_1196),
.C(n_1161),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1070),
.B(n_1097),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_SL g1311 ( 
.A(n_1186),
.B(n_1179),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1168),
.A2(n_1183),
.B(n_1189),
.C(n_1207),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_L g1313 ( 
.A1(n_1099),
.A2(n_1145),
.B(n_1104),
.C(n_1128),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1082),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1188),
.A2(n_1135),
.B(n_1202),
.Y(n_1315)
);

NAND3x1_ASAP7_75t_L g1316 ( 
.A(n_1077),
.B(n_1172),
.C(n_1091),
.Y(n_1316)
);

AOI21xp33_ASAP7_75t_L g1317 ( 
.A1(n_1147),
.A2(n_1133),
.B(n_1161),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1135),
.A2(n_1184),
.B(n_1134),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1077),
.B(n_1091),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1162),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1155),
.A2(n_1131),
.B1(n_1136),
.B2(n_1166),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1129),
.B(n_1210),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1142),
.A2(n_1157),
.B(n_1190),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1149),
.Y(n_1324)
);

OAI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1147),
.A2(n_1206),
.B(n_1111),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1152),
.B(n_1165),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1118),
.A2(n_1192),
.A3(n_1191),
.B(n_1196),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1181),
.B(n_1159),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1203),
.A2(n_1178),
.B(n_1127),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1082),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1156),
.A2(n_1181),
.B(n_1175),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1208),
.A2(n_1082),
.B(n_1175),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1204),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1150),
.A2(n_743),
.B1(n_405),
.B2(n_403),
.Y(n_1335)
);

AND2x6_ASAP7_75t_L g1336 ( 
.A(n_1075),
.B(n_1066),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1065),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1146),
.A2(n_1035),
.B1(n_1150),
.B2(n_932),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1105),
.B(n_795),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1211),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1193),
.Y(n_1341)
);

O2A1O1Ixp5_ASAP7_75t_SL g1342 ( 
.A1(n_1068),
.A2(n_1071),
.B(n_1105),
.C(n_1051),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1065),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1153),
.A2(n_1096),
.B(n_1102),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_SL g1345 ( 
.A1(n_1105),
.A2(n_1068),
.B(n_1185),
.C(n_1199),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1150),
.B(n_403),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1126),
.B(n_890),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1158),
.B(n_523),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1102),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1126),
.B(n_890),
.Y(n_1350)
);

NOR3xp33_ASAP7_75t_L g1351 ( 
.A(n_1150),
.B(n_743),
.C(n_695),
.Y(n_1351)
);

NAND2x1_ASAP7_75t_L g1352 ( 
.A(n_1180),
.B(n_987),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1193),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1193),
.Y(n_1354)
);

AOI21xp33_ASAP7_75t_L g1355 ( 
.A1(n_1081),
.A2(n_743),
.B(n_805),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1117),
.A2(n_1090),
.B(n_1107),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1126),
.B(n_890),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1309),
.B(n_1276),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1339),
.A2(n_1335),
.B1(n_1311),
.B2(n_1258),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1323),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1355),
.B(n_1351),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1319),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1346),
.A2(n_1339),
.B1(n_1310),
.B2(n_1301),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1248),
.B(n_1278),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1349),
.A2(n_1296),
.B(n_1297),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1218),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1319),
.B(n_1230),
.Y(n_1368)
);

AOI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1243),
.A2(n_1317),
.B(n_1328),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1219),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1341),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1357),
.B(n_1272),
.Y(n_1373)
);

AOI221xp5_ASAP7_75t_L g1374 ( 
.A1(n_1345),
.A2(n_1288),
.B1(n_1289),
.B2(n_1338),
.C(n_1283),
.Y(n_1374)
);

INVxp33_ASAP7_75t_SL g1375 ( 
.A(n_1220),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1349),
.A2(n_1296),
.B(n_1298),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1228),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1325),
.B(n_1280),
.C(n_1243),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1233),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1307),
.B(n_1302),
.Y(n_1380)
);

NAND2x1_ASAP7_75t_L g1381 ( 
.A(n_1336),
.B(n_1246),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1315),
.A2(n_1260),
.B(n_1235),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1282),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1253),
.B(n_1257),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1226),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1316),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1260),
.A2(n_1235),
.B(n_1216),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1287),
.A2(n_1293),
.B1(n_1325),
.B2(n_1286),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1294),
.Y(n_1390)
);

OAI221xp5_ASAP7_75t_L g1391 ( 
.A1(n_1348),
.A2(n_1293),
.B1(n_1285),
.B2(n_1311),
.C(n_1313),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1214),
.A2(n_1342),
.B(n_1275),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1331),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1236),
.Y(n_1394)
);

CKINVDCx6p67_ASAP7_75t_R g1395 ( 
.A(n_1274),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1318),
.A2(n_1268),
.B(n_1232),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1324),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1240),
.B(n_1225),
.C(n_1290),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1222),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1226),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1264),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1267),
.A2(n_1247),
.B(n_1284),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1261),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1267),
.A2(n_1266),
.B(n_1262),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1353),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1266),
.A2(n_1270),
.B(n_1276),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1237),
.A2(n_1244),
.B(n_1250),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1270),
.A2(n_1254),
.B(n_1241),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1307),
.B(n_1336),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1263),
.A2(n_1273),
.B1(n_1252),
.B2(n_1353),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1241),
.A2(n_1344),
.B(n_1326),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1281),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1321),
.A2(n_1329),
.B(n_1277),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1249),
.A2(n_1292),
.B(n_1256),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1226),
.B(n_1242),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1303),
.A2(n_1332),
.B(n_1305),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1303),
.A2(n_1306),
.B(n_1300),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1354),
.A2(n_1227),
.B1(n_1299),
.B2(n_1271),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1322),
.A2(n_1234),
.B(n_1308),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1259),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1352),
.A2(n_1343),
.B(n_1337),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1217),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1333),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1299),
.A2(n_1265),
.B1(n_1304),
.B2(n_1242),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1246),
.A2(n_1255),
.B(n_1330),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1336),
.B(n_1334),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1217),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1255),
.A2(n_1330),
.B(n_1334),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1217),
.A2(n_1245),
.B(n_1215),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1215),
.A2(n_1223),
.B(n_1327),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1333),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1223),
.A2(n_1327),
.B(n_1269),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1291),
.A2(n_1259),
.B1(n_1224),
.B2(n_1320),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1231),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1229),
.Y(n_1435)
);

AND2x6_ASAP7_75t_L g1436 ( 
.A(n_1229),
.B(n_1279),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1314),
.B(n_1340),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1327),
.A2(n_1269),
.B(n_1224),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1231),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1231),
.A2(n_1242),
.B1(n_1229),
.B2(n_1279),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1279),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1340),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1340),
.B(n_1221),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1218),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1341),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1319),
.B(n_1230),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1341),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1335),
.A2(n_1351),
.B1(n_1258),
.B2(n_1346),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1341),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1351),
.A2(n_1355),
.B(n_1317),
.C(n_1280),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1218),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1226),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1456)
);

INVx3_ASAP7_75t_SL g1457 ( 
.A(n_1274),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1458)
);

NAND2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1226),
.B(n_1231),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1221),
.B(n_1126),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1339),
.A2(n_1335),
.B1(n_1311),
.B2(n_620),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1218),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1335),
.A2(n_1351),
.B1(n_1258),
.B2(n_1346),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_SL g1465 ( 
.A1(n_1287),
.A2(n_1185),
.B(n_1239),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1341),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1355),
.B(n_1346),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1323),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1335),
.A2(n_1351),
.B1(n_1258),
.B2(n_1346),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1226),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1323),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1351),
.A2(n_1317),
.B1(n_1105),
.B2(n_1339),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1339),
.A2(n_1335),
.B1(n_1311),
.B2(n_620),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1218),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1265),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1265),
.Y(n_1486)
);

INVxp33_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1319),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1323),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_1335),
.B2(n_743),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1218),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1355),
.B(n_1346),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1221),
.B(n_1126),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1218),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1319),
.B(n_1230),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1339),
.A2(n_1335),
.B1(n_1311),
.B2(n_620),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_SL g1500 ( 
.A1(n_1317),
.A2(n_1280),
.B(n_1312),
.C(n_1105),
.Y(n_1500)
);

AOI211xp5_ASAP7_75t_L g1501 ( 
.A1(n_1351),
.A2(n_1355),
.B(n_620),
.C(n_743),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1218),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1253),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1319),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1356),
.A2(n_1295),
.B(n_1251),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1335),
.A2(n_1351),
.B1(n_1258),
.B2(n_1346),
.Y(n_1506)
);

OA22x2_ASAP7_75t_L g1507 ( 
.A1(n_1364),
.A2(n_1490),
.B1(n_1407),
.B2(n_1506),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1450),
.A2(n_1494),
.B(n_1467),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1426),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1367),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1460),
.B(n_1496),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1467),
.A2(n_1494),
.B1(n_1501),
.B2(n_1480),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1362),
.A2(n_1463),
.B(n_1448),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1362),
.A2(n_1461),
.B(n_1499),
.C(n_1474),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1370),
.Y(n_1516)
);

O2A1O1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1360),
.A2(n_1500),
.B(n_1374),
.C(n_1391),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1429),
.A2(n_1392),
.B(n_1408),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1432),
.B(n_1438),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1426),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1405),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1443),
.B(n_1452),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1409),
.B(n_1380),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1415),
.A2(n_1459),
.B(n_1434),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1389),
.A2(n_1378),
.B1(n_1479),
.B2(n_1398),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1493),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1389),
.A2(n_1479),
.B1(n_1433),
.B2(n_1464),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1432),
.B(n_1438),
.Y(n_1528)
);

NAND2xp33_ASAP7_75t_SL g1529 ( 
.A(n_1434),
.B(n_1381),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1500),
.A2(n_1369),
.B(n_1465),
.C(n_1410),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1394),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1380),
.Y(n_1532)
);

AND2x4_ASAP7_75t_SL g1533 ( 
.A(n_1409),
.B(n_1371),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1415),
.A2(n_1459),
.B(n_1434),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1487),
.A2(n_1375),
.B1(n_1418),
.B2(n_1359),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1380),
.B(n_1368),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1368),
.B(n_1446),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1368),
.B(n_1446),
.Y(n_1538)
);

O2A1O1Ixp5_ASAP7_75t_L g1539 ( 
.A1(n_1393),
.A2(n_1383),
.B(n_1427),
.C(n_1424),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1446),
.B(n_1498),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1395),
.Y(n_1541)
);

O2A1O1Ixp5_ASAP7_75t_L g1542 ( 
.A1(n_1387),
.A2(n_1439),
.B(n_1431),
.C(n_1361),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1416),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_1399),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1445),
.B(n_1447),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1375),
.A2(n_1359),
.B1(n_1466),
.B2(n_1503),
.Y(n_1546)
);

AOI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1457),
.A2(n_1384),
.B(n_1449),
.C(n_1403),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1498),
.B(n_1363),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_R g1549 ( 
.A(n_1442),
.B(n_1420),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1442),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1434),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1395),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1417),
.A2(n_1359),
.B(n_1401),
.C(n_1497),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1475),
.A2(n_1440),
.B(n_1414),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1412),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1485),
.A2(n_1486),
.B1(n_1453),
.B2(n_1462),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1444),
.A2(n_1491),
.B1(n_1502),
.B2(n_1484),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1475),
.A2(n_1414),
.B(n_1400),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1437),
.B(n_1379),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1379),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1386),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1402),
.A2(n_1396),
.B(n_1411),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1365),
.B(n_1397),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1435),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1386),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1475),
.A2(n_1414),
.B(n_1454),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1396),
.A2(n_1411),
.B(n_1404),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1390),
.B(n_1397),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1404),
.A2(n_1406),
.B(n_1413),
.Y(n_1571)
);

CKINVDCx16_ASAP7_75t_R g1572 ( 
.A(n_1436),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1365),
.Y(n_1573)
);

O2A1O1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1488),
.A2(n_1504),
.B(n_1366),
.C(n_1454),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1423),
.A2(n_1419),
.B(n_1366),
.C(n_1421),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1504),
.A2(n_1400),
.B(n_1385),
.C(n_1376),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1365),
.B(n_1441),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1441),
.B(n_1436),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1385),
.B(n_1428),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1430),
.B(n_1376),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1423),
.B(n_1428),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1430),
.B(n_1382),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1430),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1421),
.B(n_1425),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1419),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1425),
.B(n_1436),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1471),
.A2(n_1489),
.B(n_1478),
.C(n_1382),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1388),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1358),
.B(n_1473),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1451),
.B(n_1455),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1456),
.A2(n_1458),
.B(n_1468),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1458),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1470),
.B(n_1472),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1481),
.A2(n_1482),
.B1(n_1483),
.B2(n_1492),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1481),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1495),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1495),
.B(n_1505),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1505),
.B(n_1460),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1362),
.A2(n_1351),
.B(n_1355),
.C(n_1501),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1450),
.A2(n_1293),
.B(n_1105),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1362),
.A2(n_1351),
.B(n_1355),
.C(n_1501),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1422),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1450),
.A2(n_1293),
.B(n_1105),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1367),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1422),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1422),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1490),
.A2(n_1364),
.B1(n_1335),
.B2(n_1467),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1490),
.A2(n_1364),
.B1(n_1335),
.B2(n_1467),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1490),
.A2(n_1364),
.B1(n_1335),
.B2(n_1467),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1450),
.A2(n_1293),
.B(n_1105),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1467),
.B(n_1494),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1429),
.A2(n_1392),
.B(n_1408),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1460),
.B(n_1496),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1460),
.B(n_1496),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1362),
.A2(n_1351),
.B(n_1355),
.C(n_1501),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1460),
.B(n_1496),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1600),
.B(n_1518),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1573),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1616),
.A2(n_1614),
.B1(n_1612),
.B2(n_1613),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1616),
.A2(n_1525),
.B1(n_1513),
.B2(n_1508),
.Y(n_1627)
);

INVxp33_ASAP7_75t_L g1628 ( 
.A(n_1549),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1514),
.A2(n_1604),
.B(n_1601),
.Y(n_1629)
);

NOR2x1_ASAP7_75t_L g1630 ( 
.A(n_1560),
.B(n_1568),
.Y(n_1630)
);

AND2x4_ASAP7_75t_SL g1631 ( 
.A(n_1581),
.B(n_1586),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1581),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1569),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1558),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1518),
.B(n_1617),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1533),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1617),
.B(n_1580),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1519),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1519),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1507),
.A2(n_1527),
.B1(n_1535),
.B2(n_1515),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1519),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1642)
);

AOI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1591),
.A2(n_1596),
.B(n_1599),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1620),
.A2(n_1517),
.B1(n_1606),
.B2(n_1615),
.C(n_1603),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1526),
.B(n_1512),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1605),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1528),
.B(n_1609),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1609),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1507),
.A2(n_1602),
.B1(n_1608),
.B2(n_1610),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1510),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1585),
.B(n_1579),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1516),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1531),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1528),
.B(n_1583),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1528),
.B(n_1543),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1530),
.A2(n_1522),
.B(n_1511),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1569),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1533),
.Y(n_1660)
);

BUFx4f_ASAP7_75t_SL g1661 ( 
.A(n_1566),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1523),
.Y(n_1662)
);

BUFx8_ASAP7_75t_SL g1663 ( 
.A(n_1541),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1556),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1607),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1550),
.B(n_1559),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1562),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1569),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1564),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1555),
.B(n_1574),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1564),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1575),
.B(n_1589),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1544),
.B(n_1565),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1563),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1549),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1572),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1590),
.Y(n_1677)
);

AO21x2_ASAP7_75t_L g1678 ( 
.A1(n_1592),
.A2(n_1597),
.B(n_1598),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1598),
.B(n_1595),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1532),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1567),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1587),
.B(n_1536),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1523),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1546),
.B(n_1521),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1642),
.B(n_1557),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1642),
.B(n_1622),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1623),
.B(n_1576),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1623),
.B(n_1539),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1654),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1623),
.B(n_1577),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1666),
.B(n_1554),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1657),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1524),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1655),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1570),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1664),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1682),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1652),
.B(n_1547),
.Y(n_1704)
);

INVx2_ASAP7_75t_R g1705 ( 
.A(n_1635),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1682),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1636),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1681),
.B(n_1548),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1631),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1625),
.A2(n_1551),
.B(n_1540),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1627),
.A2(n_1538),
.B1(n_1537),
.B2(n_1566),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1681),
.B(n_1637),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1656),
.B(n_1645),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_1645),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1638),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1679),
.B(n_1542),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1625),
.A2(n_1553),
.B1(n_1509),
.B2(n_1520),
.Y(n_1718)
);

INVx3_ASAP7_75t_SL g1719 ( 
.A(n_1670),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1678),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1671),
.B(n_1669),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1695),
.B(n_1629),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1710),
.A2(n_1629),
.B(n_1640),
.C(n_1651),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1718),
.A2(n_1640),
.B1(n_1651),
.B2(n_1644),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1716),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1695),
.A2(n_1627),
.B(n_1644),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1711),
.A2(n_1710),
.B1(n_1704),
.B2(n_1697),
.Y(n_1728)
);

OAI31xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1690),
.A2(n_1630),
.A3(n_1658),
.B(n_1672),
.Y(n_1729)
);

AOI31xp33_ASAP7_75t_L g1730 ( 
.A1(n_1704),
.A2(n_1628),
.A3(n_1630),
.B(n_1658),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1690),
.A2(n_1634),
.B1(n_1652),
.B2(n_1646),
.C(n_1683),
.Y(n_1731)
);

INVx4_ASAP7_75t_L g1732 ( 
.A(n_1697),
.Y(n_1732)
);

OAI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1711),
.A2(n_1634),
.B(n_1686),
.C(n_1646),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1716),
.B(n_1632),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1707),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1670),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1714),
.A2(n_1643),
.B(n_1659),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1699),
.B(n_1673),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1718),
.A2(n_1686),
.B(n_1673),
.C(n_1684),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1690),
.A2(n_1683),
.B1(n_1686),
.B2(n_1680),
.C(n_1653),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1626),
.Y(n_1742)
);

AOI222xp33_ASAP7_75t_L g1743 ( 
.A1(n_1692),
.A2(n_1661),
.B1(n_1683),
.B2(n_1680),
.C1(n_1676),
.C2(n_1675),
.Y(n_1743)
);

OAI33xp33_ASAP7_75t_L g1744 ( 
.A1(n_1687),
.A2(n_1691),
.A3(n_1693),
.B1(n_1698),
.B2(n_1702),
.B3(n_1701),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1697),
.A2(n_1676),
.B1(n_1670),
.B2(n_1624),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1706),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1697),
.A2(n_1676),
.B1(n_1670),
.B2(n_1624),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1707),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1712),
.B(n_1632),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1716),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1699),
.B(n_1684),
.Y(n_1751)
);

OAI31xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1692),
.A2(n_1672),
.A3(n_1624),
.B(n_1653),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1712),
.B(n_1677),
.Y(n_1753)
);

INVx4_ASAP7_75t_L g1754 ( 
.A(n_1697),
.Y(n_1754)
);

OAI33xp33_ASAP7_75t_L g1755 ( 
.A1(n_1687),
.A2(n_1667),
.A3(n_1674),
.B1(n_1650),
.B2(n_1647),
.B3(n_1649),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1688),
.Y(n_1756)
);

OAI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1692),
.A2(n_1639),
.B(n_1641),
.C(n_1676),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1694),
.B(n_1677),
.Y(n_1758)
);

OAI211xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1687),
.A2(n_1648),
.B(n_1667),
.C(n_1578),
.Y(n_1759)
);

OAI21xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1709),
.A2(n_1670),
.B(n_1685),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1697),
.A2(n_1624),
.B1(n_1685),
.B2(n_1662),
.Y(n_1761)
);

AND2x6_ASAP7_75t_L g1762 ( 
.A(n_1753),
.B(n_1662),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1726),
.A2(n_1660),
.B(n_1636),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1727),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1727),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1721),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1750),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1737),
.A2(n_1643),
.B(n_1633),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1729),
.B(n_1661),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1753),
.B(n_1705),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1721),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1750),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1721),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1724),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1746),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1728),
.B(n_1719),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1743),
.B(n_1719),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1721),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1731),
.B(n_1717),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1717),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1705),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1705),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1741),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1752),
.B(n_1719),
.Y(n_1786)
);

INVx4_ASAP7_75t_SL g1787 ( 
.A(n_1736),
.Y(n_1787)
);

NOR2x1p5_ASAP7_75t_L g1788 ( 
.A(n_1732),
.B(n_1707),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1736),
.B(n_1709),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1732),
.B(n_1696),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1736),
.Y(n_1791)
);

INVx5_ASAP7_75t_L g1792 ( 
.A(n_1732),
.Y(n_1792)
);

NOR2xp67_ASAP7_75t_L g1793 ( 
.A(n_1786),
.B(n_1757),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1781),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1767),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1763),
.B(n_1740),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1788),
.B(n_1787),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1773),
.Y(n_1798)
);

NOR2xp67_ASAP7_75t_L g1799 ( 
.A(n_1786),
.B(n_1760),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1781),
.B(n_1730),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1768),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1770),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1770),
.B(n_1738),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1788),
.B(n_1742),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1767),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1787),
.B(n_1742),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1787),
.B(n_1749),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1787),
.B(n_1792),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1773),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1776),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1776),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1787),
.B(n_1725),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1767),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1792),
.B(n_1754),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1765),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1775),
.B(n_1723),
.C(n_1733),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1775),
.B(n_1694),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.B(n_1725),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1790),
.B(n_1754),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1765),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1735),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1778),
.A2(n_1760),
.B(n_1739),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1778),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1694),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1782),
.B(n_1713),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1790),
.B(n_1735),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1766),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1762),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1768),
.B(n_1715),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1777),
.A2(n_1759),
.B(n_1745),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1790),
.B(n_1748),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1779),
.B(n_1751),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1789),
.B(n_1748),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1777),
.A2(n_1719),
.B1(n_1747),
.B2(n_1755),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1734),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1779),
.B(n_1688),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1764),
.B(n_1789),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1816),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1809),
.B(n_1792),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_L g1841 ( 
.A(n_1817),
.B(n_1744),
.C(n_1769),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1801),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1817),
.B(n_1708),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1824),
.A2(n_1761),
.B1(n_1791),
.B2(n_1779),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1833),
.B(n_1689),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1805),
.B(n_1822),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1837),
.B(n_1689),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1816),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1821),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1798),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1821),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1828),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1818),
.B(n_1689),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1824),
.B(n_1700),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1804),
.B(n_1700),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1828),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1797),
.Y(n_1857)
);

INVxp33_ASAP7_75t_L g1858 ( 
.A(n_1793),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1809),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1795),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1800),
.B(n_1708),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1811),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1811),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1812),
.Y(n_1864)
);

AND2x4_ASAP7_75t_SL g1865 ( 
.A(n_1797),
.B(n_1789),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1794),
.B(n_1700),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1812),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1798),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1802),
.B(n_1796),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1810),
.B(n_1793),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1835),
.A2(n_1784),
.B(n_1783),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1810),
.B(n_1835),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1838),
.B(n_1779),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1830),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1795),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1850),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1850),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1870),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1839),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1805),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1868),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1842),
.B(n_1830),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1858),
.B(n_1823),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1857),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1865),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1840),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1846),
.B(n_1838),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1871),
.A2(n_1872),
.B(n_1841),
.Y(n_1888)
);

NAND2x1_ASAP7_75t_L g1889 ( 
.A(n_1873),
.B(n_1838),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1869),
.A2(n_1838),
.B(n_1831),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1859),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1841),
.A2(n_1799),
.B1(n_1838),
.B2(n_1831),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1843),
.B(n_1822),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1865),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1848),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1859),
.B(n_1809),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1849),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1851),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1852),
.Y(n_1899)
);

AO21x2_ASAP7_75t_L g1900 ( 
.A1(n_1873),
.A2(n_1799),
.B(n_1809),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1861),
.B(n_1663),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1856),
.Y(n_1902)
);

OAI21xp33_ASAP7_75t_L g1903 ( 
.A1(n_1892),
.A2(n_1844),
.B(n_1874),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1883),
.A2(n_1863),
.B(n_1862),
.Y(n_1904)
);

INVxp33_ASAP7_75t_L g1905 ( 
.A(n_1888),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1885),
.Y(n_1906)
);

INVxp67_ASAP7_75t_SL g1907 ( 
.A(n_1891),
.Y(n_1907)
);

OAI31xp33_ASAP7_75t_L g1908 ( 
.A1(n_1890),
.A2(n_1840),
.A3(n_1803),
.B(n_1813),
.Y(n_1908)
);

AOI33xp33_ASAP7_75t_L g1909 ( 
.A1(n_1878),
.A2(n_1867),
.A3(n_1864),
.B1(n_1803),
.B2(n_1815),
.B3(n_1813),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1884),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1876),
.A2(n_1803),
.B1(n_1854),
.B2(n_1815),
.C(n_1834),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1894),
.B(n_1827),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1888),
.A2(n_1853),
.B1(n_1829),
.B2(n_1803),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1896),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1888),
.A2(n_1791),
.B1(n_1829),
.B2(n_1855),
.C(n_1834),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1881),
.B(n_1866),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1877),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1877),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1894),
.A2(n_1829),
.B1(n_1807),
.B2(n_1789),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1880),
.B(n_1881),
.C(n_1882),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1882),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1893),
.B(n_1845),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1896),
.B(n_1827),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1912),
.B(n_1887),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1906),
.B(n_1887),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1920),
.B(n_1900),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1921),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1910),
.B(n_1900),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1905),
.B(n_1879),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1914),
.B(n_1901),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1905),
.B(n_1901),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1907),
.B(n_1896),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1921),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1908),
.B(n_1913),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1917),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1926),
.A2(n_1904),
.B(n_1903),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1927),
.A2(n_1918),
.B(n_1915),
.C(n_1900),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1931),
.A2(n_1911),
.B(n_1916),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1933),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1927),
.A2(n_1931),
.B1(n_1934),
.B2(n_1928),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1929),
.A2(n_1889),
.B(n_1923),
.Y(n_1941)
);

NAND4xp75_ASAP7_75t_L g1942 ( 
.A(n_1925),
.B(n_1929),
.C(n_1930),
.D(n_1935),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1932),
.Y(n_1943)
);

OAI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1924),
.A2(n_1886),
.B(n_1898),
.C(n_1902),
.Y(n_1944)
);

NOR3xp33_ASAP7_75t_L g1945 ( 
.A(n_1932),
.B(n_1909),
.C(n_1919),
.Y(n_1945)
);

OAI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1926),
.A2(n_1922),
.B1(n_1886),
.B2(n_1899),
.C(n_1897),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_R g1947 ( 
.A(n_1943),
.B(n_1939),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1946),
.Y(n_1948)
);

NAND4xp25_ASAP7_75t_L g1949 ( 
.A(n_1945),
.B(n_1936),
.C(n_1938),
.D(n_1941),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1886),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1944),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1940),
.A2(n_1815),
.B1(n_1829),
.B2(n_1895),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1937),
.A2(n_1815),
.B1(n_1832),
.B2(n_1820),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1950),
.Y(n_1954)
);

NAND2x1p5_ASAP7_75t_L g1955 ( 
.A(n_1951),
.B(n_1792),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1947),
.B(n_1948),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1953),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1949),
.B(n_1909),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1952),
.A2(n_1791),
.B1(n_1860),
.B2(n_1875),
.C(n_1792),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1950),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1947),
.Y(n_1961)
);

NOR3xp33_ASAP7_75t_L g1962 ( 
.A(n_1949),
.B(n_1875),
.C(n_1860),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1954),
.A2(n_1960),
.B(n_1958),
.C(n_1956),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1961),
.A2(n_1807),
.B(n_1808),
.Y(n_1964)
);

INVxp67_ASAP7_75t_SL g1965 ( 
.A(n_1955),
.Y(n_1965)
);

OAI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1960),
.A2(n_1791),
.B1(n_1792),
.B2(n_1820),
.C(n_1808),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_R g1967 ( 
.A(n_1957),
.B(n_1832),
.Y(n_1967)
);

NOR2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1965),
.B(n_1967),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1963),
.B(n_1962),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1964),
.B(n_1836),
.Y(n_1970)
);

AND3x1_ASAP7_75t_L g1971 ( 
.A(n_1968),
.B(n_1966),
.C(n_1959),
.Y(n_1971)
);

AOI322xp5_ASAP7_75t_L g1972 ( 
.A1(n_1971),
.A2(n_1970),
.A3(n_1969),
.B1(n_1795),
.B2(n_1814),
.C1(n_1806),
.C2(n_1819),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1972),
.Y(n_1973)
);

AOI21xp33_ASAP7_75t_L g1974 ( 
.A1(n_1972),
.A2(n_1814),
.B(n_1806),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_R g1975 ( 
.A(n_1973),
.B(n_1529),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1974),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1976),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1975),
.A2(n_1806),
.B1(n_1814),
.B2(n_1847),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1977),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_SL g1980 ( 
.A1(n_1979),
.A2(n_1978),
.B1(n_1819),
.B2(n_1792),
.Y(n_1980)
);

OA21x2_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1836),
.B(n_1825),
.Y(n_1981)
);

AOI322xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1792),
.A3(n_1772),
.B1(n_1767),
.B2(n_1774),
.C1(n_1780),
.C2(n_1771),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1826),
.B1(n_1772),
.B2(n_1785),
.Y(n_1983)
);

AOI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1534),
.B(n_1552),
.C(n_1529),
.Y(n_1984)
);


endmodule