module fake_ibex_656_n_2238 (n_151, n_85, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2238);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2238;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_399;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2162;
wire n_2236;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_1845;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_634;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_2186;
wire n_1843;
wire n_408;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_75),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_380),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_262),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_341),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_327),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_50),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_383),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_211),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_293),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_52),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_329),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_35),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_128),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_50),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_154),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_26),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_225),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_55),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_99),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_260),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_199),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_218),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_82),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_39),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_143),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_198),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_18),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_22),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_190),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_298),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_203),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_59),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_368),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_294),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_213),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_94),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_253),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_13),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_181),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_255),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_301),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_226),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_207),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_337),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_102),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_348),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_222),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_338),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_384),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_161),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_243),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_4),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_79),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_74),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_221),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_264),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_263),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_144),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_192),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_36),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_112),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_6),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_322),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_68),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_355),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_357),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_58),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_111),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_93),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_214),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_179),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_373),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_113),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_382),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_129),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_124),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_200),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_155),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_208),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_147),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_31),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_38),
.B(n_167),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_149),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_18),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_331),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_185),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_111),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_284),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_271),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_306),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_112),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_114),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_171),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_360),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_372),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_165),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_283),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_178),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_45),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_379),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_130),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_210),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_321),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_101),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_59),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_351),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_250),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_41),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_105),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_52),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_46),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_246),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_184),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_41),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_267),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_167),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_202),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_138),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_147),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_290),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_350),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_242),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_82),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_305),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_282),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_312),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_376),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_15),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_323),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_6),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_236),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_71),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_102),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_299),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_216),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_239),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_251),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_224),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_385),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_371),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_220),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_139),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_60),
.Y(n_543)
);

BUFx5_ASAP7_75t_L g544 ( 
.A(n_195),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_187),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_76),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_97),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_24),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_269),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_340),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_30),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_36),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_191),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_296),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_209),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_391),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_5),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_95),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_69),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_86),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_188),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_74),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_285),
.Y(n_563)
);

BUFx5_ASAP7_75t_L g564 ( 
.A(n_21),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_40),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_104),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_288),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_34),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_83),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_42),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_153),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_204),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_313),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_324),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_238),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_79),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_149),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_244),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_108),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_138),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_20),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_48),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_325),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_261),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_157),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_361),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_336),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_70),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_223),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_170),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_292),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_212),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_374),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_153),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_63),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_150),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_387),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_302),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_109),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_31),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_57),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_139),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_115),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_8),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_205),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_227),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_23),
.B(n_85),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_256),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_47),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_314),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_215),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_175),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_10),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_258),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_162),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_83),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_289),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_354),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_186),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_286),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_133),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_310),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_127),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_87),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_123),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_266),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_352),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_131),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_362),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_78),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_363),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_72),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_182),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_134),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_142),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_265),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_86),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_343),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_233),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_295),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_231),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_119),
.B(n_104),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_150),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_280),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_196),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_28),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_57),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_389),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_228),
.Y(n_649)
);

INVxp33_ASAP7_75t_R g650 ( 
.A(n_3),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_330),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_365),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_364),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_308),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_22),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_359),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_157),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_377),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_259),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_339),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_8),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_100),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_206),
.B(n_134),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_106),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_21),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_105),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_194),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_148),
.Y(n_668)
);

BUFx8_ASAP7_75t_SL g669 ( 
.A(n_168),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_229),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_309),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_159),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_406),
.B(n_0),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_511),
.B(n_1),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_548),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_417),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_406),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_433),
.B(n_1),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_431),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_440),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_433),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_547),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_682)
);

BUFx8_ASAP7_75t_L g683 ( 
.A(n_564),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_481),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_453),
.A2(n_492),
.B1(n_659),
.B2(n_513),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_447),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_647),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_393),
.A2(n_173),
.B(n_172),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_417),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_SL g690 ( 
.A1(n_401),
.A2(n_559),
.B1(n_590),
.B2(n_557),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_564),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_481),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_403),
.Y(n_693)
);

AOI22x1_ASAP7_75t_SL g694 ( 
.A1(n_401),
.A2(n_7),
.B1(n_2),
.B2(n_5),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_481),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_473),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_464),
.B(n_575),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_485),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_481),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_506),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_564),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_393),
.A2(n_176),
.B(n_174),
.Y(n_703)
);

BUFx12f_ASAP7_75t_L g704 ( 
.A(n_403),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_403),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_397),
.B(n_7),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_669),
.Y(n_707)
);

BUFx12f_ASAP7_75t_L g708 ( 
.A(n_552),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_552),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_661),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_396),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_564),
.Y(n_713)
);

OA21x2_ASAP7_75t_L g714 ( 
.A1(n_427),
.A2(n_180),
.B(n_177),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_661),
.B(n_9),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_506),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_464),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_669),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_462),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_506),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_462),
.B(n_9),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_476),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_575),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_628),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_664),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_504),
.B(n_10),
.Y(n_727)
);

CKINVDCx6p67_ASAP7_75t_R g728 ( 
.A(n_610),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_564),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_549),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_576),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_579),
.B(n_11),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_12),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_544),
.B(n_12),
.Y(n_735)
);

BUFx12f_ASAP7_75t_L g736 ( 
.A(n_409),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_610),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_466),
.B(n_474),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_549),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_564),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_616),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_561),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_616),
.B(n_13),
.Y(n_744)
);

INVxp33_ASAP7_75t_SL g745 ( 
.A(n_392),
.Y(n_745)
);

CKINVDCx11_ASAP7_75t_R g746 ( 
.A(n_557),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_561),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_14),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_616),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_561),
.Y(n_750)
);

BUFx12f_ASAP7_75t_L g751 ( 
.A(n_578),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_528),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_606),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_402),
.Y(n_754)
);

XOR2xp5_ASAP7_75t_L g755 ( 
.A(n_559),
.B(n_14),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_639),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_561),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_489),
.B(n_605),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_584),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_603),
.B(n_16),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_590),
.Y(n_762)
);

OA21x2_ASAP7_75t_L g763 ( 
.A1(n_614),
.A2(n_189),
.B(n_183),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_616),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_480),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_616),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_614),
.B(n_17),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_584),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_395),
.B(n_19),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_584),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_404),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_616),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_673),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_673),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_679),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_708),
.B(n_399),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_673),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_R g779 ( 
.A(n_707),
.B(n_428),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_676),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_R g781 ( 
.A(n_718),
.B(n_428),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_708),
.B(n_400),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_686),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_721),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_684),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_698),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_721),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_762),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_709),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_709),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_705),
.B(n_487),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_693),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_693),
.Y(n_794)
);

BUFx6f_ASAP7_75t_SL g795 ( 
.A(n_678),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_691),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_727),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_745),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_733),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_R g801 ( 
.A(n_704),
.B(n_701),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_746),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_733),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_746),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_762),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_748),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_687),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_772),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_772),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_704),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_678),
.B(n_663),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_711),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_705),
.B(n_419),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_748),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_711),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_754),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_R g817 ( 
.A(n_701),
.B(n_487),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_703),
.A2(n_439),
.B(n_436),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_748),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_754),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_702),
.Y(n_821)
);

CKINVDCx16_ASAP7_75t_R g822 ( 
.A(n_685),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_702),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_675),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_728),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_736),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_683),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_760),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_726),
.B(n_460),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_736),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_725),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_705),
.B(n_539),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_690),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_688),
.A2(n_455),
.B(n_449),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_751),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_683),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_767),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_751),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_767),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_755),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_767),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_726),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_696),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_696),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_674),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_713),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_732),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_694),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_682),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_697),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_R g852 ( 
.A(n_680),
.B(n_539),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_732),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_676),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_753),
.Y(n_855)
);

AOI21x1_ASAP7_75t_L g856 ( 
.A1(n_766),
.A2(n_475),
.B(n_461),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_753),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_756),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_756),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_752),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_697),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_738),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_689),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_689),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_715),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_717),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_715),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_677),
.B(n_477),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_717),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_765),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_723),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_723),
.Y(n_873)
);

INVx8_ASAP7_75t_L g874 ( 
.A(n_697),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_734),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_744),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_681),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_SL g879 ( 
.A(n_735),
.B(n_398),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_737),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_737),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_706),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_729),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_735),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_706),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_758),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_740),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_758),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_719),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_769),
.A2(n_501),
.B(n_493),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_769),
.B(n_512),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_722),
.A2(n_599),
.B1(n_609),
.B2(n_595),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_731),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_740),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_741),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_758),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_742),
.B(n_416),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_758),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_741),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_R g900 ( 
.A(n_697),
.B(n_394),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_697),
.Y(n_901)
);

CKINVDCx16_ASAP7_75t_R g902 ( 
.A(n_749),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_764),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_688),
.Y(n_904)
);

INVxp33_ASAP7_75t_SL g905 ( 
.A(n_773),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_730),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_688),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_684),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_730),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_730),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_730),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_714),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_761),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_761),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_761),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_684),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_714),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_684),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_692),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_692),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_692),
.B(n_394),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_692),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_695),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_714),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_695),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_695),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_763),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_695),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_699),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_699),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_699),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_699),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_700),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_700),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_700),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_712),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_712),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_712),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_716),
.B(n_517),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_716),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_716),
.B(n_544),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_716),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_720),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_720),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_780),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_854),
.Y(n_946)
);

BUFx6f_ASAP7_75t_SL g947 ( 
.A(n_848),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_875),
.B(n_553),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_876),
.B(n_890),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_902),
.B(n_405),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_889),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_874),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_890),
.B(n_862),
.Y(n_953)
);

AND2x6_ASAP7_75t_SL g954 ( 
.A(n_788),
.B(n_650),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_789),
.B(n_23),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_812),
.B(n_457),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_815),
.B(n_469),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_844),
.B(n_421),
.C(n_420),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_863),
.B(n_407),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_774),
.B(n_626),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_806),
.Y(n_961)
);

AND2x4_ASAP7_75t_SL g962 ( 
.A(n_837),
.B(n_398),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_845),
.B(n_425),
.C(n_422),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_874),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_867),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_866),
.B(n_869),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_775),
.B(n_778),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_892),
.B(n_508),
.C(n_632),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_806),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_819),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_822),
.B(n_832),
.C(n_879),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_830),
.B(n_429),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_874),
.B(n_430),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_L g974 ( 
.A(n_811),
.B(n_544),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_891),
.B(n_520),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_843),
.B(n_443),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_828),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_872),
.B(n_873),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_877),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_816),
.B(n_505),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_L g981 ( 
.A(n_882),
.B(n_450),
.C(n_448),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_820),
.B(n_598),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_880),
.B(n_414),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_881),
.B(n_418),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_893),
.B(n_423),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_426),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_905),
.B(n_432),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_824),
.B(n_452),
.C(n_451),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_897),
.B(n_434),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_851),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_867),
.B(n_437),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_777),
.B(n_430),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_878),
.Y(n_993)
);

AO221x1_ASAP7_75t_L g994 ( 
.A1(n_793),
.A2(n_592),
.B1(n_622),
.B2(n_587),
.C(n_524),
.Y(n_994)
);

INVxp33_ASAP7_75t_L g995 ( 
.A(n_801),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_794),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_853),
.B(n_629),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_817),
.B(n_438),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_817),
.B(n_441),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_855),
.B(n_442),
.Y(n_1000)
);

INVx8_ASAP7_75t_L g1001 ( 
.A(n_795),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_891),
.B(n_521),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_891),
.B(n_526),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_857),
.B(n_444),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_858),
.B(n_445),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_891),
.B(n_529),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_859),
.B(n_446),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_784),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_891),
.B(n_531),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_798),
.B(n_465),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_787),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_791),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_860),
.B(n_885),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_776),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_906),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_909),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_852),
.B(n_454),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_852),
.B(n_463),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_849),
.B(n_478),
.C(n_471),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_851),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_783),
.B(n_486),
.C(n_479),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_825),
.B(n_468),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_900),
.B(n_470),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_L g1024 ( 
.A(n_903),
.B(n_491),
.C(n_490),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_865),
.B(n_534),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_864),
.B(n_472),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_818),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_797),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_781),
.B(n_495),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_900),
.B(n_782),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_829),
.B(n_484),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_799),
.B(n_488),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_800),
.B(n_494),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_811),
.B(n_544),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_803),
.B(n_496),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_814),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_838),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_840),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_842),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_786),
.B(n_500),
.C(n_498),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_795),
.B(n_497),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_811),
.B(n_499),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_924),
.A2(n_554),
.B(n_535),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_811),
.B(n_502),
.Y(n_1044)
);

AO221x1_ASAP7_75t_L g1045 ( 
.A1(n_921),
.A2(n_592),
.B1(n_622),
.B2(n_587),
.C(n_524),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_927),
.B(n_514),
.C(n_503),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_811),
.B(n_572),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_790),
.B(n_516),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_899),
.B(n_573),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_868),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_801),
.B(n_507),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_781),
.B(n_519),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_901),
.B(n_515),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_SL g1054 ( 
.A(n_802),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_939),
.Y(n_1055)
);

AND2x6_ASAP7_75t_SL g1056 ( 
.A(n_805),
.B(n_642),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_813),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_792),
.B(n_522),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_833),
.B(n_525),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_827),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_813),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_810),
.B(n_20),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_796),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_821),
.B(n_611),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_831),
.B(n_532),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_836),
.B(n_527),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_821),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_839),
.B(n_826),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_823),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_823),
.B(n_536),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_904),
.A2(n_410),
.B1(n_411),
.B2(n_408),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_847),
.B(n_612),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_537),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_847),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_910),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_779),
.B(n_538),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_871),
.B(n_617),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_883),
.B(n_618),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_808),
.B(n_540),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_887),
.B(n_619),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_894),
.B(n_631),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_809),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_779),
.B(n_543),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_856),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_895),
.B(n_645),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_895),
.B(n_648),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_907),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_941),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_918),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_912),
.B(n_656),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_835),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_921),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_886),
.B(n_560),
.C(n_558),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_888),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_804),
.B(n_565),
.C(n_562),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_896),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_870),
.B(n_568),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_898),
.B(n_541),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_841),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_917),
.B(n_545),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_919),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_L g1102 ( 
.A(n_861),
.B(n_544),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_911),
.B(n_550),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_913),
.B(n_555),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_922),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_850),
.B(n_556),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_923),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_914),
.B(n_563),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_926),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_928),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_929),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_930),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_915),
.B(n_567),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_933),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_935),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_938),
.Y(n_1116)
);

BUFx8_ASAP7_75t_L g1117 ( 
.A(n_834),
.Y(n_1117)
);

INVx8_ASAP7_75t_L g1118 ( 
.A(n_940),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_942),
.B(n_570),
.C(n_569),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_944),
.B(n_574),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_908),
.B(n_660),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_936),
.B(n_581),
.C(n_571),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_936),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_931),
.B(n_671),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_932),
.B(n_583),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_943),
.B(n_586),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_785),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_920),
.B(n_589),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_934),
.B(n_591),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_916),
.B(n_593),
.Y(n_1130)
);

INVxp33_ASAP7_75t_L g1131 ( 
.A(n_785),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_925),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_925),
.B(n_597),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_L g1134 ( 
.A(n_937),
.B(n_585),
.C(n_582),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_925),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_874),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_806),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_862),
.B(n_596),
.C(n_594),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_780),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_780),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_875),
.B(n_608),
.Y(n_1141)
);

INVxp33_ASAP7_75t_L g1142 ( 
.A(n_830),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_902),
.B(n_620),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_875),
.B(n_633),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_875),
.B(n_636),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_806),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_807),
.B(n_600),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_807),
.B(n_602),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_862),
.B(n_640),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_902),
.B(n_641),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_874),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_862),
.B(n_649),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_SL g1153 ( 
.A(n_848),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_862),
.B(n_651),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_875),
.B(n_652),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_875),
.B(n_653),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_902),
.B(n_654),
.Y(n_1157)
);

BUFx5_ASAP7_75t_L g1158 ( 
.A(n_851),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_875),
.B(n_658),
.Y(n_1159)
);

AO221x1_ASAP7_75t_L g1160 ( 
.A1(n_892),
.A2(n_644),
.B1(n_638),
.B2(n_609),
.C(n_599),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_862),
.B(n_667),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_807),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_875),
.B(n_670),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_875),
.B(n_412),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_970),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1162),
.B(n_638),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_961),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_952),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_SL g1169 ( 
.A(n_1082),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1162),
.Y(n_1170)
);

OR2x2_ASAP7_75t_SL g1171 ( 
.A(n_954),
.B(n_595),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_969),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_953),
.A2(n_646),
.B1(n_644),
.B2(n_415),
.Y(n_1173)
);

CKINVDCx11_ASAP7_75t_R g1174 ( 
.A(n_1056),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_996),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_953),
.B(n_634),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_977),
.B(n_607),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1137),
.Y(n_1178)
);

AND3x2_ASAP7_75t_SL g1179 ( 
.A(n_962),
.B(n_646),
.C(n_456),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_1001),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1001),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_965),
.B(n_635),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_977),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_965),
.B(n_637),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1142),
.B(n_643),
.Y(n_1185)
);

AND2x4_ASAP7_75t_SL g1186 ( 
.A(n_1075),
.B(n_458),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_949),
.A2(n_424),
.B(n_435),
.C(n_413),
.Y(n_1187)
);

AND2x6_ASAP7_75t_SL g1188 ( 
.A(n_1068),
.B(n_1106),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_949),
.A2(n_467),
.B1(n_482),
.B2(n_459),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_972),
.B(n_657),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_992),
.B(n_995),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1075),
.B(n_483),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_976),
.B(n_662),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1097),
.B(n_665),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1147),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1146),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_SL g1197 ( 
.A(n_1014),
.B(n_510),
.C(n_509),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

NOR2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1099),
.B(n_518),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_952),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1090),
.A2(n_523),
.B1(n_533),
.B2(n_530),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1122),
.B(n_971),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1118),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1148),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1090),
.A2(n_542),
.B1(n_551),
.B2(n_546),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_979),
.B(n_566),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_964),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_974),
.A2(n_577),
.B1(n_601),
.B2(n_588),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_993),
.B(n_948),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1071),
.A2(n_604),
.B1(n_615),
.B2(n_613),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1118),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1008),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1010),
.B(n_621),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1011),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_951),
.B(n_623),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1034),
.A2(n_624),
.B1(n_655),
.B2(n_625),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1012),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1118),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_981),
.B(n_666),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1013),
.B(n_668),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1138),
.B(n_672),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1127),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1136),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1048),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1060),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_947),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1151),
.Y(n_1227)
);

AND2x6_ASAP7_75t_L g1228 ( 
.A(n_1151),
.B(n_627),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1087),
.Y(n_1229)
);

NOR2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1054),
.B(n_630),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1028),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_947),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1117),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1036),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1037),
.B(n_630),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_967),
.A2(n_630),
.B1(n_627),
.B2(n_720),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1149),
.B(n_25),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1038),
.B(n_1039),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1065),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_967),
.B(n_1057),
.Y(n_1240)
);

NOR2x2_ASAP7_75t_L g1241 ( 
.A(n_994),
.B(n_25),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1105),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1100),
.B(n_627),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_990),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1029),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_966),
.B(n_720),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1164),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_986),
.B(n_724),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1164),
.Y(n_1249)
);

AND2x2_ASAP7_75t_SL g1250 ( 
.A(n_973),
.B(n_26),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_945),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1049),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_946),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1117),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1049),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1061),
.B(n_27),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1141),
.B(n_27),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1015),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1139),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1054),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1141),
.B(n_1144),
.Y(n_1261)
);

BUFx8_ASAP7_75t_L g1262 ( 
.A(n_1153),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_990),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1153),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1140),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1087),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1152),
.Y(n_1267)
);

XOR2xp5_ASAP7_75t_L g1268 ( 
.A(n_958),
.B(n_963),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1154),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1052),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1043),
.A2(n_743),
.B(n_739),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_978),
.B(n_991),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_990),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1161),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_975),
.A2(n_747),
.B1(n_750),
.B2(n_743),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1144),
.B(n_29),
.Y(n_1276)
);

NOR2x2_ASAP7_75t_L g1277 ( 
.A(n_1045),
.B(n_1160),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1087),
.Y(n_1278)
);

OR2x6_ASAP7_75t_L g1279 ( 
.A(n_955),
.B(n_743),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1016),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_975),
.A2(n_750),
.B1(n_757),
.B2(n_747),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1145),
.B(n_30),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1020),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1050),
.B(n_32),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1073),
.B(n_1083),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1002),
.A2(n_750),
.B1(n_757),
.B2(n_747),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_SL g1287 ( 
.A1(n_997),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1145),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1155),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_988),
.B(n_42),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1105),
.Y(n_1291)
);

INVx3_ASAP7_75t_SL g1292 ( 
.A(n_1051),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1092),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1003),
.A2(n_750),
.B1(n_757),
.B2(n_747),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1006),
.A2(n_759),
.B1(n_768),
.B2(n_757),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1020),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1062),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1030),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1089),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_987),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1009),
.A2(n_768),
.B1(n_770),
.B2(n_759),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1132),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_960),
.B(n_43),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1063),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1064),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1072),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1005),
.B(n_44),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1072),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1077),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_960),
.B(n_44),
.Y(n_1310)
);

OR2x4_ASAP7_75t_L g1311 ( 
.A(n_1079),
.B(n_45),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1025),
.B(n_48),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1069),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1111),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1156),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_950),
.B(n_1143),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1074),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1101),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_968),
.B(n_49),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1025),
.B(n_49),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1066),
.B(n_51),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1055),
.A2(n_770),
.B1(n_771),
.B2(n_768),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1078),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1088),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1046),
.B(n_770),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1080),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1042),
.B(n_771),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1047),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1047),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1124),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1159),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1041),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1124),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1112),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_SL g1335 ( 
.A(n_1095),
.B(n_1040),
.C(n_1021),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1084),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1000),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1084),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1080),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1163),
.B(n_61),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1123),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_985),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1107),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_1113),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_989),
.B(n_62),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1022),
.B(n_63),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1007),
.B(n_64),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1150),
.B(n_65),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1044),
.B(n_65),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1004),
.B(n_66),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1067),
.B(n_66),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1157),
.B(n_67),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1102),
.A2(n_197),
.B(n_193),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1024),
.B(n_69),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1094),
.B(n_1096),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1081),
.B(n_1085),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1076),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1081),
.B(n_72),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1132),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1032),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1085),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1109),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_956),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1033),
.A2(n_1035),
.B1(n_1031),
.B2(n_1093),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1086),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1026),
.B(n_77),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1121),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_957),
.B(n_80),
.Y(n_1368)
);

BUFx5_ASAP7_75t_L g1369 ( 
.A(n_1135),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1121),
.A2(n_84),
.B1(n_80),
.B2(n_81),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1110),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_980),
.B(n_81),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1134),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1023),
.A2(n_87),
.B(n_84),
.C(n_85),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1125),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1114),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1130),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_982),
.Y(n_1378)
);

AND2x6_ASAP7_75t_SL g1379 ( 
.A(n_1098),
.B(n_1104),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1115),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1070),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1116),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1130),
.B(n_201),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1119),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1019),
.B(n_88),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1108),
.Y(n_1386)
);

NOR2x2_ASAP7_75t_L g1387 ( 
.A(n_1017),
.B(n_89),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_959),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1158),
.Y(n_1389)
);

AO22x1_ASAP7_75t_L g1390 ( 
.A1(n_1059),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1133),
.Y(n_1391)
);

OR2x2_ASAP7_75t_SL g1392 ( 
.A(n_1018),
.B(n_92),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1058),
.B(n_94),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1170),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1356),
.A2(n_999),
.B1(n_998),
.B2(n_1120),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1250),
.A2(n_1194),
.B1(n_1245),
.B2(n_1315),
.Y(n_1396)
);

OAI21xp33_ASAP7_75t_L g1397 ( 
.A1(n_1190),
.A2(n_984),
.B(n_983),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1222),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_SL g1399 ( 
.A1(n_1220),
.A2(n_1126),
.B(n_1129),
.C(n_1128),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1356),
.A2(n_1240),
.B(n_1209),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1240),
.A2(n_1053),
.B(n_1131),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1180),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1260),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1195),
.B(n_1103),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1247),
.A2(n_1249),
.B1(n_1255),
.B2(n_1252),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1222),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1180),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1233),
.Y(n_1408)
);

NAND3x1_ASAP7_75t_L g1409 ( 
.A(n_1179),
.B(n_96),
.C(n_98),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1187),
.A2(n_99),
.B(n_96),
.C(n_98),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_R g1411 ( 
.A(n_1180),
.B(n_100),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1175),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1195),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1238),
.A2(n_1338),
.B(n_1336),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1181),
.B(n_101),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1204),
.B(n_103),
.Y(n_1416)
);

BUFx4f_ASAP7_75t_L g1417 ( 
.A(n_1254),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1204),
.B(n_1224),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1210),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_1419)
);

AOI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1353),
.A2(n_1377),
.B1(n_1375),
.B2(n_1271),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1212),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1181),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1331),
.B(n_110),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1214),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1305),
.A2(n_219),
.B(n_217),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1306),
.A2(n_1309),
.B(n_1308),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1262),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1181),
.B(n_1198),
.Y(n_1428)
);

CKINVDCx6p67_ASAP7_75t_R g1429 ( 
.A(n_1198),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1217),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1323),
.B(n_115),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1231),
.Y(n_1432)
);

BUFx4_ASAP7_75t_SL g1433 ( 
.A(n_1348),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1225),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1326),
.B(n_116),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1234),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1171),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1173),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1189),
.A2(n_121),
.B(n_122),
.C(n_124),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1262),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1339),
.B(n_125),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1302),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1166),
.B(n_125),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1193),
.B(n_126),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1256),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1361),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1186),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1285),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1448)
);

INVx8_ASAP7_75t_L g1449 ( 
.A(n_1203),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1183),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1201),
.B(n_1367),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1365),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1383),
.A2(n_232),
.B(n_230),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1327),
.A2(n_235),
.B(n_234),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1257),
.A2(n_136),
.B(n_137),
.C(n_140),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1383),
.A2(n_240),
.B(n_237),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1270),
.B(n_140),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1198),
.B(n_141),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1192),
.B(n_141),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1201),
.B(n_142),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1330),
.A2(n_245),
.B(n_241),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1269),
.B(n_143),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1300),
.B(n_144),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1205),
.B(n_145),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1303),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1211),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1333),
.A2(n_307),
.B(n_388),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1192),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1351),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_SL g1470 ( 
.A(n_1363),
.B(n_146),
.C(n_151),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1239),
.B(n_152),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_R g1472 ( 
.A(n_1174),
.B(n_155),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1185),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1351),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1386),
.B(n_160),
.Y(n_1475)
);

AND2x2_ASAP7_75t_SL g1476 ( 
.A(n_1284),
.B(n_160),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1176),
.B(n_1213),
.Y(n_1477)
);

INVx11_ASAP7_75t_L g1478 ( 
.A(n_1228),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1324),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1165),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1169),
.Y(n_1481)
);

NOR3xp33_ASAP7_75t_SL g1482 ( 
.A(n_1335),
.B(n_163),
.C(n_164),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1303),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1191),
.B(n_164),
.Y(n_1484)
);

OA22x2_ASAP7_75t_L g1485 ( 
.A1(n_1348),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1202),
.B(n_1342),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1310),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1218),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1310),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1378),
.B(n_169),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1202),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1312),
.A2(n_252),
.B(n_254),
.C(n_257),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1381),
.B(n_268),
.Y(n_1493)
);

XNOR2xp5_ASAP7_75t_L g1494 ( 
.A(n_1268),
.B(n_270),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1359),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1359),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1229),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1229),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1313),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1341),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1337),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1312),
.A2(n_278),
.B(n_279),
.C(n_281),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1320),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1355),
.A2(n_1282),
.B(n_1276),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1226),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1167),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1169),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1272),
.B(n_390),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1388),
.B(n_287),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1272),
.B(n_1299),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1228),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1291),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1172),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1348),
.B(n_291),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1340),
.A2(n_297),
.B(n_300),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1248),
.A2(n_303),
.B(n_304),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1345),
.A2(n_315),
.B(n_316),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1352),
.B(n_317),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1352),
.B(n_1206),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1358),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1251),
.Y(n_1521)
);

AO32x1_ASAP7_75t_L g1522 ( 
.A1(n_1370),
.A2(n_326),
.A3(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1197),
.A2(n_345),
.B(n_346),
.C(n_347),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1374),
.A2(n_1216),
.B(n_1208),
.C(n_1346),
.Y(n_1524)
);

BUFx4_ASAP7_75t_SL g1525 ( 
.A(n_1188),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1267),
.B(n_349),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1274),
.B(n_353),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1362),
.Y(n_1528)
);

NAND2x2_ASAP7_75t_L g1529 ( 
.A(n_1199),
.B(n_356),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1178),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1316),
.B(n_358),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1253),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1188),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1232),
.B(n_1264),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1314),
.B(n_366),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1230),
.B(n_369),
.Y(n_1536)
);

BUFx4f_ASAP7_75t_L g1537 ( 
.A(n_1292),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1266),
.Y(n_1538)
);

INVx5_ASAP7_75t_L g1539 ( 
.A(n_1228),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1334),
.B(n_375),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1284),
.Y(n_1541)
);

OAI22x1_ASAP7_75t_L g1542 ( 
.A1(n_1354),
.A2(n_378),
.B1(n_1329),
.B2(n_1347),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1372),
.A2(n_1368),
.B(n_1373),
.C(n_1384),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1237),
.A2(n_1393),
.B(n_1364),
.C(n_1329),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1311),
.A2(n_1392),
.B1(n_1287),
.B2(n_1288),
.Y(n_1545)
);

AO21x1_ASAP7_75t_L g1546 ( 
.A1(n_1370),
.A2(n_1236),
.B(n_1235),
.Y(n_1546)
);

AOI221x1_ASAP7_75t_L g1547 ( 
.A1(n_1236),
.A2(n_1289),
.B1(n_1288),
.B2(n_1354),
.C(n_1287),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1200),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1215),
.B(n_1219),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1307),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_SL g1551 ( 
.A(n_1332),
.B(n_1357),
.C(n_1289),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1371),
.B(n_1382),
.Y(n_1552)
);

OR2x6_ASAP7_75t_L g1553 ( 
.A(n_1307),
.B(n_1347),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1290),
.A2(n_1319),
.B1(n_1219),
.B2(n_1221),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1259),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1321),
.Y(n_1556)
);

O2A1O1Ixp5_ASAP7_75t_L g1557 ( 
.A1(n_1243),
.A2(n_1325),
.B(n_1349),
.C(n_1366),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1196),
.A2(n_1350),
.B(n_1235),
.C(n_1221),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1328),
.A2(n_1360),
.B1(n_1385),
.B2(n_1380),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1318),
.B(n_1343),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1304),
.A2(n_1317),
.B1(n_1280),
.B2(n_1258),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1318),
.B(n_1242),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1242),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1341),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1296),
.B(n_1227),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1376),
.B(n_1379),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1265),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1376),
.B(n_1379),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_L g1570 ( 
.A(n_1390),
.B(n_1293),
.C(n_1298),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1317),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1391),
.B(n_1246),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1297),
.B(n_1177),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1207),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1344),
.B(n_1207),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1281),
.A2(n_1294),
.B(n_1301),
.C(n_1295),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1296),
.B(n_1168),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1344),
.B(n_1168),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1223),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1223),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1278),
.B(n_1244),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1228),
.Y(n_1582)
);

AOI221x1_ASAP7_75t_L g1583 ( 
.A1(n_1389),
.A2(n_1283),
.B1(n_1244),
.B2(n_1263),
.C(n_1273),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1279),
.A2(n_1275),
.B(n_1286),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1322),
.A2(n_1277),
.B(n_1241),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1387),
.B(n_1369),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1369),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1356),
.A2(n_1247),
.B1(n_1249),
.B2(n_1252),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1192),
.B(n_1001),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1195),
.B(n_1142),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1356),
.A2(n_1247),
.B1(n_1249),
.B2(n_1252),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1187),
.A2(n_1261),
.B(n_953),
.C(n_1210),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1170),
.Y(n_1597)
);

CKINVDCx14_ASAP7_75t_R g1598 ( 
.A(n_1174),
.Y(n_1598)
);

NOR2xp67_ASAP7_75t_SL g1599 ( 
.A(n_1180),
.B(n_1181),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1260),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1250),
.A2(n_1160),
.B1(n_1045),
.B2(n_968),
.Y(n_1603)
);

NOR3xp33_ASAP7_75t_L g1604 ( 
.A(n_1335),
.B(n_1197),
.C(n_1269),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1180),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1356),
.A2(n_1247),
.B1(n_1249),
.B2(n_1252),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1170),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1180),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1180),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1336),
.A2(n_1091),
.B(n_1027),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1613)
);

INVx5_ASAP7_75t_L g1614 ( 
.A(n_1228),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1356),
.A2(n_1247),
.B1(n_1249),
.B2(n_1252),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1261),
.A2(n_927),
.B(n_907),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1261),
.A2(n_927),
.B(n_907),
.Y(n_1618)
);

OA22x2_ASAP7_75t_L g1619 ( 
.A1(n_1170),
.A2(n_1160),
.B1(n_1162),
.B2(n_994),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1220),
.B(n_1190),
.C(n_882),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1195),
.B(n_1142),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1261),
.A2(n_927),
.B(n_907),
.Y(n_1624)
);

INVx8_ASAP7_75t_L g1625 ( 
.A(n_1203),
.Y(n_1625)
);

INVx6_ASAP7_75t_L g1626 ( 
.A(n_1180),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1170),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1180),
.B(n_1181),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1408),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1449),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1449),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1417),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1417),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1421),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1610),
.A2(n_1420),
.B(n_1414),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1453),
.A2(n_1456),
.B(n_1583),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1543),
.A2(n_1559),
.B(n_1546),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1403),
.Y(n_1641)
);

BUFx12f_ASAP7_75t_L g1642 ( 
.A(n_1427),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1593),
.A2(n_1616),
.B(n_1606),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1400),
.A2(n_1618),
.B(n_1617),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1590),
.B(n_1601),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1646)
);

BUFx4f_ASAP7_75t_SL g1647 ( 
.A(n_1429),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1447),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1449),
.Y(n_1649)
);

INVx6_ASAP7_75t_L g1650 ( 
.A(n_1625),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1591),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1554),
.B(n_1486),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1625),
.B(n_1591),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1615),
.Y(n_1654)
);

AOI22x1_ASAP7_75t_L g1655 ( 
.A1(n_1542),
.A2(n_1504),
.B1(n_1584),
.B2(n_1517),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1424),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1630),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1624),
.A2(n_1426),
.B(n_1544),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1625),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1428),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1430),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1432),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1402),
.B(n_1422),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1402),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1422),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1413),
.Y(n_1666)
);

INVx6_ASAP7_75t_SL g1667 ( 
.A(n_1514),
.Y(n_1667)
);

NAND2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1605),
.B(n_1511),
.Y(n_1668)
);

AO21x2_ASAP7_75t_L g1669 ( 
.A1(n_1570),
.A2(n_1576),
.B(n_1524),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1503),
.A2(n_1483),
.B(n_1465),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1436),
.Y(n_1671)
);

BUFx4f_ASAP7_75t_SL g1672 ( 
.A(n_1582),
.Y(n_1672)
);

INVx8_ASAP7_75t_L g1673 ( 
.A(n_1514),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1407),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1622),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1628),
.B(n_1468),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1487),
.A2(n_1489),
.B(n_1445),
.Y(n_1677)
);

BUFx12f_ASAP7_75t_L g1678 ( 
.A(n_1440),
.Y(n_1678)
);

INVx5_ASAP7_75t_L g1679 ( 
.A(n_1511),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1451),
.B(n_1405),
.Y(n_1680)
);

INVx5_ASAP7_75t_SL g1681 ( 
.A(n_1478),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1506),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1461),
.A2(n_1467),
.B(n_1515),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1605),
.B(n_1608),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1537),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1450),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1513),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1415),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1530),
.Y(n_1690)
);

BUFx12f_ASAP7_75t_L g1691 ( 
.A(n_1600),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1476),
.B(n_1586),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1497),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1594),
.B(n_1477),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1609),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1394),
.Y(n_1696)
);

AO21x2_ASAP7_75t_L g1697 ( 
.A1(n_1431),
.A2(n_1441),
.B(n_1435),
.Y(n_1697)
);

INVx8_ASAP7_75t_L g1698 ( 
.A(n_1415),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1537),
.Y(n_1699)
);

BUFx12f_ASAP7_75t_L g1700 ( 
.A(n_1528),
.Y(n_1700)
);

BUFx12f_ASAP7_75t_L g1701 ( 
.A(n_1481),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1592),
.B(n_1621),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1545),
.A2(n_1604),
.B1(n_1586),
.B2(n_1438),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1609),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1553),
.A2(n_1437),
.B1(n_1619),
.B2(n_1603),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1492),
.A2(n_1502),
.B(n_1425),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_SL g1707 ( 
.A1(n_1567),
.A2(n_1569),
.B(n_1396),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1500),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1553),
.B(n_1508),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1626),
.Y(n_1710)
);

BUFx12f_ASAP7_75t_L g1711 ( 
.A(n_1507),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1626),
.Y(n_1712)
);

INVx3_ASAP7_75t_SL g1713 ( 
.A(n_1458),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1434),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1568),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1508),
.B(n_1572),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1560),
.A2(n_1399),
.B(n_1493),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1581),
.A2(n_1516),
.B(n_1454),
.Y(n_1718)
);

CKINVDCx16_ASAP7_75t_R g1719 ( 
.A(n_1411),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1566),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1547),
.A2(n_1557),
.B(n_1452),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1597),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1548),
.Y(n_1723)
);

BUFx5_ASAP7_75t_L g1724 ( 
.A(n_1577),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1550),
.B(n_1473),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1511),
.B(n_1539),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1412),
.Y(n_1727)
);

BUFx2_ASAP7_75t_R g1728 ( 
.A(n_1533),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1418),
.B(n_1627),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1433),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1466),
.Y(n_1731)
);

BUFx4_ASAP7_75t_SL g1732 ( 
.A(n_1536),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1406),
.Y(n_1733)
);

CKINVDCx16_ASAP7_75t_R g1734 ( 
.A(n_1472),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1536),
.B(n_1458),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1574),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1519),
.B(n_1620),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1575),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1541),
.B(n_1549),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1571),
.Y(n_1740)
);

BUFx2_ASAP7_75t_SL g1741 ( 
.A(n_1539),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1536),
.B(n_1485),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1572),
.B(n_1510),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1512),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1589),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1443),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1398),
.Y(n_1747)
);

INVx4_ASAP7_75t_L g1748 ( 
.A(n_1539),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1595),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1498),
.A2(n_1520),
.B(n_1523),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1560),
.A2(n_1518),
.B(n_1455),
.Y(n_1752)
);

BUFx2_ASAP7_75t_R g1753 ( 
.A(n_1529),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1607),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1401),
.A2(n_1423),
.B(n_1522),
.Y(n_1755)
);

OAI21x1_ASAP7_75t_L g1756 ( 
.A1(n_1540),
.A2(n_1499),
.B(n_1563),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1587),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1521),
.Y(n_1758)
);

OA21x2_ASAP7_75t_L g1759 ( 
.A1(n_1491),
.A2(n_1460),
.B(n_1479),
.Y(n_1759)
);

OR2x6_ASAP7_75t_L g1760 ( 
.A(n_1505),
.B(n_1459),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1532),
.Y(n_1761)
);

BUFx8_ASAP7_75t_L g1762 ( 
.A(n_1510),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1555),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1596),
.B(n_1602),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1480),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1614),
.Y(n_1766)
);

BUFx2_ASAP7_75t_R g1767 ( 
.A(n_1494),
.Y(n_1767)
);

INVx5_ASAP7_75t_L g1768 ( 
.A(n_1614),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1579),
.A2(n_1580),
.B(n_1562),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1623),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1629),
.B(n_1551),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1488),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1446),
.Y(n_1773)
);

AO21x2_ASAP7_75t_L g1774 ( 
.A1(n_1469),
.A2(n_1474),
.B(n_1470),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1410),
.A2(n_1561),
.B(n_1395),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1564),
.B(n_1444),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1404),
.B(n_1573),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1484),
.B(n_1464),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1462),
.B(n_1397),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1552),
.B(n_1578),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1475),
.B(n_1463),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1409),
.B(n_1439),
.Y(n_1782)
);

CKINVDCx6p67_ASAP7_75t_R g1783 ( 
.A(n_1556),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1419),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1565),
.Y(n_1785)
);

AO21x2_ASAP7_75t_L g1786 ( 
.A1(n_1585),
.A2(n_1501),
.B(n_1531),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1457),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1471),
.Y(n_1788)
);

INVx6_ASAP7_75t_SL g1789 ( 
.A(n_1598),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_L g1790 ( 
.A(n_1538),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1482),
.A2(n_1535),
.B(n_1522),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1442),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1490),
.Y(n_1793)
);

BUFx4f_ASAP7_75t_L g1794 ( 
.A(n_1525),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1416),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1526),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1558),
.B(n_1509),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1495),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1448),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1527),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1534),
.Y(n_1801)
);

NAND2x1_ASAP7_75t_L g1802 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1413),
.Y(n_1803)
);

INVx4_ASAP7_75t_SL g1804 ( 
.A(n_1582),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1545),
.A2(n_1604),
.B1(n_1476),
.B2(n_1250),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1421),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1449),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_1447),
.Y(n_1808)
);

OR2x6_ASAP7_75t_L g1809 ( 
.A(n_1449),
.B(n_1625),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1449),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1449),
.Y(n_1811)
);

INVx6_ASAP7_75t_L g1812 ( 
.A(n_1449),
.Y(n_1812)
);

AO21x2_ASAP7_75t_L g1813 ( 
.A1(n_1543),
.A2(n_1559),
.B(n_1546),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1591),
.B(n_1630),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1413),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1449),
.Y(n_1816)
);

BUFx10_ASAP7_75t_L g1817 ( 
.A(n_1630),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1694),
.B(n_1680),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1636),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1656),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1735),
.B(n_1688),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1661),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1662),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1666),
.Y(n_1824)
);

CKINVDCx6p67_ASAP7_75t_R g1825 ( 
.A(n_1641),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1694),
.B(n_1680),
.Y(n_1826)
);

INVx6_ASAP7_75t_L g1827 ( 
.A(n_1816),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1742),
.A2(n_1805),
.B1(n_1673),
.B2(n_1703),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1667),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1643),
.B(n_1639),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1816),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1735),
.A2(n_1643),
.B1(n_1639),
.B2(n_1667),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1637),
.A2(n_1638),
.B(n_1755),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1647),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1647),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1682),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1809),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1687),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1671),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1809),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1675),
.B(n_1676),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1808),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1659),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1809),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1659),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1735),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1659),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_SL g1848 ( 
.A1(n_1673),
.A2(n_1688),
.B1(n_1692),
.B2(n_1709),
.Y(n_1848)
);

OAI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1673),
.A2(n_1742),
.B1(n_1675),
.B2(n_1645),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1742),
.A2(n_1805),
.B1(n_1703),
.B2(n_1652),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1690),
.Y(n_1851)
);

INVx4_ASAP7_75t_L g1852 ( 
.A(n_1810),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1808),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1631),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1806),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1810),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1709),
.B(n_1653),
.Y(n_1857)
);

INVx6_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1645),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1702),
.B(n_1793),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1715),
.Y(n_1861)
);

OA21x2_ASAP7_75t_L g1862 ( 
.A1(n_1655),
.A2(n_1644),
.B(n_1658),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1758),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1761),
.Y(n_1864)
);

CKINVDCx11_ASAP7_75t_R g1865 ( 
.A(n_1691),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1810),
.Y(n_1866)
);

INVx4_ASAP7_75t_SL g1867 ( 
.A(n_1713),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1705),
.A2(n_1782),
.B1(n_1737),
.B2(n_1779),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1646),
.A2(n_1654),
.B1(n_1713),
.B2(n_1689),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1763),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1747),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1747),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1765),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1653),
.B(n_1716),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1632),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1792),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1782),
.A2(n_1737),
.B1(n_1773),
.B2(n_1784),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1666),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1653),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1782),
.A2(n_1799),
.B1(n_1778),
.B2(n_1781),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1650),
.Y(n_1881)
);

BUFx2_ASAP7_75t_SL g1882 ( 
.A(n_1634),
.Y(n_1882)
);

NAND2x1p5_ASAP7_75t_L g1883 ( 
.A(n_1649),
.B(n_1679),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1660),
.Y(n_1884)
);

OA21x2_ASAP7_75t_L g1885 ( 
.A1(n_1658),
.A2(n_1706),
.B(n_1751),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1650),
.Y(n_1886)
);

BUFx2_ASAP7_75t_R g1887 ( 
.A(n_1730),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1631),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1646),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1654),
.B(n_1670),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1814),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1650),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1670),
.B(n_1677),
.Y(n_1893)
);

NAND2x1p5_ASAP7_75t_L g1894 ( 
.A(n_1679),
.B(n_1768),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1698),
.A2(n_1716),
.B1(n_1732),
.B2(n_1719),
.Y(n_1895)
);

AOI222xp33_ASAP7_75t_L g1896 ( 
.A1(n_1794),
.A2(n_1777),
.B1(n_1746),
.B2(n_1677),
.C1(n_1739),
.C2(n_1730),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1778),
.A2(n_1781),
.B1(n_1795),
.B2(n_1788),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_SL g1898 ( 
.A1(n_1698),
.A2(n_1732),
.B1(n_1651),
.B2(n_1707),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1698),
.A2(n_1796),
.B1(n_1722),
.B2(n_1669),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_SL g1900 ( 
.A1(n_1796),
.A2(n_1696),
.B1(n_1731),
.B2(n_1774),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_SL g1901 ( 
.A1(n_1774),
.A2(n_1740),
.B1(n_1734),
.B2(n_1760),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1729),
.B(n_1803),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1787),
.A2(n_1797),
.B1(n_1800),
.B2(n_1771),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1812),
.Y(n_1904)
);

CKINVDCx11_ASAP7_75t_R g1905 ( 
.A(n_1642),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1760),
.A2(n_1749),
.B1(n_1770),
.B2(n_1745),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1812),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1764),
.Y(n_1908)
);

CKINVDCx11_ASAP7_75t_R g1909 ( 
.A(n_1678),
.Y(n_1909)
);

CKINVDCx16_ASAP7_75t_R g1910 ( 
.A(n_1635),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1764),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1760),
.A2(n_1752),
.B1(n_1754),
.B2(n_1725),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1738),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1756),
.A2(n_1775),
.B(n_1683),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1663),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1679),
.B(n_1768),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1663),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1633),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1745),
.A2(n_1770),
.B1(n_1749),
.B2(n_1744),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1776),
.A2(n_1686),
.B1(n_1714),
.B2(n_1812),
.Y(n_1920)
);

BUFx8_ASAP7_75t_L g1921 ( 
.A(n_1700),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1776),
.A2(n_1686),
.B1(n_1780),
.B2(n_1815),
.Y(n_1922)
);

OAI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1744),
.A2(n_1815),
.B1(n_1803),
.B2(n_1794),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1772),
.Y(n_1924)
);

INVx6_ASAP7_75t_L g1925 ( 
.A(n_1817),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1801),
.A2(n_1733),
.B1(n_1786),
.B2(n_1780),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1811),
.B(n_1684),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1648),
.A2(n_1633),
.B1(n_1807),
.B2(n_1743),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1807),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1757),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1789),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1693),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1757),
.Y(n_1933)
);

OAI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1657),
.A2(n_1672),
.B1(n_1679),
.B2(n_1768),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1718),
.A2(n_1769),
.B(n_1802),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1859),
.B(n_1724),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1841),
.B(n_1727),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1902),
.B(n_1785),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1825),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1819),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1865),
.Y(n_1941)
);

AO21x1_ASAP7_75t_L g1942 ( 
.A1(n_1869),
.A2(n_1657),
.B(n_1668),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1905),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1820),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1932),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1822),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1909),
.Y(n_1947)
);

CKINVDCx16_ASAP7_75t_R g1948 ( 
.A(n_1884),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1927),
.B(n_1674),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1823),
.Y(n_1950)
);

INVx4_ASAP7_75t_L g1951 ( 
.A(n_1827),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1859),
.B(n_1664),
.Y(n_1952)
);

NAND2xp33_ASAP7_75t_R g1953 ( 
.A(n_1931),
.B(n_1648),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1871),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1852),
.Y(n_1955)
);

OR2x4_ASAP7_75t_L g1956 ( 
.A(n_1915),
.B(n_1753),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1860),
.B(n_1665),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1850),
.A2(n_1786),
.B1(n_1697),
.B2(n_1813),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1836),
.Y(n_1959)
);

CKINVDCx16_ASAP7_75t_R g1960 ( 
.A(n_1834),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1838),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1831),
.B(n_1768),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1896),
.A2(n_1704),
.B(n_1695),
.C(n_1717),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1824),
.B(n_1724),
.Y(n_1964)
);

CKINVDCx11_ASAP7_75t_R g1965 ( 
.A(n_1835),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1824),
.B(n_1724),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1878),
.B(n_1720),
.Y(n_1967)
);

CKINVDCx14_ASAP7_75t_R g1968 ( 
.A(n_1854),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1849),
.A2(n_1753),
.B1(n_1767),
.B2(n_1721),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_R g1970 ( 
.A(n_1831),
.B(n_1695),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1890),
.B(n_1640),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1851),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1871),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1855),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1896),
.A2(n_1717),
.B1(n_1721),
.B2(n_1697),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1921),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1921),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1888),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_R g1979 ( 
.A(n_1910),
.B(n_1672),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1889),
.B(n_1762),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1897),
.B(n_1762),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1849),
.A2(n_1767),
.B1(n_1668),
.B2(n_1681),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1821),
.B(n_1723),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_R g1984 ( 
.A(n_1837),
.B(n_1789),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_R g1985 ( 
.A(n_1875),
.B(n_1723),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_SL g1986 ( 
.A1(n_1832),
.A2(n_1741),
.B1(n_1791),
.B2(n_1813),
.Y(n_1986)
);

NOR3xp33_ASAP7_75t_SL g1987 ( 
.A(n_1923),
.B(n_1728),
.C(n_1783),
.Y(n_1987)
);

INVx2_ASAP7_75t_SL g1988 ( 
.A(n_1827),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1878),
.B(n_1720),
.Y(n_1989)
);

NOR3xp33_ASAP7_75t_SL g1990 ( 
.A(n_1923),
.B(n_1728),
.C(n_1804),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1821),
.B(n_1736),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1894),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1887),
.Y(n_1993)
);

OR2x6_ASAP7_75t_L g1994 ( 
.A(n_1832),
.B(n_1726),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1872),
.B(n_1736),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1887),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1872),
.B(n_1712),
.Y(n_1997)
);

NAND3xp33_ASAP7_75t_SL g1998 ( 
.A(n_1895),
.B(n_1750),
.C(n_1726),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1882),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1828),
.A2(n_1681),
.B1(n_1750),
.B2(n_1759),
.Y(n_2000)
);

CKINVDCx16_ASAP7_75t_R g2001 ( 
.A(n_1842),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1876),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_1853),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1903),
.B(n_1640),
.Y(n_2004)
);

NAND3xp33_ASAP7_75t_SL g2005 ( 
.A(n_1895),
.B(n_1798),
.C(n_1748),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1861),
.B(n_1804),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1863),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1852),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1848),
.A2(n_1699),
.B1(n_1685),
.B2(n_1701),
.Y(n_2009)
);

OAI21xp33_ASAP7_75t_L g2010 ( 
.A1(n_1900),
.A2(n_1710),
.B(n_1798),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1839),
.B(n_1868),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1864),
.Y(n_2012)
);

OR2x6_ASAP7_75t_L g2013 ( 
.A(n_1916),
.B(n_1748),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_R g2014 ( 
.A(n_1827),
.B(n_1711),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1922),
.B(n_1804),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1916),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1945),
.B(n_1830),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1945),
.B(n_1830),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1971),
.B(n_2004),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1955),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1971),
.B(n_1862),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1940),
.B(n_1944),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_2008),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_SL g2024 ( 
.A1(n_1982),
.A2(n_1846),
.B1(n_1879),
.B2(n_1844),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1946),
.B(n_1862),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1942),
.B(n_1898),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1954),
.B(n_1818),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2012),
.B(n_1930),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1950),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2007),
.B(n_1933),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1973),
.B(n_2002),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1959),
.B(n_1961),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1972),
.B(n_1926),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1974),
.B(n_1826),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1982),
.A2(n_1880),
.B1(n_1877),
.B2(n_1901),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1994),
.B(n_1935),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1957),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1958),
.B(n_1908),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1958),
.B(n_1911),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1995),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1952),
.B(n_1870),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1985),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1956),
.A2(n_1898),
.B1(n_1848),
.B2(n_1901),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1975),
.B(n_1964),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1966),
.B(n_1893),
.Y(n_2045)
);

OAI222xp33_ASAP7_75t_L g2046 ( 
.A1(n_1969),
.A2(n_1900),
.B1(n_1899),
.B2(n_1906),
.C1(n_1846),
.C2(n_1912),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1997),
.B(n_1873),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1936),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1994),
.Y(n_2049)
);

NAND4xp25_ASAP7_75t_L g2050 ( 
.A(n_1963),
.B(n_1969),
.C(n_1899),
.D(n_1981),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2009),
.A2(n_1934),
.B1(n_1867),
.B2(n_1858),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2034),
.B(n_2011),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_2020),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_2020),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2025),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2045),
.B(n_1986),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_2031),
.B(n_1938),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_2042),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2025),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2031),
.B(n_2000),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_2036),
.B(n_1994),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2024),
.A2(n_1956),
.B1(n_2009),
.B2(n_1906),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2029),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2027),
.B(n_1937),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_2023),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2034),
.B(n_1967),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2045),
.B(n_1885),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_2036),
.B(n_2049),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2027),
.B(n_1876),
.Y(n_2069)
);

NAND2x1_ASAP7_75t_SL g2070 ( 
.A(n_2051),
.B(n_1951),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2019),
.B(n_1833),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2022),
.B(n_1989),
.Y(n_2072)
);

NOR2xp67_ASAP7_75t_L g2073 ( 
.A(n_2051),
.B(n_1999),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2019),
.B(n_1833),
.Y(n_2074)
);

NAND2x1_ASAP7_75t_SL g2075 ( 
.A(n_2036),
.B(n_1951),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2022),
.B(n_1919),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2021),
.B(n_1914),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2021),
.B(n_1914),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2033),
.B(n_1919),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2055),
.B(n_2033),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2067),
.B(n_2044),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2067),
.B(n_2044),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2055),
.B(n_2018),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2063),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2077),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2077),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2071),
.B(n_2017),
.Y(n_2087)
);

AND2x4_ASAP7_75t_SL g2088 ( 
.A(n_2061),
.B(n_2049),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2063),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_2068),
.B(n_2036),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2059),
.B(n_2018),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2059),
.B(n_2048),
.Y(n_2092)
);

OR2x6_ASAP7_75t_L g2093 ( 
.A(n_2061),
.B(n_2026),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2062),
.A2(n_2050),
.B1(n_2043),
.B2(n_2035),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2052),
.B(n_2048),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2078),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2071),
.B(n_2017),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2053),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2074),
.B(n_2038),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2064),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2074),
.B(n_2038),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2078),
.B(n_2056),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2056),
.B(n_2039),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2068),
.B(n_2039),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2103),
.B(n_2079),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2092),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2102),
.B(n_2068),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_2090),
.Y(n_2108)
);

OAI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_2094),
.A2(n_2073),
.B(n_2070),
.C(n_2050),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_2090),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2083),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2084),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2084),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2102),
.B(n_2065),
.Y(n_2114)
);

OAI33xp33_ASAP7_75t_L g2115 ( 
.A1(n_2095),
.A2(n_2058),
.A3(n_2057),
.B1(n_2064),
.B2(n_2072),
.B3(n_2066),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_2090),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2083),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2091),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_L g2119 ( 
.A(n_2093),
.B(n_2058),
.C(n_2054),
.Y(n_2119)
);

A2O1A1Ixp33_ASAP7_75t_L g2120 ( 
.A1(n_2088),
.A2(n_2070),
.B(n_1987),
.C(n_1990),
.Y(n_2120)
);

NOR2x1p5_ASAP7_75t_L g2121 ( 
.A(n_2090),
.B(n_1993),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2091),
.Y(n_2122)
);

NAND2x2_ASAP7_75t_L g2123 ( 
.A(n_2093),
.B(n_2060),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2085),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2089),
.Y(n_2125)
);

NOR2x1p5_ASAP7_75t_L g2126 ( 
.A(n_2103),
.B(n_1996),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2089),
.Y(n_2127)
);

OA222x2_ASAP7_75t_L g2128 ( 
.A1(n_2093),
.A2(n_2060),
.B1(n_2057),
.B2(n_2069),
.C1(n_2085),
.C2(n_2086),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_2093),
.B(n_2061),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2085),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2100),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2128),
.B(n_2104),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2125),
.Y(n_2133)
);

OAI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2109),
.A2(n_2093),
.B1(n_2098),
.B2(n_2054),
.C(n_1984),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2115),
.A2(n_2082),
.B1(n_2081),
.B2(n_2104),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2123),
.A2(n_2088),
.B1(n_2037),
.B2(n_2040),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_2131),
.Y(n_2137)
);

OAI21xp33_ASAP7_75t_L g2138 ( 
.A1(n_2119),
.A2(n_2082),
.B(n_2081),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2127),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2107),
.B(n_2087),
.Y(n_2140)
);

NAND3xp33_ASAP7_75t_SL g2141 ( 
.A(n_2120),
.B(n_2014),
.C(n_1979),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2126),
.A2(n_2088),
.B1(n_2101),
.B2(n_2099),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2112),
.Y(n_2143)
);

NAND3xp33_ASAP7_75t_SL g2144 ( 
.A(n_2120),
.B(n_1976),
.C(n_2003),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2124),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2123),
.A2(n_2101),
.B1(n_2099),
.B2(n_2076),
.Y(n_2146)
);

OAI21xp33_ASAP7_75t_L g2147 ( 
.A1(n_2129),
.A2(n_2080),
.B(n_2086),
.Y(n_2147)
);

A2O1A1Ixp33_ASAP7_75t_L g2148 ( 
.A1(n_2121),
.A2(n_2075),
.B(n_1998),
.C(n_2096),
.Y(n_2148)
);

XOR2xp5_ASAP7_75t_L g2149 ( 
.A(n_2129),
.B(n_1977),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2135),
.B(n_2106),
.Y(n_2150)
);

OAI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2134),
.A2(n_2116),
.B1(n_2108),
.B2(n_2110),
.C(n_2122),
.Y(n_2151)
);

INVxp67_ASAP7_75t_SL g2152 ( 
.A(n_2137),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2133),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2139),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2132),
.B(n_2114),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2145),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2143),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_SL g2158 ( 
.A1(n_2134),
.A2(n_2129),
.B1(n_2110),
.B2(n_2108),
.Y(n_2158)
);

OAI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_2144),
.A2(n_2116),
.B1(n_2108),
.B2(n_2110),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_2141),
.A2(n_1980),
.B1(n_2015),
.B2(n_2116),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2148),
.B(n_2114),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2138),
.A2(n_2118),
.B1(n_2117),
.B2(n_2111),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2136),
.A2(n_2142),
.B(n_2146),
.C(n_2147),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2149),
.Y(n_2164)
);

OAI221xp5_ASAP7_75t_L g2165 ( 
.A1(n_2136),
.A2(n_2105),
.B1(n_2010),
.B2(n_2124),
.C(n_2130),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2140),
.B(n_2107),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2137),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_2137),
.Y(n_2168)
);

INVx1_ASAP7_75t_SL g2169 ( 
.A(n_2149),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2168),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2152),
.B(n_2112),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2168),
.Y(n_2172)
);

AOI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_2167),
.A2(n_2001),
.B1(n_2010),
.B2(n_1948),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_SL g2174 ( 
.A1(n_2163),
.A2(n_1939),
.B(n_1941),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_2169),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_2164),
.B(n_1943),
.Y(n_2176)
);

NOR3x1_ASAP7_75t_L g2177 ( 
.A(n_2151),
.B(n_1829),
.C(n_2005),
.Y(n_2177)
);

OA22x2_ASAP7_75t_L g2178 ( 
.A1(n_2161),
.A2(n_1947),
.B1(n_1978),
.B2(n_1920),
.Y(n_2178)
);

NAND3xp33_ASAP7_75t_L g2179 ( 
.A(n_2158),
.B(n_2159),
.C(n_2150),
.Y(n_2179)
);

AOI211xp5_ASAP7_75t_L g2180 ( 
.A1(n_2159),
.A2(n_2046),
.B(n_1934),
.C(n_2006),
.Y(n_2180)
);

NOR3x1_ASAP7_75t_L g2181 ( 
.A(n_2155),
.B(n_1968),
.C(n_1953),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2157),
.Y(n_2182)
);

AOI211xp5_ASAP7_75t_L g2183 ( 
.A1(n_2165),
.A2(n_2069),
.B(n_1988),
.C(n_1949),
.Y(n_2183)
);

NOR3x1_ASAP7_75t_L g2184 ( 
.A(n_2153),
.B(n_1965),
.C(n_1960),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2160),
.A2(n_2130),
.B(n_1962),
.Y(n_2185)
);

OAI21xp33_ASAP7_75t_L g2186 ( 
.A1(n_2179),
.A2(n_2160),
.B(n_2161),
.Y(n_2186)
);

NAND2x1_ASAP7_75t_L g2187 ( 
.A(n_2174),
.B(n_2162),
.Y(n_2187)
);

INVxp67_ASAP7_75t_SL g2188 ( 
.A(n_2175),
.Y(n_2188)
);

AND4x1_ASAP7_75t_L g2189 ( 
.A(n_2184),
.B(n_1928),
.C(n_2154),
.D(n_2166),
.Y(n_2189)
);

AOI211x1_ASAP7_75t_L g2190 ( 
.A1(n_2185),
.A2(n_2113),
.B(n_2032),
.C(n_2030),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2178),
.A2(n_2157),
.B(n_2156),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2170),
.Y(n_2192)
);

OAI21xp33_ASAP7_75t_L g2193 ( 
.A1(n_2178),
.A2(n_2075),
.B(n_2113),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_SL g2194 ( 
.A1(n_2172),
.A2(n_1886),
.B(n_2047),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2182),
.B(n_2183),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2181),
.B(n_2087),
.Y(n_2196)
);

AO22x2_ASAP7_75t_L g2197 ( 
.A1(n_2171),
.A2(n_1924),
.B1(n_1857),
.B2(n_1840),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2176),
.Y(n_2198)
);

OAI21xp33_ASAP7_75t_SL g2199 ( 
.A1(n_2173),
.A2(n_2097),
.B(n_2013),
.Y(n_2199)
);

NOR4xp25_ASAP7_75t_L g2200 ( 
.A(n_2188),
.B(n_2177),
.C(n_1913),
.D(n_1929),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2186),
.A2(n_1883),
.B(n_1886),
.Y(n_2201)
);

AO22x2_ASAP7_75t_L g2202 ( 
.A1(n_2198),
.A2(n_1867),
.B1(n_1840),
.B2(n_1844),
.Y(n_2202)
);

AOI21xp33_ASAP7_75t_L g2203 ( 
.A1(n_2192),
.A2(n_2180),
.B(n_1708),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2195),
.Y(n_2204)
);

AOI211xp5_ASAP7_75t_L g2205 ( 
.A1(n_2199),
.A2(n_1857),
.B(n_1874),
.C(n_1904),
.Y(n_2205)
);

OAI211xp5_ASAP7_75t_L g2206 ( 
.A1(n_2187),
.A2(n_1875),
.B(n_1892),
.C(n_1867),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2193),
.A2(n_2096),
.B(n_2086),
.C(n_2028),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2189),
.B(n_1843),
.Y(n_2208)
);

NAND5xp2_ASAP7_75t_L g2209 ( 
.A(n_2191),
.B(n_1883),
.C(n_1962),
.D(n_1681),
.E(n_1917),
.Y(n_2209)
);

AOI211xp5_ASAP7_75t_L g2210 ( 
.A1(n_2196),
.A2(n_2197),
.B(n_2190),
.C(n_2194),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2204),
.Y(n_2211)
);

NOR2xp67_ASAP7_75t_L g2212 ( 
.A(n_2206),
.B(n_2197),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2202),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2209),
.Y(n_2214)
);

NAND3xp33_ASAP7_75t_L g2215 ( 
.A(n_2201),
.B(n_1843),
.C(n_1766),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2208),
.A2(n_1970),
.B1(n_1991),
.B2(n_1983),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2200),
.A2(n_1991),
.B1(n_1983),
.B2(n_2096),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2207),
.B(n_1881),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_2211),
.B(n_2203),
.C(n_2210),
.Y(n_2219)
);

NAND4xp75_ASAP7_75t_L g2220 ( 
.A(n_2212),
.B(n_2202),
.C(n_2205),
.D(n_1847),
.Y(n_2220)
);

OAI221xp5_ASAP7_75t_SL g2221 ( 
.A1(n_2214),
.A2(n_2013),
.B1(n_1907),
.B2(n_1881),
.C(n_1891),
.Y(n_2221)
);

AOI221x1_ASAP7_75t_L g2222 ( 
.A1(n_2213),
.A2(n_2215),
.B1(n_2218),
.B2(n_2216),
.C(n_1907),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_SL g2223 ( 
.A1(n_2217),
.A2(n_1856),
.B(n_2013),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2219),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2222),
.B(n_1874),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_2220),
.Y(n_2226)
);

AOI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_2221),
.A2(n_1790),
.B(n_1866),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2224),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2225),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2229),
.Y(n_2230)
);

OAI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2228),
.A2(n_2226),
.B1(n_2227),
.B2(n_2223),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2230),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2231),
.A2(n_1925),
.B1(n_1858),
.B2(n_2016),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2232),
.Y(n_2234)
);

AO21x2_ASAP7_75t_L g2235 ( 
.A1(n_2234),
.A2(n_2233),
.B(n_2041),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2235),
.A2(n_1858),
.B1(n_1925),
.B2(n_1866),
.Y(n_2236)
);

OR2x6_ASAP7_75t_L g2237 ( 
.A(n_2236),
.B(n_1925),
.Y(n_2237)
);

AOI22xp33_ASAP7_75t_L g2238 ( 
.A1(n_2237),
.A2(n_1845),
.B1(n_1918),
.B2(n_1992),
.Y(n_2238)
);


endmodule