module fake_jpeg_13679_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_77),
.B1(n_80),
.B2(n_88),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_93),
.B1(n_20),
.B2(n_25),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_34),
.B1(n_19),
.B2(n_27),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_22),
.B(n_23),
.C(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_81),
.B(n_101),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_23),
.B1(n_52),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_23),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_40),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_20),
.B1(n_25),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_97),
.B1(n_35),
.B2(n_55),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_55),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_125),
.B1(n_140),
.B2(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_105),
.A2(n_86),
.B1(n_96),
.B2(n_100),
.Y(n_161)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_53),
.B1(n_39),
.B2(n_55),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_128),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_78),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_110),
.B(n_112),
.Y(n_177)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_42),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_44),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_64),
.C(n_46),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_115),
.C(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_121),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_126),
.Y(n_176)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_47),
.B1(n_57),
.B2(n_63),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_141),
.Y(n_143)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_56),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_37),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_74),
.B1(n_70),
.B2(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_139),
.Y(n_172)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_156),
.B1(n_171),
.B2(n_131),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_82),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_117),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_169),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_159),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_81),
.B(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_160),
.B(n_134),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_68),
.A3(n_70),
.B1(n_96),
.B2(n_100),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_107),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_97),
.B1(n_77),
.B2(n_91),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_91),
.B1(n_57),
.B2(n_47),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_161),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_125),
.C(n_109),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_101),
.B(n_71),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_76),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_103),
.A2(n_76),
.B1(n_45),
.B2(n_16),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_107),
.A2(n_49),
.B(n_38),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_137),
.B(n_138),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_178),
.A2(n_192),
.B(n_208),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_199),
.B1(n_209),
.B2(n_208),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_201),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_107),
.B1(n_130),
.B2(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_194),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_195),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_191),
.A2(n_202),
.B(n_178),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_128),
.B(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_127),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_126),
.B1(n_104),
.B2(n_123),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_204),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_152),
.B1(n_147),
.B2(n_146),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_124),
.B(n_108),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_49),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_38),
.B1(n_43),
.B2(n_62),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_207),
.B1(n_211),
.B2(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_171),
.B1(n_153),
.B2(n_151),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_145),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_1),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_145),
.B(n_3),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_174),
.Y(n_231)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_142),
.A3(n_175),
.B1(n_157),
.B2(n_145),
.C1(n_176),
.C2(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_219),
.B(n_226),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_240),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_160),
.B(n_150),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_215),
.B(n_163),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_201),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_181),
.A2(n_154),
.B1(n_173),
.B2(n_166),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_173),
.C(n_174),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_241),
.C(n_148),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_154),
.B1(n_173),
.B2(n_166),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_209),
.B1(n_198),
.B2(n_148),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_179),
.A2(n_162),
.B1(n_154),
.B2(n_170),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_244),
.B1(n_180),
.B2(n_205),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_203),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_170),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_200),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_245),
.A2(n_5),
.B(n_6),
.Y(n_280)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_274),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_268),
.C(n_270),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_202),
.B(n_192),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_280),
.B(n_217),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_221),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_261),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_256),
.A2(n_257),
.B1(n_264),
.B2(n_266),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_192),
.B1(n_182),
.B2(n_185),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_259),
.B(n_262),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_243),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_271),
.B(n_245),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_192),
.B1(n_206),
.B2(n_196),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_187),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_193),
.B1(n_190),
.B2(n_213),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_197),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_189),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_163),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_248),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_248),
.B1(n_230),
.B2(n_242),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_250),
.B1(n_228),
.B2(n_235),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_225),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_284),
.B(n_276),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_234),
.CI(n_222),
.CON(n_287),
.SN(n_287)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_290),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_298),
.B1(n_277),
.B2(n_260),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_301),
.B(n_280),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_292),
.A2(n_294),
.B1(n_260),
.B2(n_269),
.Y(n_326)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_230),
.B1(n_232),
.B2(n_236),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_265),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_257),
.A2(n_235),
.B1(n_232),
.B2(n_246),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_246),
.C(n_247),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_307),
.C(n_271),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_238),
.C(n_227),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_273),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_302),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_303),
.A2(n_267),
.B(n_258),
.C(n_279),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_217),
.Y(n_305)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_7),
.C(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_319),
.C(n_322),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_268),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_315),
.Y(n_336)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_266),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_282),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_253),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_325),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_317),
.A2(n_310),
.B1(n_321),
.B2(n_319),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_264),
.C(n_256),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_298),
.C(n_290),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_285),
.B(n_272),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_329),
.B(n_303),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_328),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_283),
.B(n_267),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_335),
.B(n_342),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_324),
.A2(n_291),
.B(n_305),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_300),
.C(n_304),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_339),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_300),
.C(n_304),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_322),
.A2(n_288),
.B(n_293),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_343),
.A2(n_338),
.B1(n_339),
.B2(n_345),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_292),
.C(n_288),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_346),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_326),
.B(n_313),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_344),
.A2(n_320),
.B(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_346),
.B1(n_296),
.B2(n_258),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_350),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_312),
.B(n_307),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_SL g351 ( 
.A(n_332),
.B(n_309),
.C(n_325),
.Y(n_351)
);

AOI21xp33_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_359),
.B(n_336),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_297),
.B1(n_296),
.B2(n_329),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_354),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_329),
.B(n_287),
.Y(n_356)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_340),
.B(n_287),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_340),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_297),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_329),
.C(n_289),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_342),
.C(n_330),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_366),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_336),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_370),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_360),
.A2(n_330),
.B1(n_337),
.B2(n_335),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_368),
.A2(n_362),
.B1(n_361),
.B2(n_363),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_369),
.B(n_8),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_346),
.B1(n_281),
.B2(n_10),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_281),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_365),
.A2(n_355),
.B(n_356),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_376),
.B(n_380),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_349),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_374),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_352),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_355),
.C(n_357),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_378),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_368),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_367),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_384),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_366),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_377),
.B(n_375),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_389),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_372),
.Y(n_390)
);

O2A1O1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_390),
.A2(n_382),
.B(n_9),
.C(n_10),
.Y(n_391)
);

AOI321xp33_ASAP7_75t_SL g393 ( 
.A1(n_391),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_392),
.B1(n_14),
.B2(n_13),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_387),
.B(n_13),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_14),
.Y(n_396)
);


endmodule