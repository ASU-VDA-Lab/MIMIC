module fake_ariane_2758_n_1806 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1806);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1806;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_22),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_9),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_98),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_67),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_115),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_0),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_54),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_71),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_104),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_38),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_8),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_50),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_33),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_155),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_163),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_97),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_50),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_47),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_73),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_20),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_29),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_26),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_2),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_93),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_70),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_59),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_62),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_88),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_126),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_160),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_69),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_87),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_9),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_141),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_112),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_56),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_11),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_24),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_72),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_177),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_57),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_30),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_78),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_39),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_66),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_180),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_82),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_106),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_164),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_179),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_60),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_153),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_173),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_86),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_43),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_53),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_51),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_132),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_27),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_129),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_134),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_127),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_27),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_6),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_31),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_39),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_43),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_3),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_48),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_168),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_42),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_5),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_7),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_79),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_40),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_84),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_140),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_25),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_124),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_2),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_8),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_108),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_46),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_30),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_89),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_0),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_176),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_101),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_40),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_122),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_165),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_14),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_52),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_14),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_159),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_85),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_46),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_49),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_19),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_121),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_110),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_45),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_41),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_156),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_149),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_118),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_133),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_37),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_166),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_123),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_105),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_81),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_38),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_10),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_247),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_247),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_247),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_269),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_269),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_269),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_269),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_269),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_233),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_192),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_192),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_223),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_304),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_314),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_299),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_210),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_320),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_322),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_299),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_362),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_213),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_207),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_182),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_210),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_190),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_216),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_213),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_220),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_287),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_244),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_212),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_186),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_186),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_212),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_188),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_361),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_361),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_215),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_231),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_217),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_236),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_266),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_232),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_246),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_280),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_290),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_298),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_234),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_240),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_242),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_302),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_243),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_245),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_254),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_233),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_270),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_303),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_259),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_262),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_256),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_392),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_364),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_408),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_379),
.A2(n_204),
.B1(n_307),
.B2(n_329),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_301),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_415),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_397),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_398),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_367),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_367),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_368),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_368),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_369),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_310),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_371),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_405),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_371),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_370),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_373),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_373),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_423),
.B(n_250),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_376),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_378),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_383),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_394),
.B(n_319),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_382),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_384),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_385),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_400),
.B(n_199),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_388),
.A2(n_317),
.B1(n_307),
.B2(n_308),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_387),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_403),
.B(n_277),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_449),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_433),
.A2(n_316),
.B1(n_317),
.B2(n_315),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_427),
.B(n_273),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_391),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_381),
.B(n_352),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_366),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_443),
.A2(n_321),
.B1(n_312),
.B2(n_270),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_418),
.B(n_250),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_389),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_477),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_461),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_521),
.B(n_405),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_530),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_467),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_521),
.B(n_430),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_512),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_512),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_422),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_470),
.B(n_399),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_512),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_512),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_493),
.A2(n_372),
.B1(n_426),
.B2(n_424),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_409),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_493),
.A2(n_420),
.B1(n_450),
.B2(n_416),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_477),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_493),
.B(n_411),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_458),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_467),
.B(n_429),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_467),
.B(n_434),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_514),
.B(n_439),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_517),
.B(n_440),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_515),
.B(n_441),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_390),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_484),
.B(n_436),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_460),
.B(n_444),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_447),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_484),
.B(n_448),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_453),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_520),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_460),
.B(n_454),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_493),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_484),
.B(n_425),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_460),
.B(n_183),
.Y(n_580)
);

AOI21x1_ASAP7_75t_L g581 ( 
.A1(n_465),
.A2(n_428),
.B(n_425),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_466),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_483),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_500),
.B(n_428),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_493),
.B(n_188),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

BUFx6f_ASAP7_75t_SL g589 ( 
.A(n_491),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_455),
.B(n_431),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_474),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_466),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_529),
.B(n_431),
.Y(n_593)
);

CKINVDCx6p67_ASAP7_75t_R g594 ( 
.A(n_464),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_492),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_477),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_530),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_492),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_478),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_479),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_495),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_481),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_481),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_482),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_509),
.B(n_183),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_491),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_468),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_482),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_504),
.B(n_506),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_516),
.B(n_432),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_489),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_491),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_508),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_432),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_455),
.B(n_435),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_480),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_480),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_480),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_529),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_516),
.B(n_435),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_473),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_526),
.B(n_437),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_528),
.B(n_533),
.C(n_532),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_480),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_495),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_501),
.Y(n_634)
);

HB1xp67_ASAP7_75t_SL g635 ( 
.A(n_531),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_522),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_523),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_486),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_469),
.A2(n_239),
.B1(n_329),
.B2(n_321),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_488),
.Y(n_643)
);

AO21x2_ASAP7_75t_L g644 ( 
.A1(n_509),
.A2(n_189),
.B(n_185),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_496),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_513),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_532),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_497),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_487),
.B(n_184),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_513),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_533),
.B(n_437),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_488),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_527),
.B(n_438),
.Y(n_654)
);

BUFx6f_ASAP7_75t_SL g655 ( 
.A(n_513),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_490),
.B(n_438),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_490),
.B(n_442),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_505),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_513),
.Y(n_659)
);

BUFx6f_ASAP7_75t_SL g660 ( 
.A(n_518),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_505),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_510),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_523),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_510),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_518),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_L g666 ( 
.A(n_494),
.B(n_203),
.C(n_201),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_518),
.Y(n_667)
);

NOR2x1p5_ASAP7_75t_L g668 ( 
.A(n_457),
.B(n_308),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_494),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_518),
.B(n_184),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_498),
.B(n_442),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_518),
.Y(n_672)
);

NOR2x1p5_ASAP7_75t_L g673 ( 
.A(n_457),
.B(n_309),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_459),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_524),
.Y(n_675)
);

AND2x6_ASAP7_75t_L g676 ( 
.A(n_498),
.B(n_200),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_499),
.B(n_445),
.Y(n_677)
);

BUFx8_ASAP7_75t_SL g678 ( 
.A(n_457),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_503),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_568),
.B(n_393),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_616),
.B(n_499),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_616),
.B(n_264),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_549),
.B(n_193),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_585),
.B(n_502),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_619),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_539),
.A2(n_256),
.B1(n_265),
.B2(n_360),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_539),
.A2(n_561),
.B1(n_550),
.B2(n_644),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_502),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_537),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_593),
.B(n_507),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_617),
.B(n_507),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_451),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_644),
.A2(n_525),
.B1(n_511),
.B2(n_524),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_548),
.B(n_193),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_611),
.B(n_445),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_535),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_617),
.B(n_511),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_556),
.B(n_196),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_540),
.B(n_525),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_589),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_558),
.B(n_566),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_543),
.B(n_271),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_628),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_642),
.A2(n_235),
.B(n_297),
.C(n_230),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_644),
.A2(n_265),
.B1(n_198),
.B2(n_325),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_535),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_544),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_547),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_538),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_547),
.B(n_196),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_540),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_639),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_571),
.B(n_197),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_568),
.B(n_446),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_573),
.B(n_197),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_589),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_567),
.B(n_198),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_541),
.B(n_457),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_639),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_541),
.B(n_476),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_567),
.B(n_205),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_647),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_553),
.B(n_205),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_591),
.B(n_206),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_547),
.B(n_206),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_547),
.B(n_208),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_545),
.B(n_476),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_562),
.B(n_272),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_546),
.B(n_476),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_647),
.B(n_476),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_553),
.B(n_208),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

INVxp33_ASAP7_75t_L g735 ( 
.A(n_636),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_538),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_554),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_642),
.A2(n_226),
.B(n_221),
.C(n_238),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_652),
.B(n_194),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_536),
.B(n_278),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_606),
.A2(n_357),
.B1(n_328),
.B2(n_325),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_652),
.B(n_268),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_625),
.B(n_285),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_625),
.B(n_318),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_557),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_557),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_570),
.B(n_283),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_656),
.B(n_318),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_671),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_577),
.B(n_580),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_635),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_600),
.B(n_328),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_649),
.B(n_289),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_563),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_579),
.B(n_291),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_563),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_600),
.B(n_446),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_559),
.A2(n_218),
.B(n_209),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_609),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_677),
.B(n_333),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_613),
.B(n_292),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_634),
.B(n_452),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_565),
.B(n_572),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_587),
.B(n_333),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_613),
.B(n_335),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_578),
.B(n_587),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_634),
.B(n_452),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_355),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_615),
.B(n_355),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_569),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_612),
.B(n_404),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_654),
.B(n_357),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_613),
.B(n_341),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_569),
.Y(n_774)
);

AND2x4_ASAP7_75t_SL g775 ( 
.A(n_627),
.B(n_311),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_404),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_590),
.B(n_621),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_629),
.B(n_360),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_582),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_565),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_542),
.B(n_459),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_578),
.B(n_248),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_572),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_582),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_542),
.B(n_471),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_575),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_578),
.B(n_258),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_578),
.B(n_263),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_344),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_614),
.B(n_312),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_612),
.A2(n_471),
.B1(n_475),
.B2(n_472),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_668),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_592),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_614),
.B(n_326),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_575),
.B(n_472),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_R g796 ( 
.A(n_594),
.B(n_332),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_576),
.B(n_475),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_576),
.B(n_345),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_612),
.B(n_410),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_640),
.A2(n_414),
.B1(n_413),
.B2(n_412),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_594),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_631),
.B(n_350),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_592),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_631),
.B(n_332),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_598),
.B(n_356),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_612),
.B(n_356),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_626),
.B(n_410),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_598),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_666),
.B(n_537),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_674),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_674),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_583),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_601),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_668),
.A2(n_267),
.B1(n_284),
.B2(n_305),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_601),
.B(n_219),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_603),
.B(n_222),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_603),
.B(n_224),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_604),
.B(n_225),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_604),
.B(n_228),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_672),
.B(n_323),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_666),
.B(n_188),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_537),
.B(n_202),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_673),
.A2(n_331),
.B1(n_343),
.B2(n_348),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_537),
.B(n_351),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_584),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_537),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_672),
.B(n_354),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_673),
.B(n_412),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_560),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_586),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_626),
.B(n_413),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_605),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_626),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_626),
.B(n_414),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_597),
.B(n_607),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_804),
.A2(n_630),
.B(n_605),
.C(n_610),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_800),
.A2(n_663),
.B1(n_640),
.B2(n_626),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_696),
.B(n_749),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_685),
.B(n_597),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_682),
.B(n_657),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_710),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_697),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_707),
.Y(n_843)
);

OR2x4_ASAP7_75t_L g844 ( 
.A(n_790),
.B(n_806),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_701),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_708),
.Y(n_847)
);

INVx6_ASAP7_75t_L g848 ( 
.A(n_701),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_801),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_693),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_709),
.B(n_676),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_833),
.B(n_597),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_682),
.B(n_610),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_833),
.B(n_597),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_710),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_SL g856 ( 
.A(n_725),
.B(n_670),
.C(n_641),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_763),
.A2(n_574),
.B(n_552),
.Y(n_857)
);

AOI21xp33_ASAP7_75t_L g858 ( 
.A1(n_703),
.A2(n_641),
.B(n_630),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_834),
.B(n_643),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_715),
.B(n_643),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_800),
.A2(n_676),
.B1(n_653),
.B2(n_669),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_762),
.B(n_417),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_736),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_767),
.B(n_417),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_734),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_737),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_745),
.A2(n_669),
.B1(n_560),
.B2(n_596),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_834),
.B(n_597),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_746),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_680),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_804),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_739),
.B(n_676),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_742),
.B(n_676),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_774),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_688),
.B(n_676),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_759),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_755),
.B(n_676),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_829),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_796),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_796),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_776),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_751),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_717),
.B(n_607),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_779),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_755),
.B(n_676),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_784),
.A2(n_632),
.B1(n_534),
.B2(n_624),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_775),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_717),
.B(n_665),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_751),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_701),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_720),
.B(n_665),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_690),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_799),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_690),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_735),
.B(n_672),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_720),
.B(n_607),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_754),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_829),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_800),
.A2(n_651),
.B1(n_602),
.B2(n_675),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_687),
.B(n_607),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_771),
.A2(n_651),
.B1(n_602),
.B2(n_675),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_793),
.Y(n_903)
);

OR2x2_ASAP7_75t_SL g904 ( 
.A(n_807),
.B(n_678),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_684),
.B(n_586),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_750),
.A2(n_623),
.B(n_596),
.C(n_555),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_771),
.A2(n_655),
.B1(n_659),
.B2(n_660),
.Y(n_907)
);

AND3x1_ASAP7_75t_SL g908 ( 
.A(n_803),
.B(n_813),
.C(n_808),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_690),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_SL g910 ( 
.A(n_703),
.B(n_358),
.C(n_359),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_690),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_832),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_704),
.B(n_607),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_756),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_736),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_681),
.B(n_588),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_831),
.A2(n_599),
.B1(n_633),
.B2(n_664),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_702),
.B(n_588),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_748),
.B(n_595),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_760),
.B(n_595),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_780),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_713),
.B(n_599),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_783),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_786),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_812),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_828),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_826),
.Y(n_927)
);

AND2x6_ASAP7_75t_SL g928 ( 
.A(n_730),
.B(n_1),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_831),
.B(n_667),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_689),
.A2(n_534),
.B(n_564),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_831),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_691),
.A2(n_662),
.B(n_664),
.C(n_661),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_828),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_721),
.B(n_618),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_706),
.A2(n_633),
.B1(n_638),
.B2(n_662),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_792),
.B(n_667),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_724),
.B(n_777),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_712),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_750),
.B(n_618),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_743),
.B(n_618),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_726),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_805),
.B(n_638),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_778),
.B(n_645),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_718),
.B(n_534),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_692),
.A2(n_632),
.B1(n_551),
.B2(n_555),
.Y(n_945)
);

AND3x2_ASAP7_75t_SL g946 ( 
.A(n_810),
.B(n_661),
.C(n_658),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_712),
.B(n_761),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_SL g948 ( 
.A(n_814),
.B(n_823),
.C(n_730),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_698),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_761),
.B(n_645),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_740),
.B(n_581),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_747),
.B(n_618),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_747),
.B(n_618),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_765),
.B(n_648),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_815),
.A2(n_632),
.B1(n_551),
.B2(n_564),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_765),
.B(n_648),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_825),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_744),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_752),
.Y(n_959)
);

INVxp67_ASAP7_75t_SL g960 ( 
.A(n_826),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_773),
.B(n_679),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_826),
.B(n_564),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_789),
.B(n_811),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_SL g964 ( 
.A1(n_753),
.A2(n_227),
.B1(n_202),
.B2(n_276),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_794),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_830),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_723),
.B(n_596),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_789),
.B(n_679),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_740),
.B(n_581),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_732),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_733),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_826),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_795),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_797),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_700),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_835),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_SL g977 ( 
.A1(n_787),
.A2(n_227),
.B1(n_202),
.B2(n_274),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_791),
.B(n_622),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_781),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_791),
.B(n_622),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_785),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_SL g982 ( 
.A(n_683),
.B(n_347),
.C(n_260),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_686),
.B(n_622),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_714),
.B(n_338),
.C(n_257),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_835),
.B(n_623),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_798),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_719),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_772),
.B(n_623),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_722),
.Y(n_989)
);

AND2x6_ASAP7_75t_L g990 ( 
.A(n_709),
.B(n_679),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_695),
.A2(n_660),
.B1(n_659),
.B2(n_655),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_729),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_731),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_809),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_716),
.B(n_624),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_802),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_768),
.B(n_624),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_820),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_816),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_769),
.B(n_679),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_637),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_817),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_741),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_820),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_782),
.B(n_637),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_925),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_845),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_849),
.B(n_827),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_948),
.A2(n_738),
.B(n_705),
.C(n_758),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_947),
.A2(n_766),
.B(n_764),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_842),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_838),
.B(n_818),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_998),
.A2(n_819),
.B1(n_699),
.B2(n_766),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1004),
.A2(n_711),
.B1(n_728),
.B2(n_727),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_727),
.B(n_711),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_846),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_949),
.B(n_694),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_948),
.A2(n_822),
.B1(n_728),
.B2(n_787),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_949),
.B(n_694),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_871),
.B(n_824),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_862),
.B(n_646),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_877),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_837),
.A2(n_824),
.B(n_788),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_840),
.A2(n_650),
.B(n_646),
.C(n_782),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_871),
.B(n_679),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_893),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_910),
.A2(n_650),
.B(n_646),
.C(n_788),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_910),
.A2(n_650),
.B(n_503),
.C(n_237),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_843),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_846),
.B(n_787),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_SL g1031 ( 
.A(n_888),
.Y(n_1031)
);

AND2x4_ASAP7_75t_SL g1032 ( 
.A(n_846),
.B(n_227),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_961),
.A2(n_660),
.B(n_659),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_853),
.A2(n_10),
.B(n_11),
.C(n_16),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_864),
.B(n_787),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_938),
.A2(n_620),
.B1(n_655),
.B2(n_229),
.Y(n_1036)
);

AND2x2_ASAP7_75t_SL g1037 ( 
.A(n_837),
.B(n_787),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_858),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_857),
.A2(n_938),
.B(n_886),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_860),
.B(n_620),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_878),
.A2(n_620),
.B(n_709),
.C(n_503),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_893),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_857),
.A2(n_709),
.B(n_282),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_882),
.B(n_620),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_847),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_848),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_968),
.A2(n_709),
.B(n_503),
.C(n_22),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_950),
.A2(n_709),
.B(n_286),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_941),
.B(n_249),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_848),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_877),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_863),
.A2(n_281),
.B1(n_353),
.B2(n_337),
.Y(n_1052)
);

AO32x2_ASAP7_75t_L g1053 ( 
.A1(n_867),
.A2(n_503),
.A3(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_954),
.A2(n_279),
.B(n_334),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_863),
.A2(n_915),
.B1(n_963),
.B2(n_975),
.Y(n_1055)
);

BUFx8_ASAP7_75t_L g1056 ( 
.A(n_850),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_999),
.A2(n_18),
.B(n_21),
.C(n_23),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_956),
.A2(n_275),
.B(n_296),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_894),
.B(n_1003),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_848),
.B(n_503),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_929),
.B(n_28),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_880),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_883),
.B(n_295),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_926),
.B(n_29),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_893),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_890),
.B(n_294),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_870),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_881),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_844),
.B(n_293),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_933),
.B(n_971),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_964),
.A2(n_856),
.B(n_982),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_915),
.A2(n_288),
.B(n_261),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_895),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_865),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_859),
.A2(n_255),
.B1(n_253),
.B2(n_252),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_SL g1076 ( 
.A1(n_944),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_SL g1077 ( 
.A1(n_952),
.A2(n_251),
.B(n_34),
.C(n_41),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_861),
.A2(n_32),
.B1(n_44),
.B2(n_47),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_866),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_859),
.B(n_44),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_1002),
.A2(n_48),
.B(n_51),
.C(n_58),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_SL g1082 ( 
.A1(n_967),
.A2(n_930),
.B(n_995),
.C(n_1001),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_859),
.B(n_65),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_959),
.B(n_896),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_895),
.Y(n_1085)
);

BUFx8_ASAP7_75t_SL g1086 ( 
.A(n_891),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_929),
.B(n_76),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_859),
.B(n_77),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_844),
.B(n_80),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_905),
.A2(n_988),
.B(n_1000),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_958),
.B(n_90),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_859),
.B(n_996),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_997),
.A2(n_91),
.B(n_92),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_937),
.B(n_96),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_931),
.A2(n_102),
.B1(n_109),
.B2(n_111),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_869),
.B(n_114),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_836),
.A2(n_116),
.B(n_117),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_904),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_907),
.B(n_120),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_895),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_931),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_874),
.B(n_128),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_965),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_906),
.A2(n_131),
.B(n_137),
.C(n_154),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_889),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_875),
.B(n_157),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_872),
.A2(n_158),
.B(n_169),
.C(n_170),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_885),
.B(n_171),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_951),
.A2(n_174),
.B(n_969),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_861),
.A2(n_912),
.B1(n_903),
.B2(n_902),
.Y(n_1110)
);

AO32x1_ASAP7_75t_L g1111 ( 
.A1(n_955),
.A2(n_945),
.A3(n_994),
.B1(n_887),
.B2(n_992),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_873),
.A2(n_964),
.B(n_856),
.C(n_986),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_909),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_936),
.B(n_900),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_868),
.B(n_841),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_973),
.B(n_974),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_841),
.B(n_855),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_876),
.A2(n_983),
.B(n_932),
.C(n_919),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_980),
.B(n_970),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_980),
.B(n_916),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_932),
.A2(n_942),
.B(n_993),
.C(n_989),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_892),
.B(n_936),
.Y(n_1122)
);

CKINVDCx8_ASAP7_75t_R g1123 ( 
.A(n_928),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_892),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_914),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_902),
.A2(n_917),
.B1(n_899),
.B2(n_879),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_839),
.A2(n_943),
.B(n_920),
.C(n_982),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_898),
.Y(n_1128)
);

AO32x1_ASAP7_75t_L g1129 ( 
.A1(n_979),
.A2(n_987),
.A3(n_981),
.B1(n_908),
.B2(n_921),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_960),
.A2(n_953),
.B(n_940),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_977),
.A2(n_918),
.B(n_984),
.C(n_978),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_909),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_991),
.A2(n_976),
.B1(n_899),
.B2(n_855),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_977),
.A2(n_984),
.B(n_939),
.C(n_917),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_900),
.A2(n_960),
.B(n_879),
.C(n_924),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_923),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_976),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_852),
.B(n_854),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_957),
.B(n_966),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_927),
.B(n_972),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_985),
.A2(n_934),
.B(n_913),
.C(n_901),
.Y(n_1141)
);

INVxp33_ASAP7_75t_SL g1142 ( 
.A(n_884),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_927),
.B(n_972),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_976),
.B(n_911),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_922),
.A2(n_897),
.B(n_946),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_985),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_935),
.B(n_946),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1132),
.Y(n_1148)
);

AOI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_1037),
.A2(n_935),
.B(n_1005),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1059),
.A2(n_1005),
.B1(n_911),
.B2(n_990),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1109),
.A2(n_1009),
.B(n_1118),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1145),
.A2(n_990),
.B(n_962),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1007),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1015),
.A2(n_990),
.B(n_962),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1011),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1046),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1120),
.B(n_927),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1006),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1086),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1055),
.A2(n_972),
.B(n_990),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1010),
.A2(n_1043),
.B(n_1048),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1056),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1013),
.A2(n_1012),
.B(n_1111),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1071),
.A2(n_1078),
.B(n_1038),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_SL g1165 ( 
.A(n_1062),
.B(n_1123),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1056),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1121),
.A2(n_1014),
.B(n_1131),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1111),
.A2(n_1082),
.B(n_1094),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1029),
.Y(n_1169)
);

NOR4xp25_ASAP7_75t_L g1170 ( 
.A(n_1034),
.B(n_1057),
.C(n_1134),
.D(n_1112),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1111),
.A2(n_1097),
.B(n_1024),
.Y(n_1171)
);

AOI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1018),
.A2(n_1023),
.B(n_1127),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1116),
.B(n_1022),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1093),
.A2(n_1106),
.B(n_1102),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1051),
.B(n_1008),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1130),
.A2(n_1033),
.B(n_1141),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_1095),
.A2(n_1110),
.B1(n_1028),
.B2(n_1135),
.C(n_1126),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1119),
.B(n_1017),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1021),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1096),
.A2(n_1108),
.B(n_1133),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1124),
.B(n_1067),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1061),
.B(n_1101),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_1068),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1104),
.A2(n_1146),
.B(n_1025),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1092),
.A2(n_1099),
.B(n_1143),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1061),
.A2(n_1079),
.B1(n_1045),
.B2(n_1074),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1098),
.B(n_1016),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1084),
.B(n_1105),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1140),
.A2(n_1088),
.B(n_1083),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1103),
.B(n_1064),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1046),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1087),
.A2(n_1035),
.B(n_1091),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_SL g1193 ( 
.A1(n_1080),
.A2(n_1044),
.B(n_1040),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1122),
.B(n_1087),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1036),
.A2(n_1027),
.B(n_1117),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1107),
.A2(n_1054),
.B(n_1058),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1100),
.B(n_1042),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1019),
.B(n_1114),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1139),
.A2(n_1081),
.B(n_1144),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1020),
.A2(n_1060),
.B1(n_1115),
.B2(n_1075),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1046),
.B(n_1030),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_SL g1202 ( 
.A1(n_1125),
.A2(n_1049),
.B(n_1070),
.C(n_1136),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1032),
.B(n_1050),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1132),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1089),
.A2(n_1069),
.B1(n_1137),
.B2(n_1138),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1072),
.A2(n_1076),
.B(n_1052),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1129),
.A2(n_1142),
.B(n_1113),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1030),
.B(n_1073),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1128),
.B(n_1065),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1053),
.A2(n_1129),
.B(n_1065),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1073),
.A2(n_1085),
.B(n_1113),
.C(n_1053),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1053),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1031),
.A2(n_1037),
.B1(n_837),
.B2(n_948),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1031),
.A2(n_1039),
.B(n_1041),
.Y(n_1215)
);

O2A1O1Ixp5_ASAP7_75t_L g1216 ( 
.A1(n_1109),
.A2(n_1009),
.B(n_886),
.C(n_878),
.Y(n_1216)
);

AOI221x1_ASAP7_75t_L g1217 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1009),
.B2(n_910),
.C(n_1078),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1122),
.B(n_1105),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1056),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1071),
.A2(n_948),
.B(n_910),
.C(n_1109),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1060),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1109),
.A2(n_836),
.B(n_878),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1118),
.A2(n_1039),
.A3(n_1135),
.B(n_876),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1120),
.B(n_998),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1230)
);

AOI221x1_ASAP7_75t_L g1231 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1009),
.B2(n_910),
.C(n_1078),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1080),
.A2(n_853),
.B(n_840),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_SL g1234 ( 
.A1(n_1127),
.A2(n_1080),
.B(n_1141),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1009),
.B(n_964),
.C(n_1071),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1059),
.B(n_553),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1120),
.B(n_998),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1037),
.A2(n_1071),
.B(n_1109),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1007),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1120),
.B(n_998),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1071),
.A2(n_948),
.B(n_910),
.C(n_1109),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1007),
.B(n_757),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1059),
.B(n_553),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1011),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1122),
.B(n_1105),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1056),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1109),
.A2(n_836),
.B(n_878),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1120),
.B(n_998),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1037),
.A2(n_838),
.B1(n_1004),
.B2(n_998),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1011),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1022),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1007),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1132),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1132),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1090),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1007),
.B(n_757),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1120),
.B(n_998),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1120),
.B(n_998),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1059),
.B(n_553),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1056),
.Y(n_1270)
);

BUFx4_ASAP7_75t_SL g1271 ( 
.A(n_1098),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1109),
.A2(n_836),
.B(n_878),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1007),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1120),
.B(n_998),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1087),
.B(n_929),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1086),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1122),
.B(n_1105),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1109),
.A2(n_836),
.B(n_878),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1109),
.A2(n_836),
.B(n_878),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1039),
.A2(n_947),
.B(n_851),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1059),
.B(n_553),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1225),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1155),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1214),
.A2(n_1235),
.B1(n_1238),
.B2(n_1252),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1171),
.B(n_1220),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_SL g1287 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1238),
.C(n_1151),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1164),
.A2(n_1170),
.B1(n_1151),
.B2(n_1252),
.C(n_1167),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1169),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1194),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1224),
.A2(n_1253),
.B(n_1242),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1218),
.A2(n_1226),
.B(n_1222),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1255),
.A2(n_1263),
.B(n_1261),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1219),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1225),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1236),
.A2(n_1269),
.B1(n_1281),
.B2(n_1245),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1186),
.A2(n_1231),
.B(n_1217),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1298)
);

OAI211xp5_ASAP7_75t_L g1299 ( 
.A1(n_1167),
.A2(n_1164),
.B(n_1170),
.C(n_1172),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1230),
.A2(n_1280),
.B(n_1232),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1240),
.A2(n_1246),
.B(n_1268),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1259),
.A2(n_1260),
.B(n_1266),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1172),
.A2(n_1251),
.B1(n_1229),
.B2(n_1274),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1186),
.B(n_1200),
.Y(n_1304)
);

NAND2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1159),
.B(n_1175),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1256),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1279),
.A2(n_1278),
.B(n_1250),
.C(n_1272),
.Y(n_1307)
);

INVxp33_ASAP7_75t_L g1308 ( 
.A(n_1173),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1163),
.A2(n_1180),
.B(n_1278),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_1161),
.B(n_1212),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1200),
.B(n_1229),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1227),
.A2(n_1279),
.B(n_1250),
.C(n_1272),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1153),
.B(n_1239),
.Y(n_1313)
);

OAI21xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1192),
.A2(n_1150),
.B(n_1227),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1215),
.A2(n_1176),
.B(n_1216),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1154),
.A2(n_1152),
.B(n_1174),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1149),
.A2(n_1195),
.B(n_1274),
.C(n_1237),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1189),
.A2(n_1184),
.B(n_1160),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1211),
.A2(n_1149),
.B(n_1179),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1208),
.B(n_1201),
.Y(n_1320)
);

INVx3_ASAP7_75t_SL g1321 ( 
.A(n_1276),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1271),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1237),
.A2(n_1265),
.B1(n_1267),
.B2(n_1251),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1193),
.A2(n_1233),
.B(n_1185),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1247),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1241),
.B(n_1265),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1201),
.B(n_1225),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1234),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1183),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1275),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1254),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1179),
.A2(n_1199),
.B(n_1213),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1162),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1275),
.B(n_1157),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1206),
.A2(n_1196),
.B(n_1241),
.Y(n_1335)
);

CKINVDCx6p67_ASAP7_75t_R g1336 ( 
.A(n_1166),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1209),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1267),
.A2(n_1206),
.B(n_1202),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1157),
.B(n_1188),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1210),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1210),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1147),
.A2(n_1225),
.B(n_1197),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1228),
.B(n_1273),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1187),
.A2(n_1228),
.B(n_1203),
.Y(n_1344)
);

AOI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1257),
.A2(n_1181),
.B(n_1190),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1156),
.Y(n_1346)
);

INVx8_ASAP7_75t_L g1347 ( 
.A(n_1219),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1248),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1228),
.B(n_1277),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1221),
.B(n_1249),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1191),
.A2(n_1148),
.B(n_1258),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1204),
.B(n_1258),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1262),
.A2(n_1270),
.B(n_1165),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1262),
.A2(n_837),
.B1(n_1037),
.B2(n_948),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1220),
.A2(n_1242),
.B(n_1224),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1151),
.A2(n_1167),
.B(n_1234),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1235),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1214),
.A2(n_837),
.B1(n_1037),
.B2(n_948),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_SL g1359 ( 
.A1(n_1151),
.A2(n_1167),
.B(n_1234),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1168),
.A2(n_1171),
.A3(n_1211),
.B(n_1177),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1192),
.B(n_1186),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1223),
.A2(n_1243),
.B1(n_1235),
.B2(n_1214),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1168),
.A2(n_1171),
.A3(n_1211),
.B(n_1177),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1168),
.A2(n_1171),
.B(n_1220),
.Y(n_1364)
);

O2A1O1Ixp5_ASAP7_75t_L g1365 ( 
.A1(n_1151),
.A2(n_1223),
.B(n_1243),
.C(n_1167),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1155),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1218),
.A2(n_1226),
.B(n_1222),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1223),
.A2(n_1243),
.B1(n_1235),
.B2(n_1214),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1168),
.A2(n_1171),
.A3(n_1211),
.B(n_1177),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1155),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1236),
.B(n_640),
.Y(n_1371)
);

INVx4_ASAP7_75t_SL g1372 ( 
.A(n_1194),
.Y(n_1372)
);

AOI222xp33_ASAP7_75t_L g1373 ( 
.A1(n_1214),
.A2(n_837),
.B1(n_948),
.B2(n_833),
.C1(n_640),
.C2(n_663),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1223),
.A2(n_1243),
.B1(n_1235),
.B2(n_1214),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1155),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_R g1376 ( 
.A(n_1167),
.B(n_1151),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1220),
.A2(n_1242),
.B(n_1224),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1182),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1220),
.A2(n_1242),
.B(n_1224),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1236),
.B(n_640),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1158),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1155),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1276),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1235),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1220),
.A2(n_1242),
.B(n_1224),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_SL g1387 ( 
.A(n_1223),
.B(n_1243),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1168),
.A2(n_1171),
.A3(n_1211),
.B(n_1177),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1235),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1148),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_R g1391 ( 
.A(n_1167),
.B(n_1151),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1182),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1155),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1244),
.B(n_1264),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1194),
.B(n_1208),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1183),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1225),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1214),
.A2(n_837),
.B1(n_1037),
.B2(n_948),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1387),
.A2(n_1312),
.B(n_1307),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1288),
.A2(n_1299),
.B1(n_1399),
.B2(n_1358),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1313),
.B(n_1393),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1283),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1289),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1291),
.A2(n_1355),
.B(n_1293),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1362),
.A2(n_1374),
.B(n_1368),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1387),
.A2(n_1374),
.B1(n_1368),
.B2(n_1362),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1395),
.B(n_1308),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1307),
.A2(n_1312),
.B(n_1287),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1308),
.B(n_1326),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_L g1411 ( 
.A(n_1321),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1357),
.A2(n_1385),
.B(n_1389),
.C(n_1287),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1357),
.A2(n_1389),
.B(n_1385),
.C(n_1365),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1361),
.A2(n_1288),
.B(n_1304),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1326),
.B(n_1311),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1306),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1311),
.B(n_1286),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1304),
.B(n_1345),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1383),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1299),
.A2(n_1380),
.B(n_1371),
.C(n_1356),
.Y(n_1420)
);

O2A1O1Ixp5_ASAP7_75t_L g1421 ( 
.A1(n_1338),
.A2(n_1328),
.B(n_1317),
.C(n_1343),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1345),
.B(n_1348),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1314),
.A2(n_1371),
.B(n_1380),
.C(n_1358),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1292),
.A2(n_1302),
.B(n_1367),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_SL g1425 ( 
.A1(n_1352),
.A2(n_1350),
.B(n_1343),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1399),
.A2(n_1284),
.B1(n_1354),
.B2(n_1303),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1284),
.A2(n_1354),
.B1(n_1303),
.B2(n_1297),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1296),
.A2(n_1376),
.B1(n_1391),
.B2(n_1317),
.Y(n_1428)
);

CKINVDCx16_ASAP7_75t_R g1429 ( 
.A(n_1322),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1333),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1376),
.A2(n_1391),
.B1(n_1323),
.B2(n_1384),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1323),
.B(n_1286),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1372),
.B(n_1327),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1298),
.B(n_1384),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1298),
.B(n_1392),
.Y(n_1435)
);

O2A1O1Ixp5_ASAP7_75t_L g1436 ( 
.A1(n_1338),
.A2(n_1349),
.B(n_1342),
.C(n_1305),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1377),
.A2(n_1379),
.B(n_1386),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1327),
.B(n_1396),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1321),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1325),
.B(n_1331),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_1382),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1394),
.B(n_1396),
.Y(n_1443)
);

BUFx2_ASAP7_75t_R g1444 ( 
.A(n_1329),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1359),
.A2(n_1373),
.B(n_1309),
.C(n_1310),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1337),
.B(n_1346),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1344),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1337),
.B(n_1336),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1373),
.A2(n_1335),
.B1(n_1310),
.B2(n_1319),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1332),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1341),
.B(n_1340),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_1282),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1319),
.A2(n_1334),
.B1(n_1330),
.B2(n_1339),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1334),
.A2(n_1330),
.B1(n_1290),
.B2(n_1390),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1390),
.B(n_1294),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1367),
.A2(n_1300),
.B(n_1301),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1316),
.A2(n_1318),
.B(n_1324),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1309),
.B(n_1360),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1347),
.A2(n_1282),
.B1(n_1397),
.B2(n_1295),
.Y(n_1460)
);

NOR2xp67_ASAP7_75t_L g1461 ( 
.A(n_1320),
.B(n_1381),
.Y(n_1461)
);

BUFx2_ASAP7_75t_SL g1462 ( 
.A(n_1333),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1353),
.B(n_1351),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1315),
.A2(n_1285),
.B(n_1364),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1363),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1369),
.B(n_1388),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1315),
.Y(n_1467)
);

O2A1O1Ixp5_ASAP7_75t_L g1468 ( 
.A1(n_1398),
.A2(n_1365),
.B(n_1385),
.C(n_1357),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1333),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1387),
.A2(n_1243),
.B(n_1223),
.C(n_1357),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1323),
.B(n_1311),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1291),
.A2(n_1355),
.B(n_1293),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1323),
.B(n_1311),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1288),
.A2(n_1299),
.B1(n_1399),
.B2(n_1358),
.Y(n_1474)
);

O2A1O1Ixp5_ASAP7_75t_L g1475 ( 
.A1(n_1365),
.A2(n_1385),
.B(n_1389),
.C(n_1357),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1323),
.B(n_1311),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1313),
.B(n_1378),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1387),
.A2(n_1151),
.B(n_1307),
.Y(n_1478)
);

O2A1O1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1387),
.A2(n_1243),
.B(n_1223),
.C(n_1357),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1387),
.A2(n_1151),
.B(n_1307),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1383),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1313),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1288),
.A2(n_1299),
.B1(n_1399),
.B2(n_1358),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_SL g1484 ( 
.A(n_1333),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1288),
.A2(n_1299),
.B1(n_1399),
.B2(n_1358),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1288),
.A2(n_1299),
.B1(n_1399),
.B2(n_1358),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1467),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1471),
.B(n_1473),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1403),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1405),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1439),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1405),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1437),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1404),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1466),
.B(n_1451),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1471),
.B(n_1473),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1459),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1464),
.A2(n_1424),
.B(n_1421),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1436),
.A2(n_1409),
.B(n_1480),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1441),
.B(n_1442),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1452),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1482),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1458),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1450),
.A2(n_1427),
.B(n_1445),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1432),
.B(n_1415),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1428),
.B(n_1478),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1452),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1432),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1417),
.B(n_1431),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1472),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1407),
.A2(n_1486),
.B1(n_1485),
.B2(n_1401),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1470),
.A2(n_1479),
.B1(n_1406),
.B2(n_1401),
.C(n_1483),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1427),
.A2(n_1400),
.B(n_1426),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1463),
.B(n_1453),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1447),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1431),
.B(n_1402),
.Y(n_1520)
);

AO21x2_ASAP7_75t_L g1521 ( 
.A1(n_1426),
.A2(n_1428),
.B(n_1485),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1416),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1425),
.A2(n_1454),
.B(n_1460),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1484),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1474),
.A2(n_1486),
.B(n_1483),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1477),
.B(n_1410),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1422),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1414),
.B(n_1443),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1413),
.B(n_1412),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1474),
.A2(n_1454),
.B(n_1423),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1408),
.B(n_1435),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1434),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1446),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1488),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1488),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1487),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1521),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1429),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1526),
.A2(n_1462),
.B1(n_1420),
.B2(n_1438),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1491),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1518),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1494),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1496),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1522),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1514),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1498),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1508),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_1449),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1526),
.A2(n_1438),
.B1(n_1433),
.B2(n_1461),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1506),
.Y(n_1555)
);

AOI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1509),
.A2(n_1455),
.B(n_1460),
.C(n_1456),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1493),
.B(n_1411),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1455),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1519),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1495),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1553),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1545),
.B(n_1497),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1553),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1541),
.A2(n_1521),
.B1(n_1526),
.B2(n_1516),
.C(n_1515),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1535),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1541),
.A2(n_1521),
.B1(n_1526),
.B2(n_1517),
.Y(n_1568)
);

NOR5xp2_ASAP7_75t_SL g1569 ( 
.A(n_1549),
.B(n_1516),
.C(n_1530),
.D(n_1521),
.E(n_1526),
.Y(n_1569)
);

OAI33xp33_ASAP7_75t_L g1570 ( 
.A1(n_1552),
.A2(n_1513),
.A3(n_1524),
.B1(n_1533),
.B2(n_1511),
.B3(n_1532),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1541),
.A2(n_1513),
.B1(n_1520),
.B2(n_1521),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1541),
.A2(n_1520),
.B1(n_1502),
.B2(n_1517),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1541),
.A2(n_1520),
.B1(n_1558),
.B2(n_1542),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1539),
.A2(n_1517),
.B1(n_1531),
.B2(n_1507),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1556),
.A2(n_1517),
.B(n_1531),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1525),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1540),
.B(n_1533),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1537),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1559),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1552),
.B(n_1505),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1546),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1535),
.Y(n_1584)
);

NOR4xp25_ASAP7_75t_SL g1585 ( 
.A(n_1555),
.B(n_1522),
.C(n_1506),
.D(n_1492),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1538),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1538),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1537),
.Y(n_1588)
);

OAI211xp5_ASAP7_75t_L g1589 ( 
.A1(n_1543),
.A2(n_1515),
.B(n_1530),
.C(n_1502),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1539),
.A2(n_1517),
.B1(n_1531),
.B2(n_1524),
.C(n_1510),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1543),
.A2(n_1502),
.B(n_1523),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1558),
.A2(n_1531),
.B1(n_1510),
.B2(n_1504),
.C(n_1528),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1556),
.A2(n_1502),
.B1(n_1522),
.B2(n_1534),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1536),
.Y(n_1594)
);

AOI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1551),
.A2(n_1531),
.B1(n_1504),
.B2(n_1528),
.C(n_1499),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1555),
.A2(n_1502),
.B(n_1505),
.C(n_1534),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1545),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1545),
.B(n_1497),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1542),
.A2(n_1502),
.B1(n_1529),
.B2(n_1527),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1561),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1579),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1588),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1597),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1551),
.Y(n_1605)
);

OR2x4_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1546),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1581),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1576),
.A2(n_1560),
.B(n_1544),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1587),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1548),
.Y(n_1611)
);

NOR2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1563),
.B(n_1545),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

INVx4_ASAP7_75t_SL g1614 ( 
.A(n_1569),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1568),
.A2(n_1560),
.B(n_1547),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1567),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1572),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1566),
.A2(n_1560),
.B(n_1547),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1591),
.B(n_1596),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1592),
.A2(n_1560),
.B(n_1547),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1564),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1582),
.B(n_1527),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1584),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1584),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1571),
.B(n_1580),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.B(n_1527),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1580),
.B(n_1548),
.Y(n_1628)
);

INVx5_ASAP7_75t_L g1629 ( 
.A(n_1583),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1612),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1605),
.B(n_1593),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1585),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1600),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1621),
.B(n_1564),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1619),
.B(n_1614),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1617),
.A2(n_1589),
.B1(n_1563),
.B2(n_1575),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1602),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1605),
.B(n_1565),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1606),
.Y(n_1641)
);

NAND4xp75_ASAP7_75t_L g1642 ( 
.A(n_1619),
.B(n_1569),
.C(n_1595),
.D(n_1573),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1559),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1619),
.B(n_1564),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1598),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.B(n_1594),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1617),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1614),
.B(n_1574),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.B(n_1565),
.Y(n_1653)
);

OAI33xp33_ASAP7_75t_L g1654 ( 
.A1(n_1613),
.A2(n_1599),
.A3(n_1623),
.B1(n_1624),
.B2(n_1616),
.B3(n_1626),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1565),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1615),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1629),
.B(n_1604),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1625),
.B(n_1555),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1601),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1610),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1615),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1602),
.B(n_1570),
.C(n_1550),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1629),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1633),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1644),
.B(n_1622),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1636),
.A2(n_1606),
.B1(n_1627),
.B2(n_1618),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1644),
.B(n_1622),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1635),
.B(n_1430),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1655),
.B(n_1603),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1635),
.B(n_1629),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1637),
.B(n_1628),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1647),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1655),
.B(n_1603),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1638),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1628),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1635),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1636),
.B(n_1618),
.C(n_1620),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1607),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1631),
.B(n_1611),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1653),
.B(n_1608),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1664),
.B(n_1608),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1640),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1657),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1642),
.B(n_1611),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1650),
.A2(n_1618),
.B(n_1620),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1659),
.B(n_1618),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1665),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1656),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1655),
.B(n_1557),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1645),
.A2(n_1620),
.B1(n_1615),
.B2(n_1554),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1645),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1631),
.B(n_1613),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1660),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1660),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1659),
.B(n_1620),
.Y(n_1702)
);

NOR3xp33_ASAP7_75t_L g1703 ( 
.A(n_1692),
.B(n_1680),
.C(n_1689),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1645),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1694),
.Y(n_1705)
);

AO21x2_ASAP7_75t_L g1706 ( 
.A1(n_1690),
.A2(n_1648),
.B(n_1650),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1666),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1698),
.B(n_1672),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1698),
.B(n_1630),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1654),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1681),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1688),
.B(n_1630),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1681),
.Y(n_1718)
);

AOI31xp67_ASAP7_75t_L g1719 ( 
.A1(n_1695),
.A2(n_1648),
.A3(n_1658),
.B(n_1662),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1668),
.A2(n_1620),
.B1(n_1646),
.B2(n_1658),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1699),
.B(n_1646),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1685),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1685),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1667),
.B(n_1647),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1669),
.B(n_1647),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1671),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1675),
.Y(n_1727)
);

INVx3_ASAP7_75t_SL g1728 ( 
.A(n_1672),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1673),
.B(n_1661),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1711),
.A2(n_1706),
.B(n_1708),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1703),
.A2(n_1690),
.B1(n_1686),
.B2(n_1682),
.C(n_1693),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1719),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1727),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1722),
.B(n_1676),
.Y(n_1735)
);

OAI32xp33_ASAP7_75t_L g1736 ( 
.A1(n_1708),
.A2(n_1702),
.A3(n_1678),
.B1(n_1632),
.B2(n_1700),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1696),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1717),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1723),
.B(n_1688),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1728),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1706),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1712),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1726),
.B(n_1711),
.Y(n_1744)
);

INVxp33_ASAP7_75t_L g1745 ( 
.A(n_1710),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1728),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1704),
.A2(n_1697),
.B(n_1632),
.C(n_1641),
.Y(n_1747)
);

OAI31xp33_ASAP7_75t_L g1748 ( 
.A1(n_1720),
.A2(n_1658),
.A3(n_1656),
.B(n_1662),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1710),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1715),
.A2(n_1606),
.B1(n_1649),
.B2(n_1641),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1737),
.B(n_1745),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1730),
.B(n_1714),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1732),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1744),
.B(n_1750),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1749),
.B(n_1740),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1737),
.B(n_1718),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1742),
.B(n_1721),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1745),
.B(n_1712),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1749),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1746),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_SL g1763 ( 
.A1(n_1753),
.A2(n_1731),
.B(n_1736),
.C(n_1732),
.Y(n_1763)
);

NAND2x1_ASAP7_75t_L g1764 ( 
.A(n_1756),
.B(n_1716),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1754),
.A2(n_1748),
.B(n_1747),
.C(n_1736),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1759),
.A2(n_1741),
.B(n_1734),
.C(n_1762),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1762),
.B(n_1735),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1752),
.A2(n_1757),
.B(n_1755),
.Y(n_1768)
);

NOR2xp67_ASAP7_75t_L g1769 ( 
.A(n_1760),
.B(n_1705),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1733),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1758),
.A2(n_1741),
.B(n_1739),
.C(n_1738),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1761),
.A2(n_1716),
.B(n_1733),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1767),
.B(n_1716),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1763),
.A2(n_1743),
.B1(n_1695),
.B2(n_1707),
.C(n_1713),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1765),
.A2(n_1724),
.B(n_1725),
.C(n_1663),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1764),
.B(n_1634),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1768),
.B(n_1634),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1773),
.B(n_1769),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1778),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1776),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1774),
.B(n_1770),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1775),
.A2(n_1766),
.B1(n_1771),
.B2(n_1751),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1729),
.Y(n_1785)
);

CKINVDCx16_ASAP7_75t_R g1786 ( 
.A(n_1782),
.Y(n_1786)
);

AOI32xp33_ASAP7_75t_L g1787 ( 
.A1(n_1783),
.A2(n_1781),
.A3(n_1779),
.B1(n_1784),
.B2(n_1705),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1780),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1780),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1786),
.B(n_1705),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1788),
.B(n_1469),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1787),
.A2(n_1729),
.B(n_1663),
.C(n_1656),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1790),
.B(n_1789),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1791),
.C(n_1792),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1794),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1794),
.A2(n_1785),
.B1(n_1419),
.B2(n_1481),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1677),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1795),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1663),
.B(n_1662),
.Y(n_1799)
);

OAI22x1_ASAP7_75t_SL g1800 ( 
.A1(n_1797),
.A2(n_1694),
.B1(n_1444),
.B2(n_1701),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1799),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1801),
.B(n_1694),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1800),
.B(n_1687),
.Y(n_1803)
);

AOI22x1_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1444),
.B1(n_1691),
.B2(n_1683),
.Y(n_1804)
);

AOI31xp33_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1632),
.A3(n_1657),
.B(n_1652),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1665),
.B(n_1651),
.C(n_1643),
.Y(n_1806)
);


endmodule