module fake_jpeg_22852_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_SL g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx5_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_2),
.B(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVxp33_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_14),
.B(n_15),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_6),
.B1(n_10),
.B2(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_21),
.A2(n_16),
.B(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_17),
.C(n_5),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_0),
.C(n_3),
.Y(n_26)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_11),
.CI(n_25),
.CON(n_27),
.SN(n_27)
);


endmodule