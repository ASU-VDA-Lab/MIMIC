module fake_jpeg_24494_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_1),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_50),
.A2(n_51),
.B1(n_82),
.B2(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_18),
.B1(n_36),
.B2(n_20),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_56),
.B1(n_84),
.B2(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_20),
.B1(n_36),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_20),
.B1(n_36),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_63),
.B1(n_31),
.B2(n_28),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_61),
.B(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_35),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_69),
.Y(n_121)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_17),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_SL g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_86),
.Y(n_118)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_19),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_37),
.B1(n_23),
.B2(n_32),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_33),
.C(n_28),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_61),
.C(n_77),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_50),
.B1(n_51),
.B2(n_40),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_114),
.B1(n_119),
.B2(n_73),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_103),
.B1(n_111),
.B2(n_116),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_19),
.B1(n_32),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_37),
.B1(n_32),
.B2(n_27),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_37),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_110),
.C(n_54),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_32),
.B1(n_27),
.B2(n_25),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_16),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_27),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_25),
.B1(n_23),
.B2(n_10),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_25),
.B1(n_23),
.B2(n_3),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_25),
.B1(n_9),
.B2(n_11),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_88),
.B1(n_59),
.B2(n_84),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_129),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_66),
.B(n_60),
.C(n_70),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_143),
.B(n_147),
.Y(n_177)
);

OR2x4_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_109),
.B(n_97),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_59),
.B1(n_85),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_148),
.B1(n_151),
.B2(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_60),
.C(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_144),
.C(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_62),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_152),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_54),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_140),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_153),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_74),
.B1(n_78),
.B2(n_71),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_104),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_95),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_89),
.B(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_67),
.B1(n_65),
.B2(n_72),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_1),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_58),
.C(n_2),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_91),
.A2(n_112),
.A3(n_95),
.B1(n_107),
.B2(n_113),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_9),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_7),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_4),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_113),
.B(n_109),
.C(n_118),
.Y(n_147)
);

AO21x1_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_117),
.B(n_108),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_58),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_159),
.Y(n_190)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_175),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_115),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_173),
.C(n_155),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_115),
.B1(n_100),
.B2(n_98),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_169),
.B1(n_182),
.B2(n_151),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_172),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_140),
.B1(n_144),
.B2(n_132),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_98),
.B1(n_117),
.B2(n_6),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_4),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_5),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_180),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_127),
.A2(n_5),
.B(n_7),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_170),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_126),
.B(n_145),
.C(n_141),
.D(n_123),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g225 ( 
.A(n_187),
.B(n_188),
.C(n_202),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_129),
.B1(n_148),
.B2(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_194),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_195),
.B1(n_182),
.B2(n_174),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_132),
.B1(n_14),
.B2(n_15),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_156),
.B1(n_183),
.B2(n_184),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_158),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_163),
.C(n_162),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_172),
.B1(n_177),
.B2(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_222),
.B1(n_227),
.B2(n_185),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_188),
.B1(n_185),
.B2(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_219),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_177),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_200),
.B(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_192),
.B1(n_191),
.B2(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_181),
.C(n_176),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_226),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_156),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_171),
.C(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_238),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_234),
.B(n_242),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_187),
.B(n_188),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_244),
.B1(n_237),
.B2(n_242),
.Y(n_251)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_218),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_196),
.B1(n_202),
.B2(n_204),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_219),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_221),
.B1(n_210),
.B2(n_214),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_211),
.C(n_226),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_230),
.Y(n_264)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_209),
.B(n_222),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_258),
.B(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_224),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_257),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_223),
.B1(n_217),
.B2(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_154),
.B(n_175),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_263),
.B(n_252),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_239),
.B(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_230),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_232),
.B(n_160),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_261),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_253),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_275),
.B(n_264),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_247),
.B1(n_254),
.B2(n_248),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_270),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_257),
.B1(n_252),
.B2(n_246),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_267),
.B(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_256),
.B1(n_258),
.B2(n_251),
.C(n_215),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_260),
.C(n_266),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_232),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_279),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_281),
.B1(n_202),
.B2(n_157),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_287),
.B(n_285),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_160),
.Y(n_290)
);


endmodule