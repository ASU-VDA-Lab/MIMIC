module fake_jpeg_24202_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_16),
.B1(n_26),
.B2(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_40),
.B1(n_23),
.B2(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_44),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_34),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g46 ( 
.A(n_43),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_50),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_34),
.B(n_23),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_57),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_55),
.B1(n_67),
.B2(n_24),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_64),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_34),
.A3(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_61),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_60),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_21),
.B(n_13),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_13),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_66),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_1),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_3),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_17),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_22),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_4),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_30),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_76),
.Y(n_85)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_4),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_3),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_84),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_90),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_51),
.B(n_62),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_68),
.B(n_69),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_55),
.C(n_52),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_61),
.C(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_67),
.B1(n_48),
.B2(n_7),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_83),
.B1(n_72),
.B2(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_76),
.C(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_85),
.B1(n_89),
.B2(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_68),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_113),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_92),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_94),
.B1(n_98),
.B2(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_105),
.B1(n_104),
.B2(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_120),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_107),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_115),
.B(n_112),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_110),
.C(n_8),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_125),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_6),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_10),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_10),
.B(n_11),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_11),
.B(n_12),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_120),
.B1(n_122),
.B2(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_131),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_125),
.C(n_130),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_130),
.B(n_132),
.C(n_74),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_74),
.Y(n_136)
);


endmodule