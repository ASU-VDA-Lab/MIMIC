module real_aes_256_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_0), .B(n_113), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_1), .A2(n_122), .B(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_2), .A2(n_100), .B1(n_741), .B2(n_745), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_3), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_4), .B(n_113), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_5), .B(n_129), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_6), .B(n_129), .Y(n_499) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_8), .B(n_129), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_9), .Y(n_755) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_10), .B(n_131), .Y(n_480) );
AND2x2_ASAP7_75t_L g149 ( .A(n_11), .B(n_138), .Y(n_149) );
AND2x2_ASAP7_75t_L g158 ( .A(n_12), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
AOI221x1_ASAP7_75t_L g521 ( .A1(n_14), .A2(n_25), .B1(n_113), .B2(n_122), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_15), .B(n_129), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_16), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_17), .B(n_113), .Y(n_476) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_18), .A2(n_138), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_19), .B(n_133), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_20), .B(n_129), .Y(n_459) );
AO21x1_ASAP7_75t_L g494 ( .A1(n_21), .A2(n_113), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_22), .B(n_113), .Y(n_183) );
INVx1_ASAP7_75t_L g446 ( .A(n_23), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_24), .A2(n_87), .B1(n_113), .B2(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_26), .Y(n_769) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_27), .B(n_129), .Y(n_508) );
NAND2x1_ASAP7_75t_L g469 ( .A(n_28), .B(n_131), .Y(n_469) );
OR2x2_ASAP7_75t_L g136 ( .A(n_29), .B(n_84), .Y(n_136) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_29), .A2(n_84), .B(n_135), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_30), .B(n_131), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_31), .B(n_129), .Y(n_479) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_32), .A2(n_159), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_33), .B(n_131), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_34), .A2(n_122), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_35), .B(n_129), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_36), .A2(n_122), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g119 ( .A(n_37), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g123 ( .A(n_37), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g230 ( .A(n_37), .Y(n_230) );
OR2x6_ASAP7_75t_L g444 ( .A(n_38), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_39), .B(n_113), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_40), .B(n_113), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_41), .B(n_129), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_42), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_43), .B(n_131), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_44), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_45), .A2(n_122), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_46), .A2(n_122), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_47), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_48), .B(n_131), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_49), .B(n_113), .Y(n_165) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g126 ( .A(n_50), .Y(n_126) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_51), .A2(n_99), .B1(n_748), .B2(n_759), .C1(n_770), .C2(n_772), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g761 ( .A1(n_51), .A2(n_104), .B1(n_762), .B2(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_51), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_52), .B(n_129), .Y(n_156) );
AND2x2_ASAP7_75t_L g194 ( .A(n_53), .B(n_133), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_54), .B(n_131), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_55), .B(n_129), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_56), .B(n_131), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_57), .A2(n_122), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_58), .B(n_113), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_59), .B(n_113), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_60), .A2(n_122), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g189 ( .A(n_61), .B(n_134), .Y(n_189) );
AO21x1_ASAP7_75t_L g496 ( .A1(n_62), .A2(n_122), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_63), .B(n_113), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_64), .B(n_131), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_65), .B(n_113), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_66), .B(n_131), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_67), .A2(n_92), .B1(n_122), .B2(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_68), .B(n_129), .Y(n_186) );
AND2x2_ASAP7_75t_L g544 ( .A(n_69), .B(n_134), .Y(n_544) );
INVx1_ASAP7_75t_L g118 ( .A(n_70), .Y(n_118) );
INVx1_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
AND2x2_ASAP7_75t_L g472 ( .A(n_71), .B(n_159), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_72), .B(n_131), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_73), .A2(n_122), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_74), .A2(n_122), .B(n_127), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_75), .A2(n_122), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g180 ( .A(n_76), .B(n_134), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_77), .B(n_133), .Y(n_219) );
INVx1_ASAP7_75t_L g447 ( .A(n_78), .Y(n_447) );
INVx1_ASAP7_75t_L g100 ( .A(n_79), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_80), .B(n_113), .Y(n_461) );
AND2x2_ASAP7_75t_L g482 ( .A(n_81), .B(n_159), .Y(n_482) );
AND2x2_ASAP7_75t_L g137 ( .A(n_82), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g495 ( .A(n_83), .B(n_170), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_85), .B(n_131), .Y(n_460) );
AND2x2_ASAP7_75t_L g511 ( .A(n_86), .B(n_159), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_88), .B(n_129), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_89), .A2(n_122), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_90), .B(n_131), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_91), .A2(n_122), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_93), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_94), .B(n_129), .Y(n_487) );
BUFx2_ASAP7_75t_L g188 ( .A(n_95), .Y(n_188) );
BUFx2_ASAP7_75t_L g756 ( .A(n_96), .Y(n_756) );
BUFx2_ASAP7_75t_SL g776 ( .A(n_96), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_97), .A2(n_122), .B(n_478), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_101), .B(n_740), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_439), .B1(n_448), .B2(n_738), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_104), .A2(n_441), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx5_ASAP7_75t_L g762 ( .A(n_104), .Y(n_762) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_343), .Y(n_104) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_268), .C(n_304), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_242), .Y(n_106) );
AOI211xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_160), .B(n_190), .C(n_215), .Y(n_107) );
AND2x2_ASAP7_75t_L g333 ( .A(n_108), .B(n_192), .Y(n_333) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_140), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_109), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g366 ( .A(n_109), .B(n_248), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_109), .B(n_207), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_109), .B(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_109), .B(n_416), .Y(n_415) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_SL g202 ( .A(n_110), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g237 ( .A(n_110), .Y(n_237) );
AND2x2_ASAP7_75t_L g284 ( .A(n_110), .B(n_217), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_110), .B(n_140), .Y(n_303) );
BUFx2_ASAP7_75t_L g308 ( .A(n_110), .Y(n_308) );
AND2x2_ASAP7_75t_L g352 ( .A(n_110), .B(n_150), .Y(n_352) );
AND2x4_ASAP7_75t_L g424 ( .A(n_110), .B(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_110), .B(n_206), .Y(n_436) );
OR2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_137), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_121), .B(n_133), .Y(n_111) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_119), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND2x6_ASAP7_75t_L g131 ( .A(n_115), .B(n_124), .Y(n_131) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g129 ( .A(n_117), .B(n_126), .Y(n_129) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx5_ASAP7_75t_L g132 ( .A(n_119), .Y(n_132) );
AND2x2_ASAP7_75t_L g125 ( .A(n_120), .B(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_120), .Y(n_225) );
AND2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
BUFx3_ASAP7_75t_L g226 ( .A(n_123), .Y(n_226) );
INVx2_ASAP7_75t_L g232 ( .A(n_124), .Y(n_232) );
AND2x4_ASAP7_75t_L g228 ( .A(n_125), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_130), .B(n_132), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_131), .B(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_132), .A2(n_146), .B(n_147), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_132), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_132), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_132), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_132), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_132), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_132), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_132), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_132), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_132), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_132), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_132), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_132), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_132), .A2(n_541), .B(n_542), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_133), .Y(n_142) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_227), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_133), .A2(n_484), .B(n_485), .Y(n_483) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_133), .A2(n_521), .B(n_525), .Y(n_520) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_133), .A2(n_521), .B(n_525), .Y(n_532) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x4_ASAP7_75t_L g170 ( .A(n_135), .B(n_136), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_138), .A2(n_183), .B(n_184), .Y(n_182) );
BUFx4f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_140), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g355 ( .A(n_140), .Y(n_355) );
BUFx2_ASAP7_75t_L g404 ( .A(n_140), .Y(n_404) );
INVx1_ASAP7_75t_L g426 ( .A(n_140), .Y(n_426) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_150), .Y(n_140) );
INVx3_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_141), .Y(n_392) );
AOI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_149), .Y(n_141) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_142), .A2(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
INVx2_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_150), .B(n_203), .Y(n_207) );
INVx2_ASAP7_75t_L g292 ( .A(n_150), .Y(n_292) );
OR2x2_ASAP7_75t_L g299 ( .A(n_150), .B(n_248), .Y(n_299) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_158), .Y(n_150) );
INVx4_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
INVx3_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
AND2x2_ASAP7_75t_L g254 ( .A(n_160), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g288 ( .A(n_160), .B(n_251), .Y(n_288) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_171), .Y(n_160) );
AND2x2_ASAP7_75t_L g324 ( .A(n_161), .B(n_213), .Y(n_324) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g281 ( .A(n_162), .B(n_172), .Y(n_281) );
AND2x2_ASAP7_75t_L g400 ( .A(n_162), .B(n_181), .Y(n_400) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
INVx1_ASAP7_75t_L g240 ( .A(n_163), .Y(n_240) );
AND2x2_ASAP7_75t_L g296 ( .A(n_163), .B(n_172), .Y(n_296) );
AND2x2_ASAP7_75t_L g301 ( .A(n_163), .B(n_193), .Y(n_301) );
OR2x2_ASAP7_75t_L g364 ( .A(n_163), .B(n_181), .Y(n_364) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_163), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_170), .A2(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_SL g455 ( .A(n_170), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_170), .A2(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_170), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g192 ( .A(n_171), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
NOR2x1_ASAP7_75t_SL g171 ( .A(n_172), .B(n_181), .Y(n_171) );
AO21x1_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_172) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_214) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_173), .A2(n_505), .B(n_511), .Y(n_504) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_173), .A2(n_538), .B(n_544), .Y(n_537) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_173), .A2(n_538), .B(n_544), .Y(n_573) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_173), .A2(n_505), .B(n_511), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
AND2x2_ASAP7_75t_L g209 ( .A(n_181), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_SL g267 ( .A(n_181), .Y(n_267) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_181), .B(n_193), .Y(n_277) );
OR2x2_ASAP7_75t_L g282 ( .A(n_181), .B(n_210), .Y(n_282) );
BUFx2_ASAP7_75t_L g338 ( .A(n_181), .Y(n_338) );
AND2x2_ASAP7_75t_L g374 ( .A(n_181), .B(n_253), .Y(n_374) );
AND2x2_ASAP7_75t_L g385 ( .A(n_181), .B(n_213), .Y(n_385) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_189), .Y(n_181) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_201), .B1(n_207), .B2(n_208), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_192), .A2(n_382), .B1(n_432), .B2(n_437), .Y(n_431) );
INVx4_ASAP7_75t_L g210 ( .A(n_193), .Y(n_210) );
INVx2_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_193), .Y(n_322) );
OR2x2_ASAP7_75t_L g337 ( .A(n_193), .B(n_213), .Y(n_337) );
OR2x2_ASAP7_75t_SL g363 ( .A(n_193), .B(n_364), .Y(n_363) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx2_ASAP7_75t_SL g244 ( .A(n_202), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_202), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g312 ( .A(n_202), .B(n_260), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_202), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g234 ( .A(n_203), .Y(n_234) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_203), .Y(n_259) );
AND2x2_ASAP7_75t_L g315 ( .A(n_203), .B(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g425 ( .A(n_203), .Y(n_425) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_205), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_205), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g233 ( .A(n_206), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_207), .B(n_366), .Y(n_365) );
AOI321xp33_ASAP7_75t_L g387 ( .A1(n_208), .A2(n_289), .A3(n_357), .B1(n_388), .B2(n_389), .C(n_393), .Y(n_387) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_209), .Y(n_286) );
AND2x2_ASAP7_75t_L g311 ( .A(n_209), .B(n_240), .Y(n_311) );
AND2x2_ASAP7_75t_L g386 ( .A(n_209), .B(n_296), .Y(n_386) );
INVx1_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
BUFx2_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_210), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g310 ( .A(n_211), .Y(n_310) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
BUFx2_ASAP7_75t_L g317 ( .A(n_212), .Y(n_317) );
INVx2_ASAP7_75t_L g253 ( .A(n_213), .Y(n_253) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_213), .Y(n_276) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21xp33_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_235), .B(n_238), .Y(n_215) );
NOR2xp67_ASAP7_75t_L g369 ( .A(n_216), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
INVx3_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x4_ASAP7_75t_L g248 ( .A(n_219), .B(n_220), .Y(n_248) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NOR2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
INVx1_ASAP7_75t_SL g416 ( .A(n_234), .Y(n_416) );
INVxp33_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_237), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g342 ( .A(n_237), .B(n_299), .Y(n_342) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
AND2x2_ASAP7_75t_L g346 ( .A(n_239), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_239), .B(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_240), .B(n_277), .Y(n_332) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_240), .B(n_271), .C(n_428), .D(n_429), .Y(n_427) );
OR2x2_ASAP7_75t_L g395 ( .A(n_241), .B(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B1(n_254), .B2(n_256), .C(n_261), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g270 ( .A(n_245), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g307 ( .A(n_246), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_248), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
OR2x2_ASAP7_75t_L g294 ( .A(n_251), .B(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_253), .B(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
INVx2_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_258), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g263 ( .A(n_260), .Y(n_263) );
OAI321xp33_ASAP7_75t_L g375 ( .A1(n_260), .A2(n_368), .A3(n_376), .B1(n_381), .B2(n_383), .C(n_387), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g330 ( .A(n_263), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g430 ( .A(n_266), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_267), .B(n_310), .Y(n_309) );
NAND2xp33_ASAP7_75t_SL g410 ( .A(n_267), .B(n_281), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_283), .C(n_287), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
INVx3_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
OR2x2_ASAP7_75t_L g421 ( .A(n_277), .B(n_295), .Y(n_421) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_279), .A2(n_363), .B1(n_365), .B2(n_367), .Y(n_362) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_SL g361 ( .A(n_282), .Y(n_361) );
OR2x2_ASAP7_75t_L g438 ( .A(n_282), .B(n_295), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_289), .B(n_293), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_291), .B(n_308), .Y(n_407) );
AND2x2_ASAP7_75t_L g413 ( .A(n_291), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_300), .B2(n_302), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_338), .B(n_340), .C(n_342), .Y(n_339) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_298), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_298), .B(n_390), .Y(n_412) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_303), .A2(n_335), .B(n_338), .C(n_339), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g304 ( .A(n_305), .B(n_319), .C(n_334), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B1(n_311), .B2(n_312), .C1(n_313), .C2(n_316), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_308), .B(n_341), .Y(n_394) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g328 ( .A(n_315), .Y(n_328) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OR2x2_ASAP7_75t_L g433 ( .A(n_317), .B(n_350), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_318), .A2(n_409), .B1(n_411), .B2(n_413), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B1(n_329), .B2(n_332), .C(n_333), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp5_ASAP7_75t_SL g393 ( .A1(n_326), .A2(n_394), .B(n_395), .Y(n_393) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
AND2x2_ASAP7_75t_L g435 ( .A(n_327), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g419 ( .A(n_331), .Y(n_419) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g348 ( .A(n_337), .B(n_338), .Y(n_348) );
INVx1_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_375), .C(n_397), .Y(n_343) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B(n_351), .C(n_356), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_346), .A2(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_362), .C(n_369), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_364), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_366), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g396 ( .A(n_372), .Y(n_396) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_427), .Y(n_417) );
OAI21xp33_ASAP7_75t_SL g432 ( .A1(n_389), .A2(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_408), .C(n_417), .D(n_431), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_405), .B2(n_406), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
CKINVDCx6p67_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
AND2x6_ASAP7_75t_SL g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OR2x6_ASAP7_75t_SL g738 ( .A(n_443), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g747 ( .A(n_443), .B(n_444), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_443), .B(n_739), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_444), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_L g742 ( .A(n_448), .Y(n_742) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_636), .Y(n_448) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_548), .C(n_603), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_489), .B1(n_512), .B2(n_516), .C(n_526), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_473), .Y(n_451) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_452), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
AND2x2_ASAP7_75t_L g592 ( .A(n_452), .B(n_529), .Y(n_592) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g580 ( .A(n_454), .Y(n_580) );
INVx1_ASAP7_75t_L g590 ( .A(n_454), .Y(n_590) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_462), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_455), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_455), .A2(n_456), .B(n_462), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
OR2x2_ASAP7_75t_L g569 ( .A(n_464), .B(n_474), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_464), .B(n_515), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_464), .B(n_481), .Y(n_613) );
INVx2_ASAP7_75t_L g622 ( .A(n_464), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_464), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g727 ( .A(n_464), .B(n_546), .Y(n_727) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g555 ( .A(n_465), .B(n_481), .Y(n_555) );
AND2x2_ASAP7_75t_L g688 ( .A(n_465), .B(n_515), .Y(n_688) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_465), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
AND2x4_ASAP7_75t_L g642 ( .A(n_473), .B(n_643), .Y(n_642) );
AOI321xp33_ASAP7_75t_L g656 ( .A1(n_473), .A2(n_585), .A3(n_586), .B1(n_618), .B2(n_657), .C(n_660), .Y(n_656) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_481), .Y(n_473) );
BUFx3_ASAP7_75t_L g513 ( .A(n_474), .Y(n_513) );
INVx2_ASAP7_75t_L g546 ( .A(n_474), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_474), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g579 ( .A(n_474), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g612 ( .A(n_474), .Y(n_612) );
INVx5_ASAP7_75t_L g515 ( .A(n_481), .Y(n_515) );
NOR2x1_ASAP7_75t_SL g564 ( .A(n_481), .B(n_554), .Y(n_564) );
BUFx2_ASAP7_75t_L g659 ( .A(n_481), .Y(n_659) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVxp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
NOR2xp33_ASAP7_75t_SL g557 ( .A(n_491), .B(n_558), .Y(n_557) );
NOR4xp25_ASAP7_75t_L g660 ( .A(n_491), .B(n_654), .C(n_658), .D(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g698 ( .A(n_491), .Y(n_698) );
AND2x2_ASAP7_75t_L g732 ( .A(n_491), .B(n_672), .Y(n_732) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g533 ( .A(n_492), .Y(n_533) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
OAI21x1_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g501 ( .A(n_495), .Y(n_501) );
AOI33xp33_ASAP7_75t_L g728 ( .A1(n_502), .A2(n_530), .A3(n_561), .B1(n_577), .B2(n_683), .B3(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g518 ( .A(n_503), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g528 ( .A(n_503), .B(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g535 ( .A(n_504), .Y(n_535) );
INVxp67_ASAP7_75t_L g616 ( .A(n_504), .Y(n_616) );
AND2x2_ASAP7_75t_L g672 ( .A(n_504), .B(n_537), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_512), .A2(n_694), .B(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_L g681 ( .A(n_513), .B(n_555), .Y(n_681) );
AND3x2_ASAP7_75t_L g683 ( .A(n_513), .B(n_567), .C(n_622), .Y(n_683) );
INVx3_ASAP7_75t_SL g635 ( .A(n_514), .Y(n_635) );
INVx4_ASAP7_75t_L g529 ( .A(n_515), .Y(n_529) );
AND2x2_ASAP7_75t_L g567 ( .A(n_515), .B(n_554), .Y(n_567) );
INVxp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g561 ( .A(n_519), .Y(n_561) );
AND2x4_ASAP7_75t_L g586 ( .A(n_519), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g649 ( .A(n_519), .B(n_537), .Y(n_649) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g619 ( .A(n_520), .Y(n_619) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_R g526 ( .A1(n_527), .A2(n_530), .B(n_534), .C(n_545), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g578 ( .A(n_529), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_529), .B(n_546), .Y(n_707) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g689 ( .A(n_531), .B(n_679), .Y(n_689) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g536 ( .A(n_532), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g558 ( .A(n_532), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g574 ( .A(n_532), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g607 ( .A(n_532), .B(n_587), .Y(n_607) );
AND2x4_ASAP7_75t_L g572 ( .A(n_533), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g596 ( .A(n_533), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g634 ( .A(n_533), .B(n_559), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g562 ( .A(n_535), .B(n_559), .Y(n_562) );
AND2x2_ASAP7_75t_L g577 ( .A(n_535), .B(n_537), .Y(n_577) );
BUFx2_ASAP7_75t_L g633 ( .A(n_535), .Y(n_633) );
AND2x2_ASAP7_75t_L g647 ( .A(n_535), .B(n_558), .Y(n_647) );
INVx2_ASAP7_75t_L g559 ( .A(n_537), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_539), .B(n_543), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_545), .A2(n_596), .B1(n_598), .B2(n_602), .Y(n_595) );
INVx2_ASAP7_75t_SL g626 ( .A(n_545), .Y(n_626) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_L g601 ( .A(n_546), .B(n_554), .Y(n_601) );
INVx1_ASAP7_75t_L g708 ( .A(n_547), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_581), .C(n_595), .Y(n_548) );
OAI221xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_556), .B1(n_560), .B2(n_563), .C(n_565), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g609 ( .A(n_553), .Y(n_609) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_553), .Y(n_737) );
INVx1_ASAP7_75t_L g700 ( .A(n_555), .Y(n_700) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_555), .B(n_579), .Y(n_710) );
INVxp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_559), .B(n_587), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OR2x2_ASAP7_75t_L g593 ( .A(n_561), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g671 ( .A(n_561), .Y(n_671) );
AND2x2_ASAP7_75t_L g606 ( .A(n_562), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g652 ( .A(n_564), .B(n_612), .Y(n_652) );
AND2x2_ASAP7_75t_L g729 ( .A(n_564), .B(n_727), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_570), .B1(n_577), .B2(n_578), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g588 ( .A(n_569), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx2_ASAP7_75t_L g594 ( .A(n_572), .Y(n_594) );
AND2x4_ASAP7_75t_L g618 ( .A(n_572), .B(n_619), .Y(n_618) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_572), .A2(n_649), .B(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g675 ( .A(n_572), .B(n_633), .Y(n_675) );
INVx2_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_573), .Y(n_630) );
INVx1_ASAP7_75t_SL g654 ( .A(n_574), .Y(n_654) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g585 ( .A(n_576), .Y(n_585) );
AND2x4_ASAP7_75t_SL g679 ( .A(n_576), .B(n_597), .Y(n_679) );
AND2x2_ASAP7_75t_L g676 ( .A(n_579), .B(n_622), .Y(n_676) );
AND2x2_ASAP7_75t_L g702 ( .A(n_579), .B(n_688), .Y(n_702) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
INVx1_ASAP7_75t_L g644 ( .A(n_580), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_588), .B1(n_591), .B2(n_593), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_586), .B(n_597), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_586), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g725 ( .A(n_586), .Y(n_725) );
INVx2_ASAP7_75t_SL g650 ( .A(n_588), .Y(n_650) );
AND2x2_ASAP7_75t_L g662 ( .A(n_590), .B(n_622), .Y(n_662) );
INVx2_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
INVxp33_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g627 ( .A(n_593), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_596), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g718 ( .A(n_596), .Y(n_718) );
INVx1_ASAP7_75t_L g646 ( .A(n_598), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_599), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g657 ( .A(n_601), .B(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_601), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_625), .C(n_628), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B1(n_610), .B2(n_614), .C(n_617), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g723 ( .A(n_608), .Y(n_723) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g692 ( .A(n_609), .B(n_658), .Y(n_692) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g623 ( .A(n_612), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g694 ( .A(n_614), .Y(n_694) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g691 ( .A(n_615), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_616), .Y(n_697) );
OR2x2_ASAP7_75t_L g720 ( .A(n_616), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_SL g629 ( .A(n_619), .Y(n_629) );
AND2x2_ASAP7_75t_L g699 ( .A(n_619), .B(n_679), .Y(n_699) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_619), .B(n_632), .Y(n_731) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g736 ( .A(n_622), .Y(n_736) );
INVx1_ASAP7_75t_L g686 ( .A(n_624), .Y(n_686) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_631), .C(n_635), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_629), .B(n_679), .Y(n_703) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_632), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g640 ( .A(n_634), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g721 ( .A(n_634), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g636 ( .A(n_637), .B(n_693), .C(n_709), .D(n_730), .Y(n_636) );
NOR3x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_655), .C(n_677), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_639), .B(n_645), .C(n_648), .D(n_651), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_642), .Y(n_639) );
AND2x2_ASAP7_75t_L g690 ( .A(n_641), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g715 ( .A(n_642), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_SL g704 ( .A(n_647), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .Y(n_655) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_659), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_669), .B(n_673), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI322xp33_ASAP7_75t_L g695 ( .A1(n_667), .A2(n_696), .A3(n_700), .B1(n_701), .B2(n_703), .C1(n_704), .C2(n_705), .Y(n_695) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_668), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_671), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_672), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_682), .C(n_684), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_684) );
NOR2xp33_ASAP7_75t_SL g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_699), .Y(n_696) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_702), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g712 ( .A(n_707), .B(n_713), .Y(n_712) );
O2A1O1Ixp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_716), .C(n_719), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_712), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI221xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_722), .B1(n_724), .B2(n_726), .C(n_728), .Y(n_719) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
CKINVDCx11_ASAP7_75t_R g744 ( .A(n_738), .Y(n_744) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_757), .Y(n_750) );
INVxp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_756), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_SL g771 ( .A(n_754), .B(n_756), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_754), .A2(n_774), .B(n_777), .Y(n_773) );
INVx1_ASAP7_75t_SL g765 ( .A(n_757), .Y(n_765) );
BUFx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
BUFx3_ASAP7_75t_L g768 ( .A(n_758), .Y(n_768) );
BUFx2_ASAP7_75t_L g778 ( .A(n_758), .Y(n_778) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .B(n_766), .Y(n_760) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_SL g766 ( .A(n_767), .B(n_769), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
CKINVDCx8_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
endmodule