module fake_jpeg_19572_n_189 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_21),
.B1(n_12),
.B2(n_23),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_13),
.B(n_31),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_49),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_27),
.C(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_49),
.Y(n_62)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_40),
.B1(n_32),
.B2(n_43),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_41),
.B(n_40),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_76),
.B1(n_70),
.B2(n_37),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_13),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_19),
.B(n_17),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_27),
.B1(n_24),
.B2(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_76),
.B1(n_66),
.B2(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_64),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_81),
.C(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_66),
.B1(n_73),
.B2(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_75),
.B(n_67),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_104),
.B(n_77),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_75),
.B(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_64),
.B1(n_47),
.B2(n_62),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_71),
.B1(n_37),
.B2(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_111),
.B(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_112),
.C(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_78),
.B1(n_84),
.B2(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_78),
.C(n_58),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_121),
.B1(n_39),
.B2(n_30),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_85),
.B(n_83),
.C(n_27),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_56),
.B(n_68),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_50),
.B(n_20),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_24),
.B1(n_59),
.B2(n_103),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_129),
.C(n_132),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_106),
.B1(n_93),
.B2(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_136),
.B1(n_137),
.B2(n_116),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_120),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_96),
.CI(n_50),
.CON(n_128),
.SN(n_128)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_25),
.C(n_33),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_59),
.C(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_20),
.C(n_14),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_114),
.B1(n_117),
.B2(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_145),
.B1(n_126),
.B2(n_133),
.Y(n_151)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_136),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_122),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_137),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_114),
.B(n_122),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_148),
.B1(n_113),
.B2(n_121),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_107),
.B1(n_121),
.B2(n_113),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_129),
.C(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_154),
.C(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_149),
.B1(n_148),
.B2(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_159),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_133),
.C(n_111),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_163),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_146),
.C(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_18),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_14),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_SL g174 ( 
.A(n_166),
.B(n_168),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_R g168 ( 
.A(n_159),
.B(n_7),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_152),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_175),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_167),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_174),
.A3(n_167),
.B1(n_18),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_180),
.B(n_10),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.C(n_10),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_6),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_182),
.B(n_184),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_1),
.B1(n_186),
.B2(n_164),
.Y(n_189)
);


endmodule