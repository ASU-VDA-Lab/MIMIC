module fake_jpeg_1567_n_325 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_46),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_49),
.Y(n_90)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_25),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_61),
.Y(n_117)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_53),
.Y(n_140)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_55),
.Y(n_135)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx2_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_26),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_74),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_22),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_2),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_30),
.B(n_2),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_33),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_16),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_45),
.B1(n_36),
.B2(n_29),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_91),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_36),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_95),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_23),
.C(n_38),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_65),
.C(n_53),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_36),
.B1(n_29),
.B2(n_43),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_29),
.B1(n_43),
.B2(n_27),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_117),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_42),
.B1(n_34),
.B2(n_35),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_126),
.B1(n_128),
.B2(n_71),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_27),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_114),
.B(n_96),
.Y(n_185)
);

CKINVDCx12_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_125),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_37),
.B1(n_32),
.B2(n_35),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_60),
.A2(n_42),
.B1(n_34),
.B2(n_32),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_48),
.B1(n_52),
.B2(n_55),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_4),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_137),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_62),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_54),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_56),
.B(n_6),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_91),
.B1(n_121),
.B2(n_138),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_86),
.B1(n_78),
.B2(n_67),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_147),
.A2(n_165),
.B1(n_116),
.B2(n_113),
.Y(n_193)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_46),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_7),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_168),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_95),
.B(n_9),
.CI(n_11),
.CON(n_155),
.SN(n_155)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_155),
.B(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_97),
.A2(n_9),
.B(n_12),
.C(n_14),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_170),
.B(n_175),
.Y(n_186)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_166),
.Y(n_198)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_167),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_14),
.B1(n_15),
.B2(n_133),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_15),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_174),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_92),
.A2(n_15),
.B(n_137),
.C(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_115),
.B(n_111),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_94),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_108),
.A2(n_119),
.B(n_128),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_140),
.C(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_104),
.B(n_112),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_94),
.B(n_110),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_105),
.B(n_138),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_151),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_96),
.B(n_141),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_102),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_116),
.B1(n_141),
.B2(n_102),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_149),
.B1(n_161),
.B2(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_190),
.B(n_204),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_206),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_164),
.B1(n_167),
.B2(n_163),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_124),
.B1(n_134),
.B2(n_113),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_195),
.A2(n_217),
.B1(n_213),
.B2(n_209),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_124),
.B(n_134),
.C(n_151),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_180),
.B(n_206),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_154),
.B1(n_153),
.B2(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_142),
.B(n_168),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_142),
.A2(n_151),
.B1(n_155),
.B2(n_181),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_151),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_225),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_144),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_234),
.B(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_217),
.B1(n_195),
.B2(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_159),
.C(n_166),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_235),
.C(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_198),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_243),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_231),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_210),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_194),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_186),
.A2(n_219),
.B(n_205),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_214),
.B(n_200),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_202),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_189),
.C(n_197),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_203),
.C(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_214),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_213),
.B1(n_212),
.B2(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_247),
.B1(n_259),
.B2(n_231),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_256),
.C(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_217),
.B(n_194),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_242),
.C(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_192),
.B(n_198),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_211),
.B(n_201),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_264),
.B(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_246),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_239),
.C(n_235),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_228),
.C(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_229),
.C(n_231),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_216),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_244),
.C(n_224),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_222),
.C(n_211),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_253),
.C(n_223),
.Y(n_289)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_289),
.C(n_267),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_252),
.B(n_278),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_263),
.B1(n_274),
.B2(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_258),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_302),
.B1(n_294),
.B2(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_282),
.C(n_283),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_276),
.B(n_245),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_260),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_282),
.C(n_286),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_286),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

AOI31xp67_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_289),
.A3(n_287),
.B(n_288),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_304),
.A3(n_281),
.B1(n_295),
.B2(n_302),
.C1(n_297),
.C2(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_310),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_305),
.B(n_260),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.C(n_192),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_262),
.C(n_240),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_262),
.C(n_201),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_319),
.B(n_227),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_192),
.C(n_226),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_323),
.B(n_192),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_226),
.Y(n_325)
);


endmodule