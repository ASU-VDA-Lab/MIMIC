module fake_jpeg_25126_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_45),
.Y(n_61)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_52),
.B(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_75),
.Y(n_114)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_44),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_83),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_44),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_68),
.C(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_38),
.B1(n_46),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_94),
.B1(n_56),
.B2(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_24),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_61),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_38),
.B1(n_46),
.B2(n_42),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_33),
.Y(n_107)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_62),
.B1(n_58),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_84),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_91),
.B1(n_97),
.B2(n_74),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_126),
.B(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_122),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_58),
.B1(n_20),
.B2(n_23),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_120),
.B1(n_124),
.B2(n_78),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_77),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_70),
.B(n_77),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_10),
.B(n_13),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_25),
.B1(n_29),
.B2(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_20),
.B1(n_25),
.B2(n_29),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_73),
.B1(n_93),
.B2(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_75),
.B1(n_80),
.B2(n_73),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_132),
.B1(n_135),
.B2(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_139),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_143),
.Y(n_159)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

BUFx24_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_82),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_134),
.B(n_149),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_71),
.B1(n_72),
.B2(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_137),
.B(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_79),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_99),
.B1(n_107),
.B2(n_101),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_109),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_146),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_94),
.B1(n_87),
.B2(n_88),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_88),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_153),
.Y(n_182)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_115),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_121),
.B(n_101),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_45),
.B1(n_17),
.B2(n_27),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_100),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_105),
.B1(n_119),
.B2(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_160),
.B1(n_168),
.B2(n_134),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_105),
.B1(n_120),
.B2(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_174),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_180),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_102),
.B(n_121),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_148),
.B(n_146),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_124),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_139),
.C(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_152),
.B1(n_156),
.B2(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_129),
.A2(n_132),
.B1(n_149),
.B2(n_128),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_114),
.B1(n_100),
.B2(n_113),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_114),
.B1(n_113),
.B2(n_115),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_136),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_141),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_177),
.B(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_169),
.B1(n_189),
.B2(n_179),
.Y(n_228)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_218),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_134),
.B1(n_151),
.B2(n_155),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_179),
.B(n_174),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_184),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_157),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_150),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_207),
.B(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_143),
.C(n_131),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_181),
.C(n_185),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_171),
.B(n_9),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_239),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_225),
.B(n_226),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_187),
.B(n_172),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_244),
.C(n_194),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_211),
.B1(n_217),
.B2(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_168),
.B1(n_160),
.B2(n_187),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_236),
.B1(n_205),
.B2(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_12),
.C(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_10),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_169),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_27),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_165),
.C(n_161),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_201),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_175),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_200),
.A2(n_161),
.B1(n_158),
.B2(n_30),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_204),
.B1(n_215),
.B2(n_158),
.Y(n_259)
);

FAx1_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_225),
.CI(n_203),
.CON(n_248),
.SN(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_267),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_255),
.B1(n_222),
.B2(n_234),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_253),
.B1(n_259),
.B2(n_264),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_196),
.B1(n_195),
.B2(n_202),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_211),
.B1(n_219),
.B2(n_191),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_197),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_193),
.C(n_199),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_258),
.C(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_193),
.C(n_214),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_214),
.B(n_175),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_214),
.B1(n_115),
.B2(n_175),
.Y(n_264)
);

AOI31xp33_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_17),
.A3(n_19),
.B(n_34),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_252),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_255),
.C(n_249),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_284),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_230),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_276),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_230),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_283),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_226),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_223),
.C(n_232),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_285),
.C(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_223),
.C(n_242),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_12),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_260),
.C(n_265),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_292),
.C(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_279),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_254),
.C(n_237),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_237),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_261),
.B1(n_220),
.B2(n_242),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_229),
.B1(n_248),
.B2(n_274),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_248),
.B1(n_229),
.B2(n_224),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_282),
.C(n_285),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_287),
.B(n_293),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_311),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_246),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_312),
.C(n_313),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_296),
.B1(n_300),
.B2(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_34),
.C(n_9),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_0),
.C(n_1),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_2),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_0),
.C(n_2),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_323),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_0),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_304),
.B(n_2),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_302),
.B1(n_309),
.B2(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_330),
.A3(n_318),
.B1(n_321),
.B2(n_6),
.C1(n_7),
.C2(n_4),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_3),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_3),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_317),
.B(n_333),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_332),
.C(n_324),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_326),
.B(n_316),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_316),
.C(n_329),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_6),
.CI(n_7),
.CON(n_340),
.SN(n_340)
);


endmodule