module fake_jpeg_16667_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_42),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_23),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_31),
.B1(n_34),
.B2(n_22),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_13),
.C(n_17),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_13),
.C(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_27),
.B1(n_46),
.B2(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_63),
.B1(n_21),
.B2(n_5),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_59),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_6),
.C(n_7),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_38),
.B(n_46),
.C(n_40),
.D(n_34),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_61),
.B1(n_9),
.B2(n_10),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_4),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_56),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_54),
.C(n_58),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_52),
.B(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_86),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_68),
.C(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.C(n_81),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

AO221x1_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_82),
.B1(n_60),
.B2(n_61),
.C(n_75),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_77),
.B1(n_66),
.B2(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_88),
.C(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_60),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_62),
.B(n_50),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_87),
.B(n_90),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_97),
.C(n_94),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_104),
.C(n_105),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_89),
.C(n_11),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_108),
.Y(n_110)
);


endmodule