module fake_jpeg_30129_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_12),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_SL g38 ( 
.A1(n_21),
.A2(n_1),
.B(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_42),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_19),
.C(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_29),
.B(n_28),
.Y(n_50)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_SL g59 ( 
.A(n_30),
.B(n_20),
.C(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_32),
.B1(n_26),
.B2(n_41),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_64),
.B1(n_74),
.B2(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_25),
.B1(n_23),
.B2(n_16),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_20),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_75),
.B(n_12),
.C(n_10),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_16),
.B(n_14),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_57),
.B(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_25),
.B1(n_14),
.B2(n_20),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_8),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_3),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_8),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_53),
.C(n_52),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.C(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_44),
.B1(n_55),
.B2(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_51),
.B1(n_78),
.B2(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_44),
.C(n_51),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_92),
.B(n_75),
.C(n_71),
.D(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_76),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_91),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_87),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_65),
.B1(n_70),
.B2(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_100),
.B(n_102),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_57),
.B1(n_6),
.B2(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_6),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_110),
.C(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_112),
.B1(n_94),
.B2(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_104),
.C(n_98),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.C(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_90),
.C(n_99),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_92),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_88),
.B1(n_113),
.B2(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_123),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_111),
.B(n_102),
.C(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_83),
.A3(n_93),
.B1(n_58),
.B2(n_68),
.C1(n_9),
.C2(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_115),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_83),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_121),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_129),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_68),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_45),
.Y(n_134)
);


endmodule