module fake_netlist_5_650_n_2592 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_520, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2592);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_520;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2592;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2282;
wire n_2002;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_336),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_321),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_136),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_58),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_462),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_358),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_252),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_539),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_536),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_390),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_129),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_303),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_288),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_377),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_115),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_475),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_38),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_99),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_6),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_86),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_381),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_232),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_542),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_371),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_171),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_537),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_398),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_99),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_195),
.Y(n_587)
);

CKINVDCx14_ASAP7_75t_R g588 ( 
.A(n_319),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_204),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_300),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_77),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_62),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_95),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_535),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_538),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_355),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_484),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_547),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_369),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_66),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_490),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_502),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_21),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_211),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_12),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_61),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_305),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_256),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_80),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_477),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_119),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_403),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_479),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_268),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_194),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_332),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_21),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_339),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_272),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_3),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_91),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_214),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_439),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_354),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_208),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_333),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_361),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_273),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_54),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_349),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_224),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_125),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_168),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_143),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_394),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_392),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_202),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_67),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_206),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_316),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_452),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_550),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_140),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_446),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_156),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_210),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_528),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_163),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_329),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_94),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_56),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_100),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_518),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_69),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_42),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_172),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_86),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_116),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_226),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_413),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_109),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_543),
.Y(n_662)
);

BUFx8_ASAP7_75t_SL g663 ( 
.A(n_117),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_476),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_124),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_494),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_123),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_529),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_341),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_359),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_146),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_110),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_416),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_58),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_267),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_37),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_308),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_127),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_549),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_332),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_541),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_180),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_221),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_306),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_530),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_533),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_2),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_42),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_260),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_96),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_367),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_531),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_492),
.Y(n_693)
);

INVx4_ASAP7_75t_R g694 ( 
.A(n_493),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_411),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_117),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_263),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_510),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_169),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_521),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_208),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_79),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_362),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_319),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_548),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_187),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_365),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_105),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_449),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_545),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_72),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_44),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_443),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_540),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_374),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_40),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_128),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_505),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_139),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_156),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_165),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_186),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_546),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_282),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_32),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_182),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_364),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_307),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_509),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_342),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_544),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_210),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_324),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_143),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_527),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_189),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_123),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_301),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_522),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_78),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_59),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_532),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_78),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_400),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_221),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_395),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_506),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_426),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_108),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_290),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_324),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_5),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_44),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_38),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_184),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_60),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_50),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_440),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_534),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_328),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_279),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_236),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_108),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_296),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_337),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_434),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_195),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_293),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_357),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_415),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_65),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_467),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_193),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_495),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_62),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_18),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_181),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_454),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_153),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_328),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_331),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_36),
.Y(n_782)
);

BUFx8_ASAP7_75t_SL g783 ( 
.A(n_274),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_635),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_663),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_663),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_632),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_765),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_765),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_765),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_783),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_783),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_571),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_571),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_588),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_628),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_604),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_604),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_606),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_626),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_553),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

INVxp33_ASAP7_75t_SL g803 ( 
.A(n_587),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_708),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_736),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_708),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_730),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_730),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_604),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_604),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_619),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_572),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_678),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_572),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_619),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_619),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_619),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_654),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_654),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_654),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_740),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_554),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_555),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_654),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_558),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_734),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_556),
.B(n_0),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_567),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_734),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_734),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_734),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_563),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_575),
.Y(n_833)
);

INVx4_ASAP7_75t_R g834 ( 
.A(n_557),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_586),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_575),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_589),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_767),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_561),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_590),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_579),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_593),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_608),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_569),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_582),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_574),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_611),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_614),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_579),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_615),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_617),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_556),
.B(n_0),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_561),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_591),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_592),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_600),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_605),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_633),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_645),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_650),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_651),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_564),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_657),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_621),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_658),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_581),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_661),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_665),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_675),
.Y(n_869)
);

INVxp33_ASAP7_75t_L g870 ( 
.A(n_677),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_680),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_696),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_603),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_699),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_609),
.Y(n_875)
);

CKINVDCx16_ASAP7_75t_R g876 ( 
.A(n_566),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_557),
.B(n_1),
.Y(n_877)
);

CKINVDCx14_ASAP7_75t_R g878 ( 
.A(n_576),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_706),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_558),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_713),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_576),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_621),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_656),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_712),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_716),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_811),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_809),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_812),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_795),
.Y(n_891)
);

CKINVDCx14_ASAP7_75t_R g892 ( 
.A(n_878),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_795),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_816),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_876),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_817),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_833),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_786),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_786),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_799),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_818),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_784),
.B(n_562),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_801),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_801),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_824),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_799),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_822),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_833),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_814),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_836),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_826),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_829),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_825),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_830),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_831),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_797),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_881),
.B(n_822),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_797),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_836),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_800),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_841),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_798),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_823),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_798),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_825),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_841),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_823),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_828),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_849),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_828),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_844),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_846),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_815),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_844),
.B(n_580),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_815),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_845),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_819),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_849),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_873),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_825),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_819),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_800),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_785),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_845),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_820),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_820),
.Y(n_947)
);

INVxp67_ASAP7_75t_SL g948 ( 
.A(n_825),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_R g949 ( 
.A(n_854),
.B(n_573),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_785),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_811),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_854),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_917),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_907),
.B(n_889),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_917),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_910),
.B(n_832),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_907),
.B(n_788),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_919),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_892),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_902),
.B(n_789),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_897),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_923),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_888),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_887),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_890),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_894),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_896),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_SL g968 ( 
.A(n_891),
.B(n_566),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_887),
.A2(n_862),
.B(n_790),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_914),
.B(n_855),
.Y(n_970)
);

OAI22x1_ASAP7_75t_SL g971 ( 
.A1(n_909),
.A2(n_873),
.B1(n_607),
.B2(n_631),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_901),
.Y(n_972)
);

AOI22x1_ASAP7_75t_SL g973 ( 
.A1(n_911),
.A2(n_603),
.B1(n_631),
.B2(n_607),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_905),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_925),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_912),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_920),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_935),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_933),
.A2(n_803),
.B1(n_838),
.B2(n_787),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_913),
.B(n_839),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_915),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_916),
.B(n_839),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_934),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_936),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_938),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_942),
.B(n_853),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_946),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_947),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_949),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_926),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_941),
.B(n_855),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_948),
.B(n_853),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_918),
.B(n_856),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_906),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_921),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_943),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_903),
.B(n_856),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_903),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_900),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_SL g1000 ( 
.A1(n_922),
.A2(n_669),
.B1(n_719),
.B2(n_652),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_900),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_904),
.B(n_846),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_904),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_891),
.A2(n_803),
.B1(n_875),
.B2(n_857),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_895),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_952),
.B(n_864),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_908),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_893),
.A2(n_875),
.B1(n_857),
.B2(n_773),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_908),
.B(n_864),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_924),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_924),
.B(n_881),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_928),
.B(n_883),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_928),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_895),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_929),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_893),
.A2(n_568),
.B1(n_852),
.B2(n_827),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_929),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_931),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_931),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_932),
.B(n_883),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_932),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_937),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_937),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_945),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_945),
.B(n_877),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_952),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_898),
.B(n_882),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_944),
.B(n_813),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_899),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_899),
.B(n_877),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_950),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_927),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_SL g1034 ( 
.A1(n_940),
.A2(n_669),
.B1(n_719),
.B2(n_652),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_930),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_939),
.B(n_825),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_917),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_902),
.B(n_581),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_951),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_902),
.A2(n_610),
.B1(n_636),
.B2(n_599),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_953),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1006),
.B(n_813),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1025),
.B(n_558),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1006),
.B(n_884),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_982),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_993),
.B(n_599),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1020),
.B(n_884),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_986),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_982),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_986),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_957),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_957),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_963),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_986),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_965),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_R g1056 ( 
.A(n_989),
.B(n_574),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_966),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1020),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_967),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_953),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_998),
.B(n_791),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1025),
.B(n_558),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_972),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_954),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_992),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_SL g1066 ( 
.A1(n_1034),
.A2(n_756),
.B1(n_764),
.B2(n_726),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_974),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_976),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_955),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_954),
.B(n_835),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_955),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_960),
.B(n_884),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_981),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1040),
.A2(n_1025),
.B1(n_956),
.B2(n_1031),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_980),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1037),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_980),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1009),
.B(n_598),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_964),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_964),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_964),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_960),
.B(n_851),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1009),
.B(n_598),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1037),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_954),
.A2(n_636),
.B1(n_718),
.B2(n_610),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1039),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_958),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_961),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_958),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_962),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_962),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_1028),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_1038),
.B(n_718),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_975),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_1028),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_975),
.Y(n_1096)
);

AND3x1_ASAP7_75t_L g1097 ( 
.A(n_968),
.B(n_792),
.C(n_805),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1009),
.B(n_821),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1012),
.B(n_622),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_984),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_987),
.Y(n_1101)
);

INVx6_ASAP7_75t_L g1102 ( 
.A(n_983),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1012),
.A2(n_664),
.B1(n_769),
.B2(n_641),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_990),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_990),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1000),
.A2(n_756),
.B1(n_764),
.B2(n_726),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1012),
.Y(n_1107)
);

NOR2x1_ASAP7_75t_L g1108 ( 
.A(n_1036),
.B(n_584),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_969),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_983),
.Y(n_1110)
);

BUFx3_ASAP7_75t_SL g1111 ( 
.A(n_1038),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_969),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_959),
.B(n_771),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_969),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1031),
.B(n_698),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_983),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_985),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_985),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1002),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1031),
.B(n_585),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_985),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_970),
.B(n_644),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_985),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_988),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_961),
.A2(n_771),
.B1(n_780),
.B2(n_577),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_988),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_996),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_989),
.B(n_870),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_988),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_SL g1130 ( 
.A1(n_977),
.A2(n_1033),
.B1(n_1035),
.B2(n_1032),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_988),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_991),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1011),
.B(n_698),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_978),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1011),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_996),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_994),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1013),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_995),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1013),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1017),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1017),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1016),
.A2(n_731),
.B1(n_739),
.B2(n_707),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_999),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_SL g1145 ( 
.A(n_1021),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1001),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1003),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_SL g1148 ( 
.A1(n_977),
.A2(n_577),
.B1(n_781),
.B2(n_780),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1007),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1024),
.B(n_997),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1010),
.Y(n_1151)
);

INVxp33_ASAP7_75t_L g1152 ( 
.A(n_997),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1015),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1018),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1019),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1003),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1022),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1026),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1024),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1024),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1003),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1027),
.B(n_707),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1003),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1023),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1008),
.A2(n_560),
.B1(n_565),
.B2(n_559),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_998),
.B(n_793),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1023),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1033),
.A2(n_781),
.B1(n_762),
.B2(n_649),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1023),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_998),
.B(n_794),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_979),
.B(n_731),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1023),
.B(n_796),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1030),
.Y(n_1173)
);

AND2x6_ASAP7_75t_L g1174 ( 
.A(n_1030),
.B(n_739),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1092),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1065),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1135),
.B(n_1004),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1065),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1046),
.A2(n_1030),
.B1(n_1021),
.B2(n_1029),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1041),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1046),
.A2(n_1029),
.B1(n_1014),
.B2(n_1005),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1107),
.B(n_837),
.Y(n_1182)
);

AO22x2_ASAP7_75t_L g1183 ( 
.A1(n_1074),
.A2(n_973),
.B1(n_749),
.B2(n_656),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1135),
.B(n_1032),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1041),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1127),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1082),
.B(n_959),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1060),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1088),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1111),
.A2(n_748),
.B1(n_668),
.B2(n_679),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1127),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1048),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1064),
.B(n_573),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1147),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1132),
.B(n_660),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1048),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1088),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1147),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1152),
.B(n_971),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1064),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_1145),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1060),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1050),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1050),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1141),
.B(n_695),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1147),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1172),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1147),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1093),
.A2(n_748),
.B1(n_715),
.B2(n_723),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1156),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_1113),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1141),
.B(n_710),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1164),
.B(n_840),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1069),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1054),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1164),
.B(n_842),
.Y(n_1217)
);

INVx4_ASAP7_75t_SL g1218 ( 
.A(n_1145),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1169),
.B(n_843),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1056),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1169),
.B(n_847),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1156),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1064),
.Y(n_1223)
);

AND2x2_ASAP7_75t_SL g1224 ( 
.A(n_1097),
.B(n_637),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1142),
.B(n_746),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1075),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1077),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1069),
.Y(n_1228)
);

BUFx4_ASAP7_75t_L g1229 ( 
.A(n_1144),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1167),
.B(n_848),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1064),
.B(n_1156),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1056),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1152),
.B(n_578),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1087),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1150),
.B(n_1119),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1085),
.B(n_782),
.C(n_732),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1156),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1087),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1142),
.B(n_747),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_L g1240 ( 
.A(n_1161),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1096),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1096),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1123),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1123),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1120),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1095),
.B(n_802),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1159),
.B(n_758),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1159),
.B(n_1160),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1130),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1119),
.B(n_578),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1137),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1161),
.B(n_850),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1123),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1136),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1071),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1160),
.B(n_759),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1071),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1093),
.A2(n_583),
.B1(n_594),
.B2(n_570),
.Y(n_1258)
);

AND2x2_ASAP7_75t_SL g1259 ( 
.A(n_1128),
.B(n_637),
.Y(n_1259)
);

AO22x2_ASAP7_75t_L g1260 ( 
.A1(n_1143),
.A2(n_749),
.B1(n_638),
.B2(n_648),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1079),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1044),
.B(n_804),
.Y(n_1262)
);

OR2x2_ASAP7_75t_SL g1263 ( 
.A(n_1106),
.B(n_638),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1047),
.B(n_595),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1080),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1095),
.B(n_616),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1163),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1122),
.B(n_596),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1058),
.B(n_618),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1081),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1076),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1076),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1123),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1104),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1105),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1089),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1090),
.Y(n_1277)
);

INVxp33_ASAP7_75t_L g1278 ( 
.A(n_1042),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1122),
.B(n_597),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1058),
.B(n_806),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1066),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1174),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1137),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1084),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1138),
.B(n_601),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1122),
.B(n_602),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1099),
.B(n_807),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1072),
.B(n_808),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1084),
.Y(n_1289)
);

INVx4_ASAP7_75t_SL g1290 ( 
.A(n_1174),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1163),
.B(n_858),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1149),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1146),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1091),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1138),
.B(n_620),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1094),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1070),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1134),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1126),
.Y(n_1299)
);

AND2x6_ASAP7_75t_L g1300 ( 
.A(n_1109),
.B(n_643),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1173),
.B(n_1140),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1045),
.B(n_612),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_L g1303 ( 
.A(n_1153),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1100),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1086),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1053),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1055),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1149),
.B(n_643),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1070),
.B(n_859),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1049),
.B(n_613),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1099),
.B(n_860),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1166),
.B(n_623),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1151),
.B(n_624),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1126),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1057),
.Y(n_1315)
);

INVx5_ASAP7_75t_L g1316 ( 
.A(n_1174),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1151),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1157),
.B(n_625),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1157),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1101),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1170),
.B(n_627),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1109),
.B(n_648),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1120),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1059),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1063),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1102),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1067),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1051),
.B(n_861),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1102),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1129),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1125),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1098),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1158),
.B(n_630),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1139),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1102),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1158),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1148),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1068),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1073),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1052),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1110),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1154),
.B(n_629),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1098),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1133),
.B(n_642),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1116),
.A2(n_653),
.B1(n_662),
.B2(n_647),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1117),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1118),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1155),
.B(n_576),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1168),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1121),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1120),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1165),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1124),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1174),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1171),
.B(n_863),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_R g1357 ( 
.A(n_1174),
.B(n_666),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1131),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1115),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1061),
.B(n_670),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1115),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1112),
.B(n_768),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1078),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1078),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1083),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1103),
.A2(n_779),
.B1(n_777),
.B2(n_725),
.C(n_640),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1112),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1083),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1043),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1162),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1114),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1108),
.B(n_768),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1133),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1245),
.B(n_1043),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1303),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1194),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_SL g1377 ( 
.A(n_1201),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1235),
.B(n_1114),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1259),
.B(n_1062),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1180),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1185),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1319),
.B(n_1062),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1359),
.B(n_866),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1337),
.B(n_673),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_634),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1188),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1361),
.B(n_866),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1278),
.B(n_639),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1175),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1197),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1365),
.B(n_866),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1202),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1189),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1234),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1344),
.B(n_646),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1368),
.B(n_681),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1179),
.B(n_685),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1297),
.B(n_686),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1367),
.B(n_691),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1215),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1297),
.B(n_1324),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1370),
.B(n_692),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1298),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1288),
.B(n_639),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1238),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1228),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1177),
.A2(n_700),
.B1(n_703),
.B2(n_693),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1262),
.B(n_705),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1255),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1257),
.Y(n_1411)
);

INVxp33_ASAP7_75t_L g1412 ( 
.A(n_1187),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1335),
.B(n_639),
.Y(n_1413)
);

NOR2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1353),
.B(n_834),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1184),
.B(n_655),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1186),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1220),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_L g1418 ( 
.A(n_1327),
.B(n_1330),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1207),
.A2(n_714),
.B1(n_727),
.B2(n_709),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1241),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1242),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1297),
.B(n_729),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1292),
.B(n_735),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1317),
.B(n_742),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1341),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1311),
.B(n_865),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1229),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1251),
.B(n_744),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1271),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1272),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1369),
.B(n_766),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1232),
.B(n_659),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1324),
.B(n_770),
.Y(n_1433)
);

AND2x6_ASAP7_75t_SL g1434 ( 
.A(n_1199),
.B(n_1266),
.Y(n_1434)
);

NOR3xp33_ASAP7_75t_L g1435 ( 
.A(n_1211),
.B(n_868),
.C(n_867),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1281),
.A2(n_772),
.B1(n_778),
.B2(n_774),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1371),
.B(n_879),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1201),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1371),
.B(n_885),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1342),
.B(n_886),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1283),
.B(n_667),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1209),
.A2(n_713),
.B1(n_871),
.B2(n_869),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1195),
.B(n_671),
.Y(n_1444)
);

AO221x1_ASAP7_75t_L g1445 ( 
.A1(n_1183),
.A2(n_874),
.B1(n_872),
.B2(n_880),
.C(n_672),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1327),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1194),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1226),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1366),
.B(n_1233),
.C(n_1264),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1194),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1193),
.A2(n_713),
.B1(n_674),
.B2(n_682),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1324),
.B(n_676),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1284),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1373),
.B(n_683),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1301),
.B(n_684),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1245),
.B(n_880),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_SL g1457 ( 
.A(n_1309),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1227),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1191),
.B(n_687),
.Y(n_1459)
);

OAI22x1_ASAP7_75t_R g1460 ( 
.A1(n_1332),
.A2(n_1350),
.B1(n_1338),
.B2(n_1249),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1305),
.B(n_688),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1312),
.A2(n_689),
.B1(n_697),
.B2(n_690),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1289),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1315),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1250),
.B(n_701),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1181),
.B(n_702),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1176),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1325),
.B(n_704),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1326),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1293),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1330),
.B(n_711),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1336),
.B(n_1322),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1352),
.B(n_1343),
.C(n_1360),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1287),
.B(n_717),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1340),
.B(n_720),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1218),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1336),
.B(n_721),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1318),
.B(n_722),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1190),
.A2(n_724),
.B1(n_733),
.B2(n_728),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1282),
.A2(n_880),
.B(n_694),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1240),
.B(n_737),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1280),
.B(n_738),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1304),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1269),
.B(n_672),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1246),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1321),
.B(n_741),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1328),
.A2(n_672),
.B1(n_745),
.B2(n_743),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1339),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1254),
.B(n_750),
.Y(n_1490)
);

INVx8_ASAP7_75t_L g1491 ( 
.A(n_1198),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1356),
.B(n_751),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1295),
.B(n_752),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1198),
.B(n_753),
.Y(n_1494)
);

OAI22x1_ASAP7_75t_L g1495 ( 
.A1(n_1219),
.A2(n_755),
.B1(n_757),
.B2(n_754),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_L g1496 ( 
.A(n_1349),
.B(n_761),
.C(n_760),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1198),
.B(n_763),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1219),
.B(n_775),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1214),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1309),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1214),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1268),
.A2(n_776),
.B(n_3),
.C(n_1),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1206),
.B(n_880),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1217),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1217),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1221),
.A2(n_880),
.B1(n_351),
.B2(n_352),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1276),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1248),
.B(n_350),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1206),
.B(n_353),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1261),
.B(n_356),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1265),
.B(n_360),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1206),
.B(n_363),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1270),
.B(n_366),
.Y(n_1513)
);

AO22x1_ASAP7_75t_L g1514 ( 
.A1(n_1223),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1294),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1218),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1221),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1308),
.B(n_1182),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1178),
.B(n_368),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1183),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.C(n_8),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1277),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1210),
.B(n_1222),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1308),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1296),
.B(n_370),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1329),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1252),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1192),
.B(n_372),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1224),
.B(n_7),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1182),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1230),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1196),
.B(n_373),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1210),
.B(n_375),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1203),
.B(n_376),
.Y(n_1533)
);

AND2x6_ASAP7_75t_SL g1534 ( 
.A(n_1372),
.B(n_8),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1230),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1210),
.B(n_378),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1252),
.B(n_9),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1299),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1291),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1291),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1204),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1212),
.B(n_379),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1216),
.B(n_380),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1299),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1279),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1372),
.B(n_13),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1314),
.B(n_382),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1347),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1314),
.B(n_383),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1357),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1351),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1222),
.B(n_384),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1222),
.B(n_385),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1286),
.B(n_14),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1320),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1320),
.B(n_386),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1331),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1302),
.B(n_15),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1258),
.A2(n_1310),
.B(n_1345),
.C(n_1354),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1331),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1205),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1313),
.B(n_1334),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1260),
.B(n_16),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1263),
.B(n_16),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1267),
.Y(n_1565)
);

INVx8_ASAP7_75t_L g1566 ( 
.A(n_1237),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1237),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1200),
.B(n_387),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1348),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1237),
.B(n_388),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1358),
.B(n_17),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1358),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1200),
.B(n_389),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1260),
.B(n_391),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1267),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1285),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1208),
.B(n_393),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1213),
.B(n_1225),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1346),
.B(n_17),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1426),
.B(n_1239),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1491),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1525),
.B(n_1208),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1389),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1465),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1449),
.A2(n_1247),
.B(n_1256),
.C(n_1231),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1404),
.B(n_1243),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1375),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1470),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1466),
.B(n_1236),
.Y(n_1589)
);

INVx8_ASAP7_75t_L g1590 ( 
.A(n_1491),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1491),
.B(n_1243),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1436),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1415),
.B(n_1300),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1416),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1425),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1391),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1578),
.A2(n_1316),
.B(n_1282),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1405),
.B(n_1300),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_R g1599 ( 
.A(n_1477),
.B(n_1282),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1507),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1479),
.B(n_1300),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1412),
.B(n_1243),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1474),
.A2(n_1323),
.B1(n_1362),
.B2(n_1300),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1436),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1471),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1394),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1379),
.B(n_1323),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1579),
.A2(n_1362),
.B1(n_1323),
.B2(n_1355),
.Y(n_1610)
);

AND2x6_ASAP7_75t_L g1611 ( 
.A(n_1577),
.B(n_1355),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1483),
.B(n_1244),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1439),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1528),
.A2(n_1362),
.B1(n_1323),
.B2(n_1355),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1417),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1475),
.B(n_1362),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1566),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1486),
.B(n_1244),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1432),
.B(n_1244),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1564),
.B(n_18),
.C(n_19),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1550),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1492),
.B(n_1253),
.Y(n_1623)
);

AND2x6_ASAP7_75t_L g1624 ( 
.A(n_1577),
.B(n_1253),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1517),
.B(n_1253),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_R g1626 ( 
.A(n_1516),
.B(n_1273),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1446),
.B(n_1273),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1455),
.B(n_1273),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1529),
.B(n_1518),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1485),
.A2(n_1558),
.B1(n_1554),
.B2(n_1493),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1435),
.B(n_1316),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1500),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1462),
.A2(n_1316),
.B1(n_1290),
.B2(n_22),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1460),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_SL g1635 ( 
.A(n_1496),
.B(n_1290),
.C(n_19),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_SL g1636 ( 
.A(n_1520),
.B(n_20),
.C(n_22),
.Y(n_1636)
);

AND2x6_ASAP7_75t_L g1637 ( 
.A(n_1446),
.B(n_396),
.Y(n_1637)
);

NOR3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1467),
.B(n_20),
.C(n_23),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1377),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1455),
.B(n_23),
.Y(n_1640)
);

AND2x6_ASAP7_75t_SL g1641 ( 
.A(n_1385),
.B(n_24),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1562),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1454),
.B(n_25),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1484),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1444),
.B(n_26),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1561),
.B(n_27),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1448),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1526),
.B(n_397),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1396),
.B(n_27),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1403),
.B(n_1390),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1458),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1427),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1523),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1413),
.B(n_28),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1403),
.B(n_29),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1489),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1414),
.Y(n_1657)
);

NOR2x1p5_ASAP7_75t_SL g1658 ( 
.A(n_1380),
.B(n_399),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1381),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1530),
.B(n_30),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1498),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1535),
.B(n_1499),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1501),
.B(n_31),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1454),
.B(n_1461),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1384),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1457),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1390),
.B(n_33),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1565),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1395),
.Y(n_1669)
);

INVx6_ASAP7_75t_L g1670 ( 
.A(n_1434),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1409),
.B(n_34),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1441),
.B(n_34),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1406),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1420),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1537),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1565),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_SL g1677 ( 
.A(n_1376),
.B(n_1450),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1441),
.B(n_35),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1504),
.B(n_401),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1505),
.B(n_35),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1388),
.B(n_36),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1418),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1457),
.B(n_402),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1421),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1386),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1572),
.B(n_37),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1376),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1576),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1450),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1548),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1567),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1393),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1382),
.B(n_39),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1459),
.A2(n_45),
.B1(n_41),
.B2(n_43),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1539),
.A2(n_1540),
.B1(n_1488),
.B2(n_1495),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1438),
.B(n_43),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1551),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1559),
.A2(n_405),
.B(n_404),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1567),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1452),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1438),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1440),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1571),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1401),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1515),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1546),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1440),
.B(n_48),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1575),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1378),
.B(n_49),
.Y(n_1709)
);

AND2x6_ASAP7_75t_L g1710 ( 
.A(n_1563),
.B(n_406),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1456),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1378),
.B(n_1397),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1407),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1397),
.B(n_49),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1410),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1411),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1429),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1430),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1453),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1490),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1464),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1469),
.B(n_51),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1569),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1456),
.B(n_1472),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1541),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1456),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1574),
.B(n_1538),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1544),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1383),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1476),
.B(n_52),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1374),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1408),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1377),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1437),
.B(n_53),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1442),
.B(n_55),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1383),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1402),
.Y(n_1737)
);

INVx5_ASAP7_75t_L g1738 ( 
.A(n_1374),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1374),
.B(n_552),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1482),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1555),
.Y(n_1741)
);

BUFx4f_ASAP7_75t_L g1742 ( 
.A(n_1557),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1560),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1494),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1468),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1387),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_R g1747 ( 
.A(n_1568),
.B(n_407),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1387),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1445),
.A2(n_61),
.B1(n_57),
.B2(n_60),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1487),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1423),
.B(n_63),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1522),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1398),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1392),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1480),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1392),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1400),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1480),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1534),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1424),
.B(n_68),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1428),
.B(n_70),
.Y(n_1761)
);

AND3x2_ASAP7_75t_SL g1762 ( 
.A(n_1514),
.B(n_71),
.C(n_72),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1400),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1463),
.B(n_71),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1510),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1431),
.B(n_73),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1510),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1431),
.B(n_73),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1497),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1508),
.A2(n_409),
.B(n_408),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1511),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1447),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1524),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1630),
.B(n_1473),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_L g1775 ( 
.A(n_1611),
.B(n_1511),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1650),
.B(n_1513),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1592),
.B(n_1443),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1664),
.B(n_1419),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1623),
.B(n_1513),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1589),
.B(n_1399),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1757),
.B(n_1422),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1605),
.B(n_1451),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1649),
.B(n_1502),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1763),
.B(n_1478),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1750),
.B(n_1524),
.Y(n_1785)
);

NAND2xp33_ASAP7_75t_SL g1786 ( 
.A(n_1626),
.B(n_1574),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1580),
.B(n_1433),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1769),
.B(n_1506),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1701),
.B(n_1519),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1615),
.B(n_1519),
.Y(n_1790)
);

NAND2xp33_ASAP7_75t_SL g1791 ( 
.A(n_1607),
.B(n_1527),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1702),
.B(n_1712),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1655),
.B(n_1740),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1628),
.B(n_1527),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1598),
.B(n_1531),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1734),
.B(n_1531),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1612),
.B(n_1533),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1617),
.B(n_1533),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1634),
.B(n_1542),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1751),
.B(n_1542),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1739),
.B(n_1509),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1739),
.B(n_1543),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1640),
.B(n_1543),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1714),
.B(n_1568),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1766),
.B(n_1573),
.Y(n_1805)
);

NAND2xp33_ASAP7_75t_SL g1806 ( 
.A(n_1638),
.B(n_1573),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_SL g1807 ( 
.A(n_1665),
.B(n_1512),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1731),
.B(n_1570),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1768),
.B(n_1593),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1731),
.B(n_1508),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1583),
.B(n_1532),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1731),
.B(n_1547),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1738),
.B(n_1547),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1672),
.B(n_1545),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1738),
.B(n_1549),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1738),
.B(n_1549),
.Y(n_1816)
);

NAND2xp33_ASAP7_75t_R g1817 ( 
.A(n_1622),
.B(n_1556),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1695),
.B(n_1556),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1645),
.B(n_1536),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1646),
.B(n_1552),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1724),
.B(n_1553),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1722),
.B(n_1481),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1730),
.B(n_1503),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1678),
.B(n_1765),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1671),
.B(n_1643),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1620),
.B(n_74),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1767),
.B(n_74),
.Y(n_1827)
);

NAND2xp33_ASAP7_75t_SL g1828 ( 
.A(n_1581),
.B(n_75),
.Y(n_1828)
);

NAND2xp33_ASAP7_75t_SL g1829 ( 
.A(n_1581),
.B(n_75),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1581),
.B(n_76),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1771),
.B(n_76),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1679),
.B(n_77),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1679),
.B(n_79),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1629),
.B(n_80),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1629),
.B(n_81),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1760),
.B(n_81),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1761),
.B(n_82),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1675),
.B(n_82),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1596),
.B(n_83),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1681),
.B(n_1706),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1735),
.B(n_83),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1742),
.B(n_84),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1742),
.B(n_1595),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1746),
.B(n_84),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1773),
.B(n_85),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1667),
.B(n_85),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1754),
.B(n_87),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1618),
.B(n_87),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1729),
.B(n_88),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1696),
.B(n_88),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1618),
.B(n_89),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1707),
.B(n_89),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1693),
.B(n_90),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1764),
.B(n_90),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1648),
.B(n_91),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1621),
.B(n_92),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1648),
.B(n_92),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1752),
.B(n_93),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1752),
.B(n_93),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1752),
.B(n_94),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1736),
.B(n_95),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1748),
.B(n_96),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1683),
.B(n_97),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1756),
.B(n_97),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1632),
.B(n_98),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1737),
.B(n_98),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1584),
.B(n_100),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_SL g1868 ( 
.A(n_1618),
.B(n_101),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1588),
.B(n_101),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1600),
.B(n_102),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1616),
.B(n_102),
.Y(n_1871)
);

NAND2xp33_ASAP7_75t_SL g1872 ( 
.A(n_1587),
.B(n_103),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1631),
.B(n_103),
.Y(n_1873)
);

NAND2xp33_ASAP7_75t_SL g1874 ( 
.A(n_1606),
.B(n_104),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1709),
.B(n_1644),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1747),
.B(n_104),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1586),
.B(n_105),
.Y(n_1877)
);

AND3x1_ASAP7_75t_L g1878 ( 
.A(n_1657),
.B(n_106),
.C(n_107),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1656),
.B(n_106),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1723),
.B(n_1594),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1609),
.B(n_107),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1602),
.B(n_109),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1614),
.B(n_110),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1715),
.B(n_111),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1713),
.B(n_410),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1745),
.B(n_111),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1717),
.B(n_1718),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1721),
.B(n_112),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1610),
.B(n_112),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1772),
.B(n_113),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1728),
.B(n_1743),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1705),
.B(n_113),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1654),
.B(n_114),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1603),
.B(n_114),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1585),
.B(n_115),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1713),
.B(n_412),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1659),
.B(n_1685),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1692),
.B(n_116),
.Y(n_1898)
);

NAND2xp33_ASAP7_75t_SL g1899 ( 
.A(n_1601),
.B(n_118),
.Y(n_1899)
);

NAND2xp33_ASAP7_75t_SL g1900 ( 
.A(n_1601),
.B(n_118),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1759),
.B(n_414),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1704),
.B(n_1716),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1719),
.B(n_119),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1708),
.B(n_120),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1608),
.B(n_120),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1759),
.B(n_417),
.Y(n_1906)
);

NAND2xp33_ASAP7_75t_SL g1907 ( 
.A(n_1608),
.B(n_121),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1708),
.B(n_121),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_SL g1909 ( 
.A(n_1677),
.B(n_122),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1604),
.B(n_124),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1639),
.B(n_125),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1661),
.B(n_126),
.Y(n_1912)
);

NAND2xp33_ASAP7_75t_SL g1913 ( 
.A(n_1733),
.B(n_127),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1647),
.B(n_130),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1651),
.B(n_130),
.Y(n_1915)
);

NAND2xp33_ASAP7_75t_SL g1916 ( 
.A(n_1666),
.B(n_131),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1690),
.B(n_131),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1697),
.B(n_132),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1669),
.B(n_132),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1673),
.B(n_133),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1674),
.B(n_133),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1758),
.B(n_134),
.Y(n_1922)
);

NAND2xp33_ASAP7_75t_SL g1923 ( 
.A(n_1689),
.B(n_134),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1684),
.B(n_135),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_SL g1925 ( 
.A(n_1689),
.B(n_135),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1725),
.B(n_136),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1689),
.B(n_137),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1662),
.B(n_137),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1582),
.B(n_138),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1619),
.B(n_138),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1694),
.B(n_139),
.Y(n_1931)
);

NAND2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1652),
.B(n_1726),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1660),
.B(n_140),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1711),
.B(n_1633),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1597),
.B(n_141),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1686),
.B(n_141),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1663),
.B(n_142),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1732),
.B(n_142),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1680),
.B(n_144),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1653),
.B(n_144),
.Y(n_1940)
);

NAND2xp33_ASAP7_75t_SL g1941 ( 
.A(n_1703),
.B(n_145),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1741),
.B(n_145),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1700),
.B(n_146),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1670),
.B(n_418),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1688),
.B(n_147),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1817),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1885),
.Y(n_1947)
);

O2A1O1Ixp33_ASAP7_75t_L g1948 ( 
.A1(n_1783),
.A2(n_1642),
.B(n_1636),
.C(n_1635),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1793),
.B(n_1778),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1843),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1880),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1786),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1887),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1840),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1891),
.Y(n_1955)
);

O2A1O1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1796),
.A2(n_1770),
.B(n_1698),
.C(n_1755),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1792),
.B(n_1727),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1824),
.B(n_1727),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1897),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1788),
.B(n_1670),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1902),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1790),
.B(n_1749),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1886),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1797),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1885),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1875),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1844),
.Y(n_1967)
);

AOI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1895),
.A2(n_1591),
.B(n_1625),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1776),
.B(n_1727),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1885),
.Y(n_1970)
);

OR2x6_ASAP7_75t_L g1971 ( 
.A(n_1810),
.B(n_1812),
.Y(n_1971)
);

OR2x6_ASAP7_75t_L g1972 ( 
.A(n_1813),
.B(n_1658),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1784),
.Y(n_1973)
);

NOR2x1_ASAP7_75t_SL g1974 ( 
.A(n_1815),
.B(n_1591),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1910),
.A2(n_1753),
.B1(n_1720),
.B2(n_1744),
.Y(n_1975)
);

AOI221xp5_ASAP7_75t_L g1976 ( 
.A1(n_1941),
.A2(n_1762),
.B1(n_1641),
.B2(n_1613),
.C(n_1590),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1896),
.Y(n_1977)
);

NOR2xp67_ASAP7_75t_L g1978 ( 
.A(n_1811),
.B(n_1687),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1910),
.A2(n_1625),
.B1(n_1676),
.B2(n_1668),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1856),
.B(n_1710),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1801),
.Y(n_1981)
);

CKINVDCx11_ASAP7_75t_R g1982 ( 
.A(n_1801),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1775),
.A2(n_1682),
.B(n_1676),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1776),
.B(n_1727),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1847),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1854),
.A2(n_1668),
.B1(n_1710),
.B2(n_1691),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1896),
.Y(n_1987)
);

AO21x2_ASAP7_75t_L g1988 ( 
.A1(n_1798),
.A2(n_1710),
.B(n_1627),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1896),
.Y(n_1989)
);

CKINVDCx8_ASAP7_75t_R g1990 ( 
.A(n_1801),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1808),
.B(n_1687),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1849),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1861),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1782),
.B(n_1710),
.Y(n_1994)
);

O2A1O1Ixp5_ASAP7_75t_L g1995 ( 
.A1(n_1818),
.A2(n_1682),
.B(n_1699),
.C(n_1691),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1825),
.B(n_1699),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1785),
.B(n_1637),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1791),
.B(n_1590),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1938),
.A2(n_1637),
.B1(n_1611),
.B2(n_1624),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1808),
.B(n_1624),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1862),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1922),
.B(n_1637),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1779),
.B(n_1624),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1943),
.A2(n_1611),
.B1(n_1624),
.B2(n_1637),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1864),
.Y(n_2005)
);

BUFx4f_ASAP7_75t_L g2006 ( 
.A(n_1808),
.Y(n_2006)
);

INVx4_ASAP7_75t_L g2007 ( 
.A(n_1838),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1802),
.A2(n_1599),
.B(n_1611),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1781),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1809),
.B(n_147),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1800),
.B(n_1627),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1921),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1799),
.Y(n_2014)
);

INVxp67_ASAP7_75t_L g2015 ( 
.A(n_1865),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1931),
.Y(n_2016)
);

INVx4_ASAP7_75t_L g2017 ( 
.A(n_1945),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1944),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1926),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1787),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1780),
.B(n_419),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_1774),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1876),
.B(n_420),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1804),
.B(n_1627),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1912),
.A2(n_1627),
.B1(n_150),
.B2(n_148),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1789),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1937),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1777),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1816),
.Y(n_2029)
);

AOI21xp33_ASAP7_75t_L g2030 ( 
.A1(n_1814),
.A2(n_148),
.B(n_149),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1878),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1794),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1845),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1827),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1901),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1831),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1846),
.B(n_1850),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1853),
.B(n_421),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1823),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1863),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1774),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2041)
);

O2A1O1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1836),
.A2(n_155),
.B(n_152),
.C(n_154),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1858),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1821),
.Y(n_2044)
);

AOI21xp33_ASAP7_75t_L g2045 ( 
.A1(n_1803),
.A2(n_154),
.B(n_155),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1884),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1888),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1879),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1855),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1805),
.A2(n_423),
.B(n_422),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1934),
.B(n_424),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1807),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1906),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1837),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1806),
.B(n_425),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1898),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1932),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1882),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1852),
.B(n_160),
.Y(n_2059)
);

OR2x6_ASAP7_75t_L g2060 ( 
.A(n_1795),
.B(n_427),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_1935),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1881),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1867),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1903),
.Y(n_2064)
);

A2O1A1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_1909),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1951),
.B(n_1841),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_1948),
.A2(n_1916),
.B(n_1828),
.C(n_1830),
.Y(n_2067)
);

O2A1O1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_1975),
.A2(n_1842),
.B(n_1857),
.C(n_1866),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1973),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1956),
.A2(n_1829),
.B(n_1851),
.C(n_1848),
.Y(n_2070)
);

OAI22x1_ASAP7_75t_L g2071 ( 
.A1(n_1946),
.A2(n_1940),
.B1(n_1890),
.B2(n_1859),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1975),
.A2(n_1822),
.B(n_1819),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_2035),
.B(n_1839),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_1983),
.A2(n_1820),
.B(n_1904),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2057),
.A2(n_1883),
.B1(n_1832),
.B2(n_1833),
.Y(n_2075)
);

AO31x2_ASAP7_75t_L g2076 ( 
.A1(n_1974),
.A2(n_1899),
.A3(n_1905),
.B(n_1900),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1954),
.Y(n_2077)
);

AOI221xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2049),
.A2(n_1893),
.B1(n_1860),
.B2(n_1915),
.C(n_1914),
.Y(n_2078)
);

OAI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1995),
.A2(n_1908),
.B(n_1928),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_1969),
.A2(n_1870),
.B(n_1869),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1949),
.A2(n_1868),
.B1(n_1925),
.B2(n_1923),
.Y(n_2081)
);

INVx6_ASAP7_75t_SL g2082 ( 
.A(n_1971),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_1950),
.Y(n_2083)
);

BUFx8_ASAP7_75t_SL g2084 ( 
.A(n_2018),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_1969),
.A2(n_1871),
.B(n_1826),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2053),
.B(n_1834),
.Y(n_2086)
);

CKINVDCx11_ASAP7_75t_R g2087 ( 
.A(n_2007),
.Y(n_2087)
);

INVx3_ASAP7_75t_SL g2088 ( 
.A(n_2007),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1953),
.Y(n_2089)
);

O2A1O1Ixp33_ASAP7_75t_SL g2090 ( 
.A1(n_2065),
.A2(n_1873),
.B(n_1918),
.C(n_1917),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1964),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1951),
.B(n_1966),
.Y(n_2092)
);

AOI21x1_ASAP7_75t_L g2093 ( 
.A1(n_1962),
.A2(n_1920),
.B(n_1919),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_2006),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2016),
.B(n_1924),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2021),
.A2(n_1936),
.B(n_1933),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_2042),
.A2(n_1927),
.B(n_1907),
.C(n_1874),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_1982),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2032),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2029),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1981),
.B(n_1835),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1955),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2009),
.Y(n_2103)
);

A2O1A1Ixp33_ASAP7_75t_L g2104 ( 
.A1(n_2054),
.A2(n_1911),
.B(n_1913),
.C(n_1872),
.Y(n_2104)
);

OR2x6_ASAP7_75t_L g2105 ( 
.A(n_1971),
.B(n_1889),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2028),
.B(n_1894),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2016),
.B(n_1877),
.Y(n_2107)
);

OA21x2_ASAP7_75t_L g2108 ( 
.A1(n_1984),
.A2(n_1930),
.B(n_1929),
.Y(n_2108)
);

AO31x2_ASAP7_75t_L g2109 ( 
.A1(n_1979),
.A2(n_1939),
.A3(n_1892),
.B(n_166),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2061),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2026),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1960),
.A2(n_168),
.B1(n_164),
.B2(n_167),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2004),
.A2(n_429),
.B(n_428),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2004),
.A2(n_431),
.B(n_430),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_L g2115 ( 
.A1(n_1984),
.A2(n_433),
.B(n_432),
.Y(n_2115)
);

A2O1A1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_2052),
.A2(n_170),
.B(n_167),
.C(n_169),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2060),
.A2(n_436),
.B(n_435),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_1957),
.A2(n_438),
.B(n_437),
.Y(n_2118)
);

A2O1A1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_2023),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_SL g2120 ( 
.A(n_1952),
.B(n_442),
.Y(n_2120)
);

AO31x2_ASAP7_75t_L g2121 ( 
.A1(n_1979),
.A2(n_175),
.A3(n_173),
.B(n_174),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2049),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2122)
);

OAI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_2055),
.A2(n_445),
.B(n_444),
.Y(n_2123)
);

NAND3xp33_ASAP7_75t_L g2124 ( 
.A(n_2041),
.B(n_176),
.C(n_177),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_2060),
.A2(n_450),
.B(n_448),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1957),
.A2(n_453),
.B(n_451),
.Y(n_2126)
);

AO31x2_ASAP7_75t_L g2127 ( 
.A1(n_1986),
.A2(n_178),
.A3(n_176),
.B(n_177),
.Y(n_2127)
);

AO31x2_ASAP7_75t_L g2128 ( 
.A1(n_1986),
.A2(n_180),
.A3(n_178),
.B(n_179),
.Y(n_2128)
);

BUFx2_ASAP7_75t_R g2129 ( 
.A(n_1990),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_1991),
.B(n_455),
.Y(n_2130)
);

AO31x2_ASAP7_75t_L g2131 ( 
.A1(n_1958),
.A2(n_182),
.A3(n_179),
.B(n_181),
.Y(n_2131)
);

AO32x2_ASAP7_75t_L g2132 ( 
.A1(n_2017),
.A2(n_185),
.A3(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_R g2133 ( 
.A(n_2031),
.B(n_457),
.Y(n_2133)
);

OAI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_2050),
.A2(n_459),
.B(n_458),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1947),
.B(n_460),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1958),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2039),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1993),
.B(n_183),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2040),
.A2(n_463),
.B(n_461),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1950),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1967),
.B(n_185),
.Y(n_2141)
);

OAI21x1_ASAP7_75t_L g2142 ( 
.A1(n_2074),
.A2(n_1968),
.B(n_2024),
.Y(n_2142)
);

OA21x2_ASAP7_75t_L g2143 ( 
.A1(n_2072),
.A2(n_1994),
.B(n_2022),
.Y(n_2143)
);

CKINVDCx6p67_ASAP7_75t_R g2144 ( 
.A(n_2087),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_SL g2145 ( 
.A1(n_2093),
.A2(n_2044),
.B(n_1997),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2069),
.Y(n_2146)
);

OAI21x1_ASAP7_75t_L g2147 ( 
.A1(n_2115),
.A2(n_2024),
.B(n_2008),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_L g2148 ( 
.A1(n_2118),
.A2(n_2003),
.B(n_1998),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2091),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_2088),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2089),
.Y(n_2151)
);

CKINVDCx6p67_ASAP7_75t_R g2152 ( 
.A(n_2098),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2136),
.B(n_2020),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2092),
.B(n_2020),
.Y(n_2154)
);

OAI21x1_ASAP7_75t_L g2155 ( 
.A1(n_2126),
.A2(n_2003),
.B(n_2012),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_2103),
.B(n_1971),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2080),
.A2(n_2061),
.B(n_1965),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2099),
.Y(n_2158)
);

AOI221xp5_ASAP7_75t_L g2159 ( 
.A1(n_2122),
.A2(n_2119),
.B1(n_2040),
.B2(n_2068),
.C(n_2116),
.Y(n_2159)
);

BUFx10_ASAP7_75t_L g2160 ( 
.A(n_2073),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2100),
.B(n_1988),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2102),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2111),
.B(n_1988),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_2085),
.A2(n_1965),
.B(n_1947),
.Y(n_2164)
);

CKINVDCx20_ASAP7_75t_R g2165 ( 
.A(n_2084),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_2079),
.A2(n_2022),
.B(n_2030),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2137),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2095),
.B(n_2010),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_2082),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2066),
.B(n_1992),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2131),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_SL g2172 ( 
.A1(n_2139),
.A2(n_2037),
.B(n_2036),
.Y(n_2172)
);

OAI21x1_ASAP7_75t_L g2173 ( 
.A1(n_2113),
.A2(n_2114),
.B(n_2117),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2140),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_2125),
.A2(n_1977),
.B(n_1970),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2134),
.A2(n_2060),
.B(n_2006),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2131),
.Y(n_2177)
);

OAI21x1_ASAP7_75t_L g2178 ( 
.A1(n_2108),
.A2(n_1977),
.B(n_1970),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2140),
.Y(n_2179)
);

OAI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2067),
.A2(n_2030),
.B(n_2045),
.Y(n_2180)
);

OAI22x1_ASAP7_75t_L g2181 ( 
.A1(n_2112),
.A2(n_2031),
.B1(n_2014),
.B2(n_2081),
.Y(n_2181)
);

BUFx12f_ASAP7_75t_L g2182 ( 
.A(n_2130),
.Y(n_2182)
);

AO21x2_ASAP7_75t_L g2183 ( 
.A1(n_2096),
.A2(n_2045),
.B(n_1978),
.Y(n_2183)
);

AOI21x1_ASAP7_75t_L g2184 ( 
.A1(n_2071),
.A2(n_1980),
.B(n_2001),
.Y(n_2184)
);

BUFx3_ASAP7_75t_L g2185 ( 
.A(n_2077),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2121),
.Y(n_2186)
);

OAI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2070),
.A2(n_1952),
.B(n_2059),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2123),
.A2(n_1972),
.B(n_1987),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2151),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2146),
.B(n_2083),
.Y(n_2190)
);

AOI22xp33_ASAP7_75t_L g2191 ( 
.A1(n_2159),
.A2(n_2124),
.B1(n_2075),
.B2(n_2025),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_2180),
.A2(n_2110),
.B1(n_2051),
.B2(n_2105),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2153),
.B(n_2154),
.Y(n_2193)
);

OR2x6_ASAP7_75t_L g2194 ( 
.A(n_2188),
.B(n_2105),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2176),
.A2(n_2097),
.B1(n_2104),
.B2(n_2082),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2187),
.A2(n_1999),
.B1(n_2129),
.B2(n_2086),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2149),
.B(n_2101),
.Y(n_2197)
);

AO31x2_ASAP7_75t_L g2198 ( 
.A1(n_2186),
.A2(n_2177),
.A3(n_2171),
.B(n_2151),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_2181),
.A2(n_2051),
.B1(n_2183),
.B2(n_2172),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2153),
.B(n_2015),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2158),
.Y(n_2201)
);

INVxp67_ASAP7_75t_SL g2202 ( 
.A(n_2149),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2168),
.B(n_2121),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2167),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2177),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2181),
.A2(n_2062),
.B1(n_2058),
.B2(n_2034),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2162),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2183),
.A2(n_2047),
.B1(n_2046),
.B2(n_2063),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_2150),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2156),
.B(n_2107),
.Y(n_2210)
);

INVx1_ASAP7_75t_SL g2211 ( 
.A(n_2152),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2186),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2201),
.Y(n_2213)
);

AOI222xp33_ASAP7_75t_L g2214 ( 
.A1(n_2191),
.A2(n_1976),
.B1(n_1985),
.B2(n_2005),
.C1(n_2019),
.C2(n_2013),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2210),
.B(n_2161),
.Y(n_2215)
);

INVx2_ASAP7_75t_SL g2216 ( 
.A(n_2209),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2198),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2191),
.A2(n_2144),
.B1(n_2169),
.B2(n_2184),
.Y(n_2218)
);

AO31x2_ASAP7_75t_L g2219 ( 
.A1(n_2212),
.A2(n_2170),
.A3(n_2141),
.B(n_2138),
.Y(n_2219)
);

OAI221xp5_ASAP7_75t_L g2220 ( 
.A1(n_2199),
.A2(n_2169),
.B1(n_2078),
.B2(n_2150),
.C(n_2043),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_2195),
.A2(n_2173),
.B1(n_2156),
.B2(n_2145),
.Y(n_2221)
);

OR2x6_ASAP7_75t_L g2222 ( 
.A(n_2209),
.B(n_2169),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2202),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_R g2224 ( 
.A(n_2216),
.B(n_2165),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2213),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2219),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2217),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_2222),
.Y(n_2228)
);

XNOR2xp5_ASAP7_75t_L g2229 ( 
.A(n_2218),
.B(n_2211),
.Y(n_2229)
);

INVxp67_ASAP7_75t_L g2230 ( 
.A(n_2222),
.Y(n_2230)
);

NAND2xp33_ASAP7_75t_R g2231 ( 
.A(n_2215),
.B(n_2133),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2230),
.B(n_2228),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2228),
.B(n_2215),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2225),
.Y(n_2234)
);

NOR2x1_ASAP7_75t_L g2235 ( 
.A(n_2229),
.B(n_2165),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2224),
.B(n_2223),
.Y(n_2236)
);

AO31x2_ASAP7_75t_L g2237 ( 
.A1(n_2227),
.A2(n_2205),
.A3(n_2196),
.B(n_2204),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_2225),
.B(n_2209),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2226),
.B(n_2219),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2227),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2229),
.B(n_2207),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2236),
.B(n_2144),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2235),
.A2(n_2220),
.B1(n_2194),
.B2(n_2199),
.Y(n_2243)
);

NAND4xp25_ASAP7_75t_L g2244 ( 
.A(n_2232),
.B(n_2214),
.C(n_2221),
.D(n_2206),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2238),
.B(n_2200),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2238),
.B(n_2206),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2233),
.B(n_2209),
.Y(n_2247)
);

NAND3xp33_ASAP7_75t_SL g2248 ( 
.A(n_2241),
.B(n_2208),
.C(n_2192),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2239),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2241),
.A2(n_2208),
.B(n_2192),
.Y(n_2250)
);

NAND4xp25_ASAP7_75t_L g2251 ( 
.A(n_2234),
.B(n_2231),
.C(n_2185),
.D(n_2120),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2237),
.B(n_2160),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2237),
.B(n_2160),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2242),
.B(n_2237),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2247),
.B(n_2237),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_2249),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2245),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2246),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2243),
.A2(n_2194),
.B1(n_2152),
.B2(n_2240),
.Y(n_2259)
);

AO21x2_ASAP7_75t_L g2260 ( 
.A1(n_2248),
.A2(n_2011),
.B(n_2132),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_2250),
.B(n_2185),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2252),
.B(n_2210),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2254),
.B(n_2253),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2256),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2254),
.B(n_2197),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2257),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2264),
.B(n_2258),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2263),
.B(n_2261),
.Y(n_2268)
);

NAND4xp25_ASAP7_75t_L g2269 ( 
.A(n_2266),
.B(n_2261),
.C(n_2259),
.D(n_2262),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2263),
.B(n_2261),
.Y(n_2270)
);

AO221x2_ASAP7_75t_L g2271 ( 
.A1(n_2268),
.A2(n_2251),
.B1(n_2260),
.B2(n_2244),
.C(n_2262),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2270),
.B(n_2265),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2267),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2269),
.B(n_2265),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2267),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_SL g2276 ( 
.A(n_2268),
.B(n_2255),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2272),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2274),
.B(n_2260),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2275),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2273),
.B(n_2255),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2271),
.B(n_2193),
.Y(n_2281)
);

AND3x2_ASAP7_75t_L g2282 ( 
.A(n_2276),
.B(n_2038),
.C(n_2094),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2275),
.B(n_2160),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2275),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_2272),
.B(n_2194),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2272),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_2281),
.B(n_2190),
.Y(n_2287)
);

OR2x2_ASAP7_75t_L g2288 ( 
.A(n_2278),
.B(n_2203),
.Y(n_2288)
);

INVxp67_ASAP7_75t_SL g2289 ( 
.A(n_2280),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2279),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2284),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2277),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2282),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2277),
.B(n_2189),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_2283),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2286),
.B(n_2143),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2285),
.B(n_2198),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2280),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2280),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2289),
.B(n_2198),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2299),
.B(n_2198),
.Y(n_2301)
);

OAI221xp5_ASAP7_75t_SL g2302 ( 
.A1(n_2293),
.A2(n_2027),
.B1(n_2132),
.B2(n_1996),
.C(n_2106),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2287),
.A2(n_2174),
.B1(n_2179),
.B2(n_2182),
.Y(n_2303)
);

OAI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2290),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2304)
);

OAI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2298),
.A2(n_2179),
.B1(n_2174),
.B2(n_2182),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2291),
.Y(n_2306)
);

OAI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2295),
.A2(n_2090),
.B1(n_2166),
.B2(n_2033),
.C(n_1963),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2288),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2295),
.A2(n_2132),
.B1(n_2135),
.B2(n_2205),
.C(n_2161),
.Y(n_2309)
);

INVxp67_ASAP7_75t_L g2310 ( 
.A(n_2292),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2294),
.B(n_188),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2296),
.B(n_2156),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2297),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2297),
.B(n_190),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2311),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2304),
.Y(n_2316)
);

OAI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2310),
.A2(n_2173),
.B(n_2142),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2306),
.B(n_2143),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2308),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2303),
.B(n_2143),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2314),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2312),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2305),
.B(n_2174),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2313),
.B(n_2142),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2309),
.B(n_2300),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2301),
.B(n_2166),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2307),
.Y(n_2327)
);

AOI21xp33_ASAP7_75t_SL g2328 ( 
.A1(n_2302),
.A2(n_190),
.B(n_191),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2319),
.Y(n_2329)
);

O2A1O1Ixp33_ASAP7_75t_L g2330 ( 
.A1(n_2316),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_2330)
);

XNOR2xp5_ASAP7_75t_L g2331 ( 
.A(n_2322),
.B(n_192),
.Y(n_2331)
);

AOI322xp5_ASAP7_75t_L g2332 ( 
.A1(n_2327),
.A2(n_2002),
.A3(n_2161),
.B1(n_2135),
.B2(n_2056),
.C1(n_2064),
.C2(n_2048),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2315),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2321),
.B(n_2174),
.Y(n_2334)
);

AO22x2_ASAP7_75t_L g2335 ( 
.A1(n_2325),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.Y(n_2335)
);

NAND4xp25_ASAP7_75t_L g2336 ( 
.A(n_2323),
.B(n_198),
.C(n_196),
.D(n_197),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2318),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2328),
.B(n_198),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2324),
.Y(n_2339)
);

AOI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_2320),
.A2(n_2179),
.B1(n_2166),
.B2(n_1950),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2326),
.B(n_2076),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2317),
.Y(n_2342)
);

AOI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_2317),
.A2(n_199),
.B(n_200),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_2319),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_2319),
.Y(n_2345)
);

AOI221x1_ASAP7_75t_SL g2346 ( 
.A1(n_2316),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2319),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2319),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2319),
.B(n_2179),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2319),
.A2(n_201),
.B(n_203),
.Y(n_2350)
);

INVx2_ASAP7_75t_SL g2351 ( 
.A(n_2349),
.Y(n_2351)
);

INVxp33_ASAP7_75t_SL g2352 ( 
.A(n_2331),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2336),
.B(n_203),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2335),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2344),
.B(n_204),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2335),
.Y(n_2356)
);

INVx1_ASAP7_75t_SL g2357 ( 
.A(n_2338),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2346),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_2350),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2334),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2330),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2329),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2347),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2348),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2333),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2345),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2337),
.Y(n_2367)
);

INVx3_ASAP7_75t_SL g2368 ( 
.A(n_2339),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2342),
.Y(n_2369)
);

CKINVDCx6p67_ASAP7_75t_R g2370 ( 
.A(n_2341),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2343),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2341),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2340),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2332),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2346),
.B(n_205),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2335),
.Y(n_2376)
);

INVxp33_ASAP7_75t_SL g2377 ( 
.A(n_2331),
.Y(n_2377)
);

CKINVDCx20_ASAP7_75t_R g2378 ( 
.A(n_2344),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2335),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2349),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2335),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2346),
.B(n_205),
.Y(n_2382)
);

INVx2_ASAP7_75t_SL g2383 ( 
.A(n_2349),
.Y(n_2383)
);

INVxp33_ASAP7_75t_SL g2384 ( 
.A(n_2331),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2335),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2349),
.Y(n_2386)
);

AOI31xp33_ASAP7_75t_L g2387 ( 
.A1(n_2375),
.A2(n_209),
.A3(n_206),
.B(n_207),
.Y(n_2387)
);

OAI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_2382),
.A2(n_2365),
.B1(n_2362),
.B2(n_2367),
.Y(n_2388)
);

OAI21xp33_ASAP7_75t_L g2389 ( 
.A1(n_2352),
.A2(n_2147),
.B(n_2148),
.Y(n_2389)
);

OAI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_2369),
.A2(n_2356),
.B1(n_2381),
.B2(n_2379),
.C(n_2376),
.Y(n_2390)
);

OAI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2355),
.A2(n_2147),
.B(n_2148),
.Y(n_2391)
);

A2O1A1Ixp33_ASAP7_75t_L g2392 ( 
.A1(n_2353),
.A2(n_211),
.B(n_207),
.C(n_209),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_2354),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2378),
.A2(n_2163),
.B1(n_2108),
.B2(n_2000),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2385),
.B(n_212),
.Y(n_2395)
);

AOI32xp33_ASAP7_75t_L g2396 ( 
.A1(n_2380),
.A2(n_2000),
.A3(n_2175),
.B1(n_2163),
.B2(n_2157),
.Y(n_2396)
);

OAI221xp5_ASAP7_75t_L g2397 ( 
.A1(n_2363),
.A2(n_2364),
.B1(n_2359),
.B2(n_2358),
.C(n_2366),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2377),
.A2(n_2163),
.B1(n_2155),
.B2(n_1991),
.Y(n_2398)
);

AOI221xp5_ASAP7_75t_L g2399 ( 
.A1(n_2361),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.C(n_215),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_2351),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2384),
.A2(n_2155),
.B1(n_2157),
.B2(n_1961),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2370),
.Y(n_2402)
);

OAI221xp5_ASAP7_75t_L g2403 ( 
.A1(n_2359),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.C(n_217),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2383),
.Y(n_2404)
);

AOI221xp5_ASAP7_75t_L g2405 ( 
.A1(n_2374),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.C(n_219),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2360),
.Y(n_2406)
);

AO22x1_ASAP7_75t_L g2407 ( 
.A1(n_2386),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_2407)
);

A2O1A1Ixp33_ASAP7_75t_L g2408 ( 
.A1(n_2373),
.A2(n_2372),
.B(n_2371),
.C(n_2357),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2357),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2368),
.A2(n_1972),
.B1(n_1959),
.B2(n_1989),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2375),
.Y(n_2411)
);

OAI21xp33_ASAP7_75t_SL g2412 ( 
.A1(n_2356),
.A2(n_2175),
.B(n_2164),
.Y(n_2412)
);

AOI322xp5_ASAP7_75t_L g2413 ( 
.A1(n_2358),
.A2(n_2128),
.A3(n_2127),
.B1(n_223),
.B2(n_224),
.C1(n_225),
.C2(n_226),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2375),
.Y(n_2414)
);

A2O1A1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2355),
.A2(n_223),
.B(n_220),
.C(n_222),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2358),
.B(n_2127),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2402),
.A2(n_1972),
.B1(n_2164),
.B2(n_2178),
.Y(n_2417)
);

OAI21xp33_ASAP7_75t_SL g2418 ( 
.A1(n_2405),
.A2(n_222),
.B(n_225),
.Y(n_2418)
);

OAI21xp33_ASAP7_75t_SL g2419 ( 
.A1(n_2393),
.A2(n_227),
.B(n_228),
.Y(n_2419)
);

INVxp67_ASAP7_75t_L g2420 ( 
.A(n_2400),
.Y(n_2420)
);

AOI221xp5_ASAP7_75t_L g2421 ( 
.A1(n_2390),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.C(n_230),
.Y(n_2421)
);

NAND4xp75_ASAP7_75t_L g2422 ( 
.A(n_2395),
.B(n_231),
.C(n_229),
.D(n_230),
.Y(n_2422)
);

AOI211xp5_ASAP7_75t_L g2423 ( 
.A1(n_2388),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2423)
);

OAI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2402),
.A2(n_2406),
.B1(n_2404),
.B2(n_2397),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2416),
.B(n_2128),
.Y(n_2425)
);

OAI321xp33_ASAP7_75t_L g2426 ( 
.A1(n_2409),
.A2(n_233),
.A3(n_234),
.B1(n_235),
.B2(n_236),
.C(n_237),
.Y(n_2426)
);

OAI221xp5_ASAP7_75t_L g2427 ( 
.A1(n_2408),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.C(n_238),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2387),
.Y(n_2428)
);

AOI321xp33_ASAP7_75t_L g2429 ( 
.A1(n_2411),
.A2(n_238),
.A3(n_239),
.B1(n_240),
.B2(n_241),
.C(n_242),
.Y(n_2429)
);

NAND5xp2_ASAP7_75t_L g2430 ( 
.A(n_2414),
.B(n_239),
.C(n_240),
.D(n_241),
.E(n_242),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2403),
.Y(n_2431)
);

NOR3xp33_ASAP7_75t_SL g2432 ( 
.A(n_2392),
.B(n_243),
.C(n_244),
.Y(n_2432)
);

INVx1_ASAP7_75t_SL g2433 ( 
.A(n_2407),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2415),
.B(n_243),
.Y(n_2434)
);

AOI311xp33_ASAP7_75t_L g2435 ( 
.A1(n_2399),
.A2(n_244),
.A3(n_245),
.B(n_246),
.C(n_247),
.Y(n_2435)
);

AOI221xp5_ASAP7_75t_L g2436 ( 
.A1(n_2410),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.C(n_248),
.Y(n_2436)
);

NOR3xp33_ASAP7_75t_L g2437 ( 
.A(n_2412),
.B(n_248),
.C(n_249),
.Y(n_2437)
);

O2A1O1Ixp33_ASAP7_75t_L g2438 ( 
.A1(n_2389),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_2438)
);

AOI211xp5_ASAP7_75t_L g2439 ( 
.A1(n_2391),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_2439)
);

AOI322xp5_ASAP7_75t_L g2440 ( 
.A1(n_2401),
.A2(n_253),
.A3(n_254),
.B1(n_255),
.B2(n_256),
.C1(n_257),
.C2(n_258),
.Y(n_2440)
);

OAI211xp5_ASAP7_75t_L g2441 ( 
.A1(n_2396),
.A2(n_253),
.B(n_254),
.C(n_255),
.Y(n_2441)
);

AOI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2398),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.C(n_260),
.Y(n_2442)
);

AOI221xp5_ASAP7_75t_L g2443 ( 
.A1(n_2394),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.C(n_263),
.Y(n_2443)
);

NAND3xp33_ASAP7_75t_SL g2444 ( 
.A(n_2413),
.B(n_261),
.C(n_262),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2400),
.Y(n_2445)
);

O2A1O1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2400),
.A2(n_264),
.B(n_265),
.C(n_266),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_SL g2447 ( 
.A1(n_2390),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C(n_267),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2400),
.Y(n_2448)
);

NOR4xp75_ASAP7_75t_L g2449 ( 
.A(n_2390),
.B(n_268),
.C(n_269),
.D(n_270),
.Y(n_2449)
);

INVx2_ASAP7_75t_SL g2450 ( 
.A(n_2402),
.Y(n_2450)
);

A2O1A1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2393),
.A2(n_269),
.B(n_270),
.C(n_271),
.Y(n_2451)
);

INVx1_ASAP7_75t_SL g2452 ( 
.A(n_2407),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2402),
.B(n_271),
.Y(n_2453)
);

AOI211xp5_ASAP7_75t_L g2454 ( 
.A1(n_2390),
.A2(n_272),
.B(n_273),
.C(n_274),
.Y(n_2454)
);

NAND3xp33_ASAP7_75t_SL g2455 ( 
.A(n_2405),
.B(n_275),
.C(n_276),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2402),
.B(n_275),
.Y(n_2456)
);

OA211x2_ASAP7_75t_L g2457 ( 
.A1(n_2421),
.A2(n_276),
.B(n_277),
.C(n_278),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2453),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2450),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_2459)
);

NAND5xp2_ASAP7_75t_L g2460 ( 
.A(n_2445),
.B(n_280),
.C(n_281),
.D(n_282),
.E(n_283),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2419),
.Y(n_2461)
);

AOI211xp5_ASAP7_75t_L g2462 ( 
.A1(n_2424),
.A2(n_280),
.B(n_281),
.C(n_283),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2456),
.A2(n_284),
.B(n_285),
.Y(n_2463)
);

O2A1O1Ixp33_ASAP7_75t_L g2464 ( 
.A1(n_2420),
.A2(n_284),
.B(n_285),
.C(n_286),
.Y(n_2464)
);

AOI211x1_ASAP7_75t_SL g2465 ( 
.A1(n_2444),
.A2(n_286),
.B(n_287),
.C(n_288),
.Y(n_2465)
);

AOI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2448),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2447),
.B(n_289),
.Y(n_2467)
);

OAI221xp5_ASAP7_75t_L g2468 ( 
.A1(n_2454),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.C(n_294),
.Y(n_2468)
);

AOI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2434),
.A2(n_291),
.B(n_292),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2429),
.B(n_2423),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2451),
.B(n_294),
.Y(n_2471)
);

NAND4xp25_ASAP7_75t_L g2472 ( 
.A(n_2435),
.B(n_295),
.C(n_296),
.D(n_297),
.Y(n_2472)
);

OAI221xp5_ASAP7_75t_L g2473 ( 
.A1(n_2436),
.A2(n_2443),
.B1(n_2442),
.B2(n_2418),
.C(n_2437),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2433),
.A2(n_2452),
.B1(n_2428),
.B2(n_2455),
.Y(n_2474)
);

OAI211xp5_ASAP7_75t_L g2475 ( 
.A1(n_2427),
.A2(n_295),
.B(n_297),
.C(n_298),
.Y(n_2475)
);

NAND2x1p5_ASAP7_75t_L g2476 ( 
.A(n_2431),
.B(n_2449),
.Y(n_2476)
);

O2A1O1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_2446),
.A2(n_298),
.B(n_299),
.C(n_300),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2430),
.Y(n_2478)
);

AOI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2438),
.A2(n_299),
.B(n_301),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2422),
.B(n_302),
.Y(n_2480)
);

OAI211xp5_ASAP7_75t_SL g2481 ( 
.A1(n_2432),
.A2(n_302),
.B(n_303),
.C(n_304),
.Y(n_2481)
);

OAI311xp33_ASAP7_75t_L g2482 ( 
.A1(n_2440),
.A2(n_304),
.A3(n_305),
.B1(n_306),
.C1(n_307),
.Y(n_2482)
);

OAI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2426),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2425),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_2484)
);

NOR3x1_ASAP7_75t_L g2485 ( 
.A(n_2441),
.B(n_311),
.C(n_312),
.Y(n_2485)
);

NOR3xp33_ASAP7_75t_L g2486 ( 
.A(n_2439),
.B(n_312),
.C(n_313),
.Y(n_2486)
);

AO221x1_ASAP7_75t_L g2487 ( 
.A1(n_2417),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.C(n_316),
.Y(n_2487)
);

OAI211xp5_ASAP7_75t_L g2488 ( 
.A1(n_2419),
.A2(n_314),
.B(n_315),
.C(n_317),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2453),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2480),
.Y(n_2490)
);

NOR2x1_ASAP7_75t_L g2491 ( 
.A(n_2461),
.B(n_317),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2485),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2484),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2488),
.Y(n_2494)
);

OAI22xp5_ASAP7_75t_L g2495 ( 
.A1(n_2474),
.A2(n_318),
.B1(n_320),
.B2(n_322),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2478),
.B(n_2109),
.Y(n_2496)
);

INVxp67_ASAP7_75t_SL g2497 ( 
.A(n_2464),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2457),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2476),
.Y(n_2499)
);

AO22x2_ASAP7_75t_L g2500 ( 
.A1(n_2458),
.A2(n_322),
.B1(n_323),
.B2(n_325),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2483),
.B(n_323),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2471),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2487),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2460),
.B(n_325),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2489),
.Y(n_2505)
);

NOR2xp67_ASAP7_75t_L g2506 ( 
.A(n_2472),
.B(n_326),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2477),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2465),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2467),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_2462),
.B(n_326),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2468),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2475),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2459),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2470),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2481),
.A2(n_327),
.B1(n_329),
.B2(n_330),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2486),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2463),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2479),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2466),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2469),
.B(n_327),
.Y(n_2520)
);

AOI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2473),
.A2(n_330),
.B1(n_331),
.B2(n_333),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2482),
.B(n_334),
.Y(n_2522)
);

OR3x1_ASAP7_75t_L g2523 ( 
.A(n_2504),
.B(n_334),
.C(n_335),
.Y(n_2523)
);

XNOR2xp5_ASAP7_75t_L g2524 ( 
.A(n_2514),
.B(n_2499),
.Y(n_2524)
);

NOR2x1p5_ASAP7_75t_L g2525 ( 
.A(n_2522),
.B(n_335),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2491),
.B(n_336),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2498),
.Y(n_2527)
);

NAND4xp75_ASAP7_75t_L g2528 ( 
.A(n_2494),
.B(n_337),
.C(n_338),
.D(n_339),
.Y(n_2528)
);

AND4x1_ASAP7_75t_L g2529 ( 
.A(n_2512),
.B(n_338),
.C(n_340),
.D(n_341),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2495),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2500),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2509),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2515),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2505),
.Y(n_2534)
);

NAND2x1p5_ASAP7_75t_L g2535 ( 
.A(n_2503),
.B(n_340),
.Y(n_2535)
);

NAND4xp25_ASAP7_75t_L g2536 ( 
.A(n_2506),
.B(n_342),
.C(n_343),
.D(n_344),
.Y(n_2536)
);

AOI321xp33_ASAP7_75t_L g2537 ( 
.A1(n_2501),
.A2(n_343),
.A3(n_344),
.B1(n_345),
.B2(n_346),
.C(n_347),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_SL g2538 ( 
.A(n_2492),
.B(n_345),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_R g2539 ( 
.A(n_2508),
.B(n_346),
.Y(n_2539)
);

NOR2x1_ASAP7_75t_L g2540 ( 
.A(n_2518),
.B(n_347),
.Y(n_2540)
);

NOR2x1_ASAP7_75t_L g2541 ( 
.A(n_2517),
.B(n_2507),
.Y(n_2541)
);

NAND3xp33_ASAP7_75t_L g2542 ( 
.A(n_2524),
.B(n_2516),
.C(n_2511),
.Y(n_2542)
);

XNOR2xp5_ASAP7_75t_L g2543 ( 
.A(n_2523),
.B(n_2521),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_R g2544 ( 
.A(n_2532),
.B(n_2519),
.Y(n_2544)
);

NAND2xp33_ASAP7_75t_SL g2545 ( 
.A(n_2539),
.B(n_2520),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2535),
.B(n_2496),
.Y(n_2546)
);

XNOR2x1_ASAP7_75t_L g2547 ( 
.A(n_2525),
.B(n_2513),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_SL g2548 ( 
.A(n_2526),
.B(n_2493),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2537),
.B(n_2490),
.Y(n_2549)
);

NAND2xp33_ASAP7_75t_SL g2550 ( 
.A(n_2534),
.B(n_2510),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_R g2551 ( 
.A(n_2534),
.B(n_2502),
.Y(n_2551)
);

NAND3xp33_ASAP7_75t_L g2552 ( 
.A(n_2527),
.B(n_2497),
.C(n_2500),
.Y(n_2552)
);

NAND2xp33_ASAP7_75t_SL g2553 ( 
.A(n_2531),
.B(n_2533),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_SL g2554 ( 
.A(n_2530),
.B(n_348),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2543),
.B(n_2540),
.Y(n_2555)
);

NAND4xp25_ASAP7_75t_L g2556 ( 
.A(n_2542),
.B(n_2541),
.C(n_2536),
.D(n_2538),
.Y(n_2556)
);

NOR2x1_ASAP7_75t_L g2557 ( 
.A(n_2552),
.B(n_2528),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2554),
.Y(n_2558)
);

HB1xp67_ASAP7_75t_L g2559 ( 
.A(n_2544),
.Y(n_2559)
);

NOR3xp33_ASAP7_75t_L g2560 ( 
.A(n_2553),
.B(n_2529),
.C(n_348),
.Y(n_2560)
);

NOR3xp33_ASAP7_75t_SL g2561 ( 
.A(n_2550),
.B(n_464),
.C(n_465),
.Y(n_2561)
);

NOR3xp33_ASAP7_75t_L g2562 ( 
.A(n_2549),
.B(n_466),
.C(n_468),
.Y(n_2562)
);

OR5x1_ASAP7_75t_L g2563 ( 
.A(n_2547),
.B(n_469),
.C(n_470),
.D(n_471),
.E(n_472),
.Y(n_2563)
);

NOR3xp33_ASAP7_75t_L g2564 ( 
.A(n_2545),
.B(n_473),
.C(n_474),
.Y(n_2564)
);

INVx2_ASAP7_75t_SL g2565 ( 
.A(n_2557),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2563),
.Y(n_2566)
);

XNOR2xp5_ASAP7_75t_L g2567 ( 
.A(n_2559),
.B(n_2546),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2555),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2560),
.Y(n_2569)
);

AO21x2_ASAP7_75t_L g2570 ( 
.A1(n_2567),
.A2(n_2551),
.B(n_2558),
.Y(n_2570)
);

HB1xp67_ASAP7_75t_L g2571 ( 
.A(n_2566),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2565),
.A2(n_2568),
.B1(n_2561),
.B2(n_2569),
.Y(n_2572)
);

OAI21x1_ASAP7_75t_L g2573 ( 
.A1(n_2567),
.A2(n_2556),
.B(n_2548),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2571),
.A2(n_2562),
.B1(n_2564),
.B2(n_482),
.Y(n_2574)
);

OAI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2572),
.A2(n_478),
.B1(n_480),
.B2(n_483),
.Y(n_2575)
);

OA22x2_ASAP7_75t_L g2576 ( 
.A1(n_2573),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_2576)
);

AOI211xp5_ASAP7_75t_L g2577 ( 
.A1(n_2574),
.A2(n_2575),
.B(n_2570),
.C(n_2576),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2574),
.Y(n_2578)
);

OAI22xp5_ASAP7_75t_SL g2579 ( 
.A1(n_2574),
.A2(n_488),
.B1(n_489),
.B2(n_491),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2578),
.A2(n_2579),
.B1(n_2577),
.B2(n_498),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2578),
.A2(n_496),
.B1(n_497),
.B2(n_499),
.Y(n_2581)
);

AOI31xp33_ASAP7_75t_L g2582 ( 
.A1(n_2577),
.A2(n_500),
.A3(n_501),
.B(n_503),
.Y(n_2582)
);

A2O1A1Ixp33_ASAP7_75t_L g2583 ( 
.A1(n_2580),
.A2(n_504),
.B(n_507),
.C(n_508),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2582),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2584),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2583),
.A2(n_2581),
.B(n_512),
.Y(n_2586)
);

OAI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2585),
.A2(n_511),
.B1(n_513),
.B2(n_514),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2587),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2588),
.Y(n_2589)
);

OAI221xp5_ASAP7_75t_R g2590 ( 
.A1(n_2589),
.A2(n_2586),
.B1(n_517),
.B2(n_519),
.C(n_520),
.Y(n_2590)
);

AOI21xp33_ASAP7_75t_SL g2591 ( 
.A1(n_2590),
.A2(n_515),
.B(n_523),
.Y(n_2591)
);

AOI211xp5_ASAP7_75t_L g2592 ( 
.A1(n_2591),
.A2(n_524),
.B(n_525),
.C(n_526),
.Y(n_2592)
);


endmodule