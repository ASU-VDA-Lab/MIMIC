module fake_jpeg_15912_n_201 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_36),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_56),
.B1(n_32),
.B2(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_3),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_3),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_23),
.B(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_25),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_19),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_61),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_88),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_47),
.B1(n_44),
.B2(n_42),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_81),
.B1(n_78),
.B2(n_69),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_29),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_79),
.B(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_80),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_22),
.B1(n_21),
.B2(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_16),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_14),
.CI(n_17),
.CON(n_91),
.SN(n_91)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_93),
.B(n_103),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_100),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_12),
.B(n_13),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_115),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_14),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_49),
.B1(n_5),
.B2(n_13),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_104),
.B(n_106),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_48),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_14),
.B1(n_70),
.B2(n_66),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_73),
.B(n_79),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_74),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_63),
.B(n_71),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_113),
.B(n_95),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_77),
.C(n_63),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_116),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_84),
.B(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_60),
.B1(n_75),
.B2(n_87),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_62),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_103),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_126),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_131),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_137),
.B(n_105),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_135),
.Y(n_146)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_101),
.B1(n_94),
.B2(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_118),
.B1(n_124),
.B2(n_140),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_92),
.B1(n_100),
.B2(n_115),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_147),
.B1(n_157),
.B2(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_91),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_154),
.C(n_155),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_97),
.B1(n_105),
.B2(n_128),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_153),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_133),
.C(n_125),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_133),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_129),
.B1(n_121),
.B2(n_120),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_142),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_137),
.B1(n_123),
.B2(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_122),
.B(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_154),
.C(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_172),
.C(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_145),
.C(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_173),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_182),
.C(n_171),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_144),
.B1(n_148),
.B2(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_146),
.B1(n_165),
.B2(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_165),
.C(n_160),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_146),
.B1(n_167),
.B2(n_170),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AOI21x1_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_162),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_176),
.B1(n_174),
.B2(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_161),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_187),
.B(n_189),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_193),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_177),
.B1(n_179),
.B2(n_190),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_192),
.C(n_191),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_196),
.B(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_197),
.Y(n_201)
);


endmodule