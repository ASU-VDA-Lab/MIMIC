module fake_jpeg_6699_n_39 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_16),
.B1(n_8),
.B2(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI21x1_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_4),
.B(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_0),
.B(n_13),
.C(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_0),
.B1(n_20),
.B2(n_19),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_31),
.B(n_32),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);


endmodule