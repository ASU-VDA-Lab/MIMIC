module fake_jpeg_11278_n_455 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_57),
.B(n_62),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_59),
.B(n_44),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_14),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_64),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_67),
.B(n_78),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_74),
.Y(n_127)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_13),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_0),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_91),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_98),
.Y(n_144)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_96),
.B(n_32),
.Y(n_166)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_19),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_105),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_1),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_110),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_5),
.B(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_39),
.B1(n_29),
.B2(n_42),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_113),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_40),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_19),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_20),
.B(n_5),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_55),
.B1(n_27),
.B2(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_119),
.A2(n_122),
.B1(n_177),
.B2(n_112),
.Y(n_200)
);

AND2x4_ASAP7_75t_SL g120 ( 
.A(n_77),
.B(n_40),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_120),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_55),
.B1(n_27),
.B2(n_49),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_121),
.A2(n_159),
.B1(n_180),
.B2(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_55),
.B1(n_27),
.B2(n_21),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_51),
.B1(n_35),
.B2(n_21),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_124),
.A2(n_133),
.B1(n_136),
.B2(n_140),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_60),
.A2(n_50),
.B1(n_46),
.B2(n_56),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g230 ( 
.A1(n_126),
.A2(n_131),
.B1(n_161),
.B2(n_167),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_50),
.B1(n_46),
.B2(n_56),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_50),
.B1(n_42),
.B2(n_34),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_135),
.A2(n_162),
.B1(n_184),
.B2(n_102),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_59),
.A2(n_42),
.B1(n_39),
.B2(n_29),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_42),
.B1(n_39),
.B2(n_29),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_47),
.CON(n_142),
.SN(n_142)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_51),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_145),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_75),
.B(n_76),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_69),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_32),
.B1(n_48),
.B2(n_45),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_71),
.A2(n_39),
.B1(n_29),
.B2(n_47),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_166),
.B(n_168),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_20),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_52),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_172),
.B(n_173),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_65),
.B(n_37),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_103),
.A2(n_37),
.B1(n_48),
.B2(n_45),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_147),
.B1(n_176),
.B2(n_148),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_73),
.A2(n_52),
.B1(n_47),
.B2(n_9),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_149),
.B(n_137),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_65),
.B(n_7),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_181),
.B(n_185),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_80),
.A2(n_11),
.B1(n_12),
.B2(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_90),
.B(n_11),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_186),
.B(n_242),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_90),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_187),
.B(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_201),
.Y(n_250)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_121),
.A2(n_97),
.B1(n_72),
.B2(n_81),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_191),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_12),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_192),
.B(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_12),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g285 ( 
.A(n_195),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_196),
.A2(n_221),
.B1(n_234),
.B2(n_226),
.Y(n_291)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_104),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_82),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_199),
.B(n_217),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

BUFx16f_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_230),
.B1(n_191),
.B2(n_209),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_135),
.A2(n_83),
.B1(n_100),
.B2(n_106),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_206),
.A2(n_211),
.B(n_214),
.Y(n_273)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_120),
.A2(n_107),
.A3(n_104),
.B1(n_92),
.B2(n_12),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_208),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_138),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_222),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_142),
.A2(n_146),
.B(n_120),
.C(n_145),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_141),
.B(n_139),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_238),
.C(n_215),
.Y(n_252)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_163),
.B1(n_158),
.B2(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

CKINVDCx9p33_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_117),
.B(n_134),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_132),
.B1(n_126),
.B2(n_131),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_183),
.B1(n_178),
.B2(n_118),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_132),
.A2(n_137),
.B1(n_156),
.B2(n_160),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_165),
.B1(n_167),
.B2(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_224),
.B(n_237),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_240),
.Y(n_269)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_183),
.A2(n_178),
.B1(n_160),
.B2(n_164),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_236),
.B1(n_206),
.B2(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_141),
.A2(n_169),
.B1(n_130),
.B2(n_143),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_165),
.A2(n_170),
.B1(n_182),
.B2(n_143),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_128),
.B(n_170),
.Y(n_238)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_155),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_243),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_155),
.B(n_169),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_151),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_245),
.Y(n_277)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_116),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_216),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_260),
.B1(n_282),
.B2(n_236),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_192),
.C(n_194),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_254),
.B(n_266),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_291),
.B1(n_236),
.B2(n_218),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_209),
.B1(n_230),
.B2(n_191),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_211),
.C(n_193),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_207),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_267),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_234),
.C(n_196),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_281),
.B(n_284),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_230),
.A2(n_191),
.B1(n_236),
.B2(n_240),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_202),
.B(n_222),
.C(n_208),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_230),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_188),
.B(n_243),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_265),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_231),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_245),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_317),
.B1(n_280),
.B2(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_227),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_296),
.B(n_301),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_229),
.B(n_195),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_303),
.B(n_305),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_298),
.A2(n_307),
.B1(n_308),
.B2(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_235),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

AOI22x1_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_267),
.B1(n_284),
.B2(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_312),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_195),
.B(n_201),
.C(n_213),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_255),
.A2(n_228),
.B1(n_203),
.B2(n_241),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_255),
.A2(n_244),
.B1(n_197),
.B2(n_204),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_201),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_309),
.B(n_310),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_263),
.B(n_195),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_315),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_273),
.A2(n_258),
.B1(n_281),
.B2(n_252),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_277),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_273),
.B(n_266),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_319),
.Y(n_346)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_247),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_259),
.B(n_286),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_323),
.B(n_251),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_250),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_261),
.A2(n_269),
.B(n_278),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_327),
.B(n_262),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_262),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_328),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_254),
.B(n_265),
.C(n_271),
.D(n_261),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_329),
.B(n_311),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_330),
.B(n_351),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_336),
.A2(n_341),
.B1(n_307),
.B2(n_308),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_314),
.A2(n_251),
.B1(n_264),
.B2(n_275),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_345),
.B1(n_352),
.B2(n_328),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_317),
.B1(n_306),
.B2(n_303),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_343),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_298),
.A2(n_275),
.B1(n_288),
.B2(n_278),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g347 ( 
.A1(n_294),
.A2(n_288),
.A3(n_275),
.B1(n_285),
.B2(n_256),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_338),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_320),
.A2(n_276),
.B(n_285),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_349),
.A2(n_326),
.B(n_316),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_276),
.C(n_256),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_305),
.C(n_325),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_285),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_303),
.A2(n_293),
.B1(n_317),
.B2(n_297),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_326),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_355),
.A2(n_334),
.B1(n_348),
.B2(n_332),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_372),
.B(n_329),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_346),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_358),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_361),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_334),
.A2(n_313),
.B1(n_324),
.B2(n_315),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_342),
.B(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_364),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_370),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_327),
.Y(n_366)
);

XOR2x1_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_375),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_299),
.B1(n_300),
.B2(n_305),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_374),
.B1(n_377),
.B2(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_369),
.Y(n_381)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_371),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_337),
.B(n_312),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_376),
.C(n_350),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_305),
.B1(n_318),
.B2(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_337),
.B(n_302),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_330),
.C(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_305),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_342),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_391),
.C(n_392),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_373),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_362),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_347),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_373),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_331),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_349),
.C(n_339),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_331),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_393),
.A2(n_363),
.B1(n_367),
.B2(n_345),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_329),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_370),
.C(n_360),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_396),
.A2(n_364),
.B1(n_368),
.B2(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_404),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_401),
.A2(n_408),
.B1(n_379),
.B2(n_389),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g405 ( 
.A1(n_395),
.A2(n_358),
.A3(n_362),
.B1(n_332),
.B2(n_365),
.C1(n_372),
.C2(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_405),
.B(n_406),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_367),
.C(n_366),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_340),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_339),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_392),
.B(n_340),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_381),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_411),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_414),
.B(n_422),
.Y(n_431)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_411),
.Y(n_415)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_415),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_406),
.Y(n_417)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_408),
.A2(n_389),
.B1(n_380),
.B2(n_381),
.Y(n_422)
);

BUFx4f_ASAP7_75t_SL g424 ( 
.A(n_421),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_413),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_348),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_426),
.B(n_430),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_407),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_418),
.C(n_407),
.Y(n_436)
);

OAI211xp5_ASAP7_75t_L g430 ( 
.A1(n_423),
.A2(n_410),
.B(n_388),
.C(n_387),
.Y(n_430)
);

OAI21xp33_ASAP7_75t_L g432 ( 
.A1(n_412),
.A2(n_399),
.B(n_402),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_382),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_428),
.A2(n_412),
.B(n_419),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_433),
.A2(n_434),
.B(n_439),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_420),
.B(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_437),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_397),
.C(n_390),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_413),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_396),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_SL g446 ( 
.A(n_438),
.B(n_383),
.C(n_359),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_391),
.B1(n_420),
.B2(n_388),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_440),
.A2(n_431),
.B(n_424),
.Y(n_444)
);

OAI21x1_ASAP7_75t_SL g447 ( 
.A1(n_444),
.A2(n_445),
.B(n_446),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_414),
.B(n_393),
.Y(n_445)
);

AOI21xp33_ASAP7_75t_L g452 ( 
.A1(n_448),
.A2(n_450),
.B(n_394),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_443),
.A2(n_383),
.B1(n_369),
.B2(n_371),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

AOI21x1_ASAP7_75t_SL g450 ( 
.A1(n_442),
.A2(n_386),
.B(n_361),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_SL g453 ( 
.A1(n_452),
.A2(n_447),
.B(n_450),
.C(n_445),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_451),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_353),
.Y(n_455)
);


endmodule