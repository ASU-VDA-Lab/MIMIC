module fake_netlist_5_389_n_70 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_70);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_70;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_46;
wire n_28;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_38;
wire n_61;
wire n_68;
wire n_32;
wire n_41;
wire n_35;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_20;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_39;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_2),
.B(n_3),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_0),
.Y(n_22)
);

AND2x6_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_5),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp67_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_30),
.Y(n_42)
);

OAI21x1_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_21),
.B(n_31),
.Y(n_43)
);

AO31x2_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_36),
.A3(n_41),
.B(n_37),
.Y(n_44)
);

OA21x2_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_24),
.B(n_25),
.Y(n_45)
);

AO31x2_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_23),
.A3(n_24),
.B(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_47),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_46),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_51),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_57),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_20),
.C(n_43),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_58),
.B(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_24),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_R g67 ( 
.A(n_66),
.B(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_25),
.B(n_28),
.Y(n_69)
);

NOR2x1_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_28),
.Y(n_70)
);


endmodule