module fake_jpeg_29551_n_146 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_34),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_42),
.B1(n_14),
.B2(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_22),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_23),
.B(n_26),
.C(n_15),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_29),
.A2(n_28),
.B1(n_17),
.B2(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_38),
.B1(n_14),
.B2(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_18),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_24),
.B1(n_15),
.B2(n_20),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_73),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_45),
.B1(n_55),
.B2(n_63),
.Y(n_91)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_70),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_51),
.B1(n_47),
.B2(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_17),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_54),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_37),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_72),
.C(n_85),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_40),
.B1(n_27),
.B2(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_51),
.B1(n_47),
.B2(n_54),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_100),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_78),
.B(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_83),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_55),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_77),
.C(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2x1p5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_78),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_96),
.A3(n_102),
.B1(n_95),
.B2(n_74),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_75),
.B(n_99),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_93),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_84),
.B(n_85),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_114),
.B(n_97),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_71),
.B(n_82),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_90),
.B1(n_89),
.B2(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_113),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_109),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_113),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_127),
.B(n_129),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_119),
.B(n_121),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_122),
.A3(n_116),
.B1(n_120),
.B2(n_87),
.C1(n_70),
.C2(n_86),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_104),
.C(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_94),
.C(n_3),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_128),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_120),
.B1(n_73),
.B2(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_1),
.C(n_4),
.D(n_5),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_137),
.B1(n_134),
.B2(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

OAI221xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_6),
.Y(n_143)
);

AOI21x1_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_141),
.B(n_6),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_7),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_145),
.Y(n_146)
);


endmodule