module fake_jpeg_16849_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_32),
.B1(n_33),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_56),
.B1(n_61),
.B2(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_17),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_33),
.B1(n_18),
.B2(n_21),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_21),
.B1(n_18),
.B2(n_47),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_98),
.B1(n_44),
.B2(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_69),
.A2(n_72),
.B1(n_100),
.B2(n_27),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_44),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_20),
.B1(n_22),
.B2(n_39),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_24),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_16),
.B(n_37),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_22),
.B(n_27),
.Y(n_114)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_37),
.B1(n_61),
.B2(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_28),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_23),
.B1(n_16),
.B2(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_24),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_109),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_87),
.B1(n_91),
.B2(n_80),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_126),
.B1(n_74),
.B2(n_98),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_39),
.C(n_30),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_123),
.C(n_93),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_0),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_20),
.CI(n_22),
.CON(n_119),
.SN(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_96),
.B(n_85),
.C(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_30),
.C(n_25),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_153),
.B1(n_25),
.B2(n_29),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_84),
.B1(n_85),
.B2(n_83),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_143),
.B1(n_151),
.B2(n_121),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_141),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_122),
.B(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_95),
.B1(n_86),
.B2(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_73),
.C(n_68),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_117),
.C(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_88),
.B1(n_71),
.B2(n_76),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_68),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_164),
.C(n_165),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_111),
.B1(n_119),
.B2(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_158),
.B1(n_180),
.B2(n_130),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_107),
.B1(n_106),
.B2(n_121),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_113),
.B(n_107),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_160),
.C(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_106),
.C(n_108),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_108),
.C(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_112),
.C(n_127),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_102),
.C(n_4),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_115),
.B1(n_97),
.B2(n_78),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_172),
.B(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_128),
.B(n_115),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_25),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_149),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_20),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_30),
.B(n_25),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_177),
.B(n_168),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_151),
.B(n_153),
.C(n_147),
.D(n_138),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_197),
.B1(n_199),
.B2(n_158),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_200),
.C(n_201),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_171),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_198),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_140),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_202),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_136),
.B1(n_29),
.B2(n_132),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_132),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_29),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_3),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_218),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.C(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_166),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_190),
.B1(n_203),
.B2(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_165),
.C(n_175),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_170),
.B(n_175),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_193),
.B(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_170),
.C(n_167),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_167),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_193),
.C(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_174),
.B1(n_159),
.B2(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_210),
.B1(n_191),
.B2(n_157),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_226),
.B1(n_236),
.B2(n_208),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_187),
.B1(n_196),
.B2(n_203),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_189),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_179),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_159),
.B1(n_183),
.B2(n_157),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_241),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_212),
.C(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_220),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_247),
.B(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_208),
.C(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_246),
.Y(n_254)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_240),
.B(n_230),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_229),
.B(n_234),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_256),
.B(n_257),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_224),
.B1(n_236),
.B2(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_189),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_3),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_244),
.C(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.C(n_261),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_242),
.C(n_238),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_7),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_253),
.C(n_11),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_10),
.C(n_12),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_264),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_269),
.C(n_14),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_15),
.Y(n_274)
);


endmodule