module fake_jpeg_1805_n_536 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_536);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_32),
.Y(n_52)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_58),
.Y(n_140)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_63),
.Y(n_119)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_77),
.Y(n_128)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_35),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_8),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_36),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_36),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_99),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_51),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_35),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_111),
.B(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_113),
.B(n_20),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_123),
.B(n_144),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_142),
.Y(n_170)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_24),
.CON(n_133),
.SN(n_133)
);

OR2x2_ASAP7_75t_SL g189 ( 
.A(n_133),
.B(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_84),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_23),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_155),
.Y(n_192)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_46),
.Y(n_155)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_R g159 ( 
.A(n_62),
.Y(n_159)
);

CKINVDCx9p33_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_73),
.B(n_35),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_165),
.A2(n_0),
.B(n_1),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_46),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_49),
.B(n_41),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_67),
.B(n_23),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_53),
.B1(n_59),
.B2(n_57),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_171),
.A2(n_173),
.B1(n_164),
.B2(n_150),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_40),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_172),
.B(n_178),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_66),
.B1(n_77),
.B2(n_79),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_100),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_93),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_182),
.B(n_183),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_91),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_124),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_187),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_195),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_199),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_144),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_200),
.B(n_208),
.Y(n_279)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_120),
.A2(n_50),
.B1(n_41),
.B2(n_49),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_210),
.B1(n_223),
.B2(n_224),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_221),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_76),
.Y(n_208)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_87),
.B1(n_50),
.B2(n_82),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_216),
.A2(n_115),
.B1(n_150),
.B2(n_139),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_225),
.Y(n_248)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_136),
.B(n_89),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_160),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_228),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_109),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_134),
.A2(n_27),
.B1(n_22),
.B2(n_86),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_106),
.B(n_10),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_107),
.A2(n_85),
.B1(n_1),
.B2(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_156),
.B1(n_130),
.B2(n_164),
.Y(n_254)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_108),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_185),
.B1(n_124),
.B2(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_112),
.B(n_11),
.Y(n_230)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_116),
.C(n_165),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_207),
.C(n_202),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_110),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_264),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_254),
.A2(n_273),
.B1(n_196),
.B2(n_191),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_256),
.A2(n_210),
.B1(n_4),
.B2(n_5),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_192),
.B(n_140),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_133),
.B(n_159),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_265),
.A2(n_282),
.B(n_235),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_138),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_270),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_184),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_222),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_216),
.B1(n_201),
.B2(n_179),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_190),
.A2(n_130),
.B1(n_148),
.B2(n_161),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_170),
.B(n_118),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_186),
.B(n_168),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_194),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_187),
.B(n_124),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_189),
.B(n_0),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_0),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_108),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_220),
.Y(n_318)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

XOR2x2_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_226),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_258),
.Y(n_339)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_248),
.C(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_296),
.C(n_315),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_290),
.A2(n_305),
.B1(n_321),
.B2(n_324),
.Y(n_349)
);

AO22x1_ASAP7_75t_SL g291 ( 
.A1(n_254),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_300),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_292),
.B(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

CKINVDCx12_ASAP7_75t_R g295 ( 
.A(n_283),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_308),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_297),
.B(n_311),
.Y(n_338)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_298),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_256),
.A2(n_197),
.B1(n_206),
.B2(n_177),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_299),
.A2(n_329),
.B1(n_269),
.B2(n_260),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_176),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_303),
.A2(n_276),
.B(n_244),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_175),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_306),
.Y(n_365)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_236),
.Y(n_308)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

OR2x4_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_231),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_326),
.Y(n_347)
);

OAI221xp5_ASAP7_75t_L g311 ( 
.A1(n_232),
.A2(n_175),
.B1(n_205),
.B2(n_162),
.C(n_209),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_196),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_271),
.B(n_16),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_314),
.B(n_317),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_209),
.C(n_227),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_239),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_249),
.B(n_218),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_319),
.B(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_234),
.B(n_13),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_233),
.B(n_1),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_331),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_273),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_283),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_233),
.B(n_17),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_237),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_233),
.B(n_14),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_262),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_250),
.B(n_4),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_286),
.A2(n_270),
.B1(n_250),
.B2(n_255),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_334),
.A2(n_346),
.B1(n_356),
.B2(n_358),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_339),
.B(n_362),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_331),
.Y(n_341)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_305),
.A2(n_255),
.B1(n_266),
.B2(n_258),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_234),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_354),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_314),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_310),
.A2(n_267),
.B(n_261),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_364),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_257),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_307),
.Y(n_355)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_327),
.A2(n_257),
.B1(n_245),
.B2(n_261),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_262),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_357),
.B(n_303),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_323),
.A2(n_245),
.B1(n_269),
.B2(n_247),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_243),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_267),
.C(n_260),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_309),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_368),
.B(n_308),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_243),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_302),
.B(n_300),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_328),
.B(n_304),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_372),
.A2(n_379),
.B(n_385),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_316),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_374),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_394),
.C(n_402),
.Y(n_418)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_380),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_335),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_387),
.Y(n_430)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_332),
.A2(n_330),
.B1(n_324),
.B2(n_291),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_384),
.A2(n_397),
.B1(n_334),
.B2(n_344),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_328),
.B(n_370),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_348),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_393),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_396),
.Y(n_410)
);

BUFx12_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_392),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_361),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_306),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_332),
.A2(n_291),
.B1(n_299),
.B2(n_301),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_343),
.Y(n_416)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_400),
.Y(n_412)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_312),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_404),
.Y(n_415)
);

CKINVDCx12_ASAP7_75t_R g402 ( 
.A(n_333),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_338),
.A2(n_329),
.B1(n_297),
.B2(n_326),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_403),
.A2(n_360),
.B(n_340),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_381),
.B(n_343),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_385),
.A2(n_372),
.B(n_375),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_420),
.B(n_433),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_368),
.Y(n_419)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_421),
.A2(n_425),
.B1(n_433),
.B2(n_398),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_388),
.A2(n_364),
.B1(n_350),
.B2(n_339),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_421),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_388),
.A2(n_349),
.B1(n_342),
.B2(n_355),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_403),
.B1(n_390),
.B2(n_386),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_397),
.A2(n_346),
.B1(n_342),
.B2(n_365),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_371),
.Y(n_427)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_381),
.B(n_360),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_429),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_371),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_431),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_340),
.C(n_344),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_320),
.C(n_313),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_375),
.A2(n_365),
.B1(n_353),
.B2(n_367),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_435),
.A2(n_390),
.B(n_400),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_377),
.B(n_353),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_298),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_438),
.A2(n_434),
.B1(n_428),
.B2(n_407),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_426),
.B(n_394),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_440),
.B(n_430),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_441),
.A2(n_448),
.B(n_431),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_405),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_447),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_443),
.A2(n_422),
.B1(n_413),
.B2(n_427),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_410),
.B(n_423),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_446),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_SL g445 ( 
.A(n_418),
.B(n_375),
.C(n_384),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_461),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_379),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_378),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_459),
.B1(n_419),
.B2(n_422),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_383),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_456),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_414),
.A2(n_380),
.B1(n_404),
.B2(n_399),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_457),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_429),
.B(n_358),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_420),
.B(n_292),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_460),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_416),
.A2(n_389),
.B1(n_406),
.B2(n_363),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_363),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_408),
.C(n_417),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_462),
.B(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_465),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_408),
.C(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_469),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_441),
.A2(n_411),
.B(n_415),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_470),
.B(n_478),
.Y(n_484)
);

AO21x1_ASAP7_75t_L g488 ( 
.A1(n_473),
.A2(n_480),
.B(n_459),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_476),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_415),
.C(n_411),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_446),
.C(n_460),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_412),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_434),
.B1(n_428),
.B2(n_407),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_479),
.A2(n_449),
.B1(n_456),
.B2(n_406),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_452),
.B(n_276),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_392),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_466),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_488),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_473),
.A2(n_453),
.B(n_451),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_487),
.B(n_490),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_462),
.C(n_468),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_491),
.B(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_492),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_458),
.C(n_392),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_392),
.C(n_278),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_497),
.C(n_481),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_278),
.C(n_244),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_508),
.Y(n_516)
);

AOI21xp33_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_471),
.B(n_479),
.Y(n_501)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_471),
.B(n_475),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_503),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_476),
.C(n_467),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_287),
.Y(n_504)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_504),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_506),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_472),
.B(n_238),
.Y(n_507)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_472),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_247),
.C(n_275),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_496),
.C(n_497),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_493),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_519),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_503),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_516),
.C(n_505),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_523),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_498),
.B1(n_511),
.B2(n_487),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_514),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_525),
.C(n_516),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_500),
.Y(n_525)
);

AOI322xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_513),
.A3(n_517),
.B1(n_488),
.B2(n_500),
.C1(n_520),
.C2(n_492),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_524),
.B(n_485),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_526),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_529),
.B(n_508),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_532),
.B(n_519),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_533),
.B(n_509),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_495),
.Y(n_535)
);

AOI311xp33_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_7),
.A3(n_274),
.B(n_275),
.C(n_532),
.Y(n_536)
);


endmodule