module fake_jpeg_4096_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_41),
.B1(n_35),
.B2(n_12),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_27),
.B1(n_16),
.B2(n_28),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_50),
.B1(n_61),
.B2(n_15),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_56),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_27),
.B1(n_16),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_16),
.B1(n_20),
.B2(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_53),
.B1(n_64),
.B2(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_20),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_24),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_29),
.B1(n_15),
.B2(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_25),
.B1(n_13),
.B2(n_10),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_15),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_46),
.B(n_47),
.C(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_45),
.B1(n_52),
.B2(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_61),
.B1(n_47),
.B2(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_54),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_60),
.B1(n_49),
.B2(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_92),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_18),
.B(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_69),
.B1(n_83),
.B2(n_82),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_104),
.B(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_97),
.B1(n_82),
.B2(n_79),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_44),
.B1(n_62),
.B2(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_52),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_65),
.B1(n_77),
.B2(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_124),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_75),
.C(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_125),
.C(n_97),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_111),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_67),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_67),
.B1(n_81),
.B2(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_82),
.B1(n_79),
.B2(n_65),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_122),
.B(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_48),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_1),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_99),
.B(n_100),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_59),
.C(n_65),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_133),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_96),
.B(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_136),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_146),
.C(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_142),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_91),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_112),
.B(n_95),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_89),
.B1(n_84),
.B2(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_87),
.B1(n_105),
.B2(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_108),
.B(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_97),
.B(n_89),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_59),
.B(n_25),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_151),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_156),
.B(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_110),
.B(n_123),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_114),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_85),
.C(n_126),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_130),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_85),
.B(n_112),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_86),
.B1(n_87),
.B2(n_94),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_144),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_87),
.B1(n_76),
.B2(n_63),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_107),
.B(n_63),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_63),
.B1(n_72),
.B2(n_107),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_127),
.B1(n_137),
.B2(n_107),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_184),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_148),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_188),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_189),
.B1(n_164),
.B2(n_154),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.C(n_143),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.C(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_138),
.C(n_129),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_138),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_140),
.B1(n_133),
.B2(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_165),
.B1(n_153),
.B2(n_156),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_153),
.B1(n_150),
.B2(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_189),
.B1(n_186),
.B2(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_206),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_157),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_167),
.B(n_152),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_185),
.B(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_72),
.B1(n_25),
.B2(n_18),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.C(n_205),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_171),
.C(n_101),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_101),
.C(n_72),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_101),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_187),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_210),
.B(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_189),
.B1(n_172),
.B2(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_179),
.B(n_186),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_213),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_187),
.C(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_194),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_18),
.B(n_8),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_173),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_205),
.C(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_228),
.C(n_25),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_226),
.B(n_227),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_203),
.B(n_200),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_191),
.C(n_204),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_221),
.A2(n_215),
.B1(n_209),
.B2(n_217),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_211),
.B1(n_219),
.B2(n_213),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_13),
.B(n_12),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_13),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_11),
.B(n_9),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_1),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_224),
.C(n_220),
.Y(n_239)
);

OAI21x1_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_242),
.B(n_2),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_223),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_229),
.C(n_11),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_232),
.A3(n_231),
.B1(n_11),
.B2(n_9),
.C1(n_8),
.C2(n_6),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_240),
.B1(n_6),
.B2(n_7),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_249),
.B(n_6),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_248),
.B(n_7),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_7),
.Y(n_252)
);


endmodule