module fake_jpeg_7560_n_200 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_16),
.B1(n_34),
.B2(n_32),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_34),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_26),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_51),
.B1(n_14),
.B2(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_26),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

OA21x2_ASAP7_75t_R g62 ( 
.A1(n_41),
.A2(n_19),
.B(n_20),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_48),
.B1(n_36),
.B2(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_24),
.B1(n_14),
.B2(n_22),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_42),
.B1(n_43),
.B2(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_84),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_59),
.B1(n_67),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_67),
.B1(n_53),
.B2(n_36),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_68),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_57),
.B(n_56),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_15),
.B(n_22),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_90),
.B1(n_102),
.B2(n_67),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_62),
.B(n_65),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_91),
.B(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_63),
.B1(n_36),
.B2(n_68),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_70),
.B1(n_40),
.B2(n_39),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_60),
.B(n_27),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_75),
.C(n_72),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_117),
.C(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_114),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_77),
.B(n_75),
.C(n_78),
.D(n_76),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_74),
.A3(n_72),
.B1(n_69),
.B2(n_82),
.C1(n_27),
.C2(n_17),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_74),
.C(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_40),
.B1(n_39),
.B2(n_47),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_40),
.B1(n_39),
.B2(n_32),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_23),
.B(n_22),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_13),
.B(n_21),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_130),
.C(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_21),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_0),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_133),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_30),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_113),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_146),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_110),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_107),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_114),
.CI(n_109),
.CON(n_145),
.SN(n_145)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_2),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_66),
.B1(n_52),
.B2(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_131),
.B1(n_120),
.B2(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_154),
.B1(n_35),
.B2(n_30),
.Y(n_166)
);

OAI321xp33_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_125),
.A3(n_52),
.B1(n_20),
.B2(n_80),
.C(n_5),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_3),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_1),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_141),
.C(n_139),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_156),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_27),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_35),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_160),
.B(n_2),
.Y(n_165)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_138),
.C(n_35),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_169),
.C(n_171),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_168),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_150),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_3),
.C(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_4),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_3),
.C(n_4),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_153),
.B(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_177),
.Y(n_183)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_7),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_158),
.B1(n_7),
.B2(n_8),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_5),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_178),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_184),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_175),
.B(n_174),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_186),
.C1(n_188),
.C2(n_163),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_181),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_9),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_193),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_194),
.C(n_195),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_196),
.B(n_191),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);


endmodule