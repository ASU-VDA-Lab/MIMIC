module fake_jpeg_11906_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_46),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_20),
.Y(n_80)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_16),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_68),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_76),
.B(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_20),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_37),
.B1(n_32),
.B2(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_108),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_34),
.B1(n_28),
.B2(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_26),
.B1(n_22),
.B2(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_57),
.B1(n_53),
.B2(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_103),
.B1(n_101),
.B2(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_2),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_99),
.B1(n_81),
.B2(n_100),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_64),
.C(n_48),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_79),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_116),
.B1(n_84),
.B2(n_128),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_43),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_51),
.B1(n_58),
.B2(n_53),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_130),
.B1(n_113),
.B2(n_138),
.Y(n_161)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_4),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_72),
.A2(n_58),
.B1(n_57),
.B2(n_52),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_138),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_47),
.B1(n_8),
.B2(n_9),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_84),
.B(n_87),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_11),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_11),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_157),
.B1(n_159),
.B2(n_123),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_78),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_84),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_161),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_83),
.B1(n_92),
.B2(n_100),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_83),
.B1(n_92),
.B2(n_87),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_12),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_91),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_127),
.A3(n_140),
.B1(n_129),
.B2(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_178),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_114),
.B(n_111),
.C(n_133),
.D(n_139),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_175),
.B(n_182),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_130),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_174),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_110),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_133),
.B1(n_118),
.B2(n_125),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_150),
.B1(n_146),
.B2(n_158),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_131),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_122),
.B1(n_123),
.B2(n_91),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_149),
.B1(n_158),
.B2(n_153),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_197),
.B1(n_171),
.B2(n_148),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_165),
.B(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_144),
.B1(n_160),
.B2(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_177),
.C(n_179),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_170),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_144),
.B1(n_146),
.B2(n_160),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_183),
.C(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_143),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_197),
.B1(n_204),
.B2(n_208),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_176),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_208),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_210)
);

OA21x2_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_193),
.B(n_186),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.C(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_215),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_198),
.B1(n_185),
.B2(n_179),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_198),
.B(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_185),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

AND3x1_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_203),
.C(n_192),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_148),
.B(n_188),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_214),
.C(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_226),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_216),
.B1(n_215),
.B2(n_211),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_223),
.Y(n_230)
);

OAI221xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_145),
.B1(n_148),
.B2(n_153),
.C(n_224),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_145),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_231),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_233),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_227),
.Y(n_236)
);


endmodule