module fake_jpeg_27689_n_272 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_39),
.Y(n_77)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_25),
.B1(n_29),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_73),
.B1(n_48),
.B2(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_65),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_35),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_63),
.C(n_75),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_26),
.B1(n_21),
.B2(n_33),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_18),
.B1(n_30),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_30),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_1),
.B(n_2),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_39),
.Y(n_104)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_48),
.B1(n_30),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_80),
.B1(n_90),
.B2(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_48),
.B1(n_47),
.B2(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_97),
.B1(n_104),
.B2(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_23),
.B1(n_47),
.B2(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_47),
.B1(n_37),
.B2(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_54),
.B1(n_62),
.B2(n_67),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_44),
.B1(n_28),
.B2(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_110),
.B1(n_62),
.B2(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_39),
.B1(n_34),
.B2(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_54),
.Y(n_113)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_59),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_69),
.A3(n_71),
.B1(n_77),
.B2(n_52),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_63),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_68),
.B(n_64),
.C(n_59),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_53),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_85),
.B1(n_96),
.B2(n_99),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_70),
.B1(n_34),
.B2(n_28),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_131),
.B1(n_93),
.B2(n_92),
.Y(n_160)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_70),
.B1(n_34),
.B2(n_19),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_19),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_87),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_150),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_116),
.B(n_119),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_145),
.B(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_159),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_95),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_120),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_87),
.B(n_94),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_157),
.Y(n_170)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_165),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_107),
.B1(n_105),
.B2(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_84),
.B1(n_109),
.B2(n_94),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_3),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_115),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_175),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_180),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_114),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_187),
.C(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_145),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_118),
.C(n_136),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_111),
.C(n_133),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_154),
.C(n_153),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_128),
.B(n_121),
.C(n_137),
.D(n_9),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_156),
.B(n_155),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_153),
.B1(n_165),
.B2(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_200),
.B1(n_211),
.B2(n_183),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_172),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_162),
.B1(n_158),
.B2(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_199),
.B1(n_206),
.B2(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_138),
.B1(n_145),
.B2(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_151),
.B1(n_142),
.B2(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_146),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_147),
.B1(n_121),
.B2(n_8),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_147),
.B1(n_7),
.B2(n_8),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_175),
.C(n_187),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_216),
.C(n_224),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_178),
.B(n_188),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_206),
.B(n_211),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_222),
.B(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_189),
.C(n_178),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_226),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_181),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_221),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_174),
.Y(n_221)
);

AOI321xp33_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_171),
.A3(n_170),
.B1(n_177),
.B2(n_172),
.C(n_179),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_179),
.C(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_185),
.C(n_12),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_225),
.B1(n_202),
.B2(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_238),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_239),
.B(n_227),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_205),
.B1(n_198),
.B2(n_193),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_197),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_R g239 ( 
.A(n_224),
.B(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_212),
.C(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_234),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_234),
.B(n_14),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_216),
.B(n_12),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_11),
.C(n_12),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_11),
.CI(n_13),
.CON(n_250),
.SN(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

OAI221xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_230),
.B1(n_231),
.B2(n_235),
.C(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_241),
.C(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_242),
.C(n_257),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_249),
.B(n_247),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_262),
.B(n_250),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_242),
.C(n_256),
.Y(n_264)
);

OAI21x1_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_250),
.B(n_15),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_266),
.B(n_11),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_15),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.C(n_16),
.Y(n_271)
);

OAI311xp33_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_15),
.A3(n_16),
.B1(n_261),
.C1(n_239),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_261),
.Y(n_272)
);


endmodule