module fake_jpeg_31173_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_1),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_18),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_32),
.C(n_15),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_16),
.C(n_20),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_57),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_44),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_33),
.B(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_19),
.Y(n_78)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_78),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_24),
.Y(n_76)
);

AOI31xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_92),
.A3(n_23),
.B(n_71),
.Y(n_116)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_96),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_16),
.B(n_47),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_89),
.B(n_20),
.Y(n_111)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_43),
.B1(n_26),
.B2(n_46),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_69),
.B1(n_38),
.B2(n_72),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_72),
.B1(n_69),
.B2(n_23),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_109),
.B1(n_88),
.B2(n_79),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_89),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_118),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_7),
.C(n_12),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_2),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_123),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_92),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_132),
.C(n_103),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_74),
.C(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_133),
.C(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_76),
.B1(n_85),
.B2(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_128),
.B1(n_136),
.B2(n_110),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_93),
.B(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_96),
.B1(n_73),
.B2(n_53),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_109),
.B1(n_102),
.B2(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_100),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_14),
.C(n_7),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_13),
.C(n_12),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_143),
.Y(n_156)
);

NOR4xp25_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_115),
.C(n_106),
.D(n_13),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_122),
.C(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_113),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_122),
.B(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_154),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_121),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_156),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_144),
.B1(n_132),
.B2(n_136),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_170),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_107),
.C(n_99),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_166),
.B(n_164),
.C(n_160),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_100),
.A3(n_99),
.B1(n_105),
.B2(n_4),
.C1(n_3),
.C2(n_5),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_161),
.B(n_100),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_105),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_175),
.B(n_173),
.C(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B1(n_105),
.B2(n_5),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);


endmodule