module fake_ibex_2080_n_62 (n_21, n_14, n_12, n_13, n_5, n_20, n_2, n_9, n_8, n_7, n_17, n_10, n_24, n_11, n_18, n_3, n_1, n_4, n_16, n_19, n_6, n_0, n_23, n_22, n_15, n_62);

input n_21;
input n_14;
input n_12;
input n_13;
input n_5;
input n_20;
input n_2;
input n_9;
input n_8;
input n_7;
input n_17;
input n_10;
input n_24;
input n_11;
input n_18;
input n_3;
input n_1;
input n_4;
input n_16;
input n_19;
input n_6;
input n_0;
input n_23;
input n_22;
input n_15;

output n_62;



endmodule