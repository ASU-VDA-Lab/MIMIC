module fake_jpeg_5010_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_SL g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

OA22x2_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_11),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_7),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_10),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_9),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_25),
.C(n_29),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_30),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_33),
.Y(n_38)
);


endmodule