module fake_netlist_1_9326_n_667 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_667);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_667;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_SL g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_0), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_82), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_54), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_36), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_86), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_2), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_84), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_19), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_76), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_26), .B(n_61), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_77), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_3), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_27), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_80), .B(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_57), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_53), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_17), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_18), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_0), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_5), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_33), .Y(n_126) );
CKINVDCx14_ASAP7_75t_R g127 ( .A(n_1), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_10), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_12), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
INVxp33_ASAP7_75t_SL g131 ( .A(n_116), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_127), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_106), .B(n_1), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_92), .B(n_2), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_106), .B(n_3), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_119), .B(n_4), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_96), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_102), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_92), .B(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_102), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_108), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_111), .B(n_5), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_108), .B(n_6), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_124), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_109), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_152), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_130), .A2(n_129), .B1(n_121), .B2(n_105), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_138), .B(n_107), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_130), .A2(n_129), .B1(n_112), .B2(n_113), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_132), .B(n_98), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_131), .B(n_107), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_137), .B(n_112), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_132), .B(n_113), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_138), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_152), .B(n_115), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_138), .B(n_115), .Y(n_178) );
INVx5_ASAP7_75t_L g179 ( .A(n_134), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_157), .B(n_120), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_137), .B(n_118), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_157), .B(n_118), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_134), .Y(n_186) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_156), .B(n_101), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_135), .A2(n_123), .B1(n_114), .B2(n_125), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_163), .B(n_153), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_175), .B(n_136), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_158), .B(n_135), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_163), .B(n_153), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_158), .B(n_146), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_163), .B(n_153), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_191), .B(n_146), .Y(n_200) );
INVx5_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_190), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_191), .B(n_148), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_168), .B(n_143), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_181), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_181), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_166), .B(n_148), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_166), .B(n_150), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_168), .A2(n_150), .B(n_144), .C(n_149), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_166), .B(n_143), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_181), .A2(n_154), .B1(n_149), .B2(n_142), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_177), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_190), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_180), .B(n_154), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_176), .B(n_143), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_176), .B(n_154), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_181), .A2(n_144), .B1(n_139), .B2(n_147), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_180), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_168), .B(n_141), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_181), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_180), .B(n_133), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_181), .B(n_136), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_181), .A2(n_155), .B1(n_122), .B2(n_110), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_184), .B(n_133), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_187), .Y(n_230) );
INVxp67_ASAP7_75t_SL g231 ( .A(n_173), .Y(n_231) );
NOR2x1p5_ASAP7_75t_L g232 ( .A(n_187), .B(n_155), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_189), .A2(n_128), .B1(n_151), .B2(n_145), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_164), .A2(n_123), .B1(n_89), .B2(n_104), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_190), .B(n_151), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_205), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_194), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_208), .B(n_173), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_233), .A2(n_160), .B(n_178), .C(n_168), .Y(n_241) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_217), .A2(n_189), .B1(n_159), .B2(n_169), .C(n_161), .Y(n_242) );
OA22x2_ASAP7_75t_L g243 ( .A1(n_227), .A2(n_162), .B1(n_178), .B2(n_160), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_213), .A2(n_161), .B1(n_159), .B2(n_169), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_193), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_206), .A2(n_173), .B(n_167), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_224), .Y(n_247) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_208), .B(n_151), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_217), .B(n_151), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_211), .A2(n_141), .B1(n_145), .B2(n_147), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_194), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_194), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_217), .B(n_90), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_206), .A2(n_188), .B(n_167), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_197), .B(n_95), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_192), .A2(n_188), .B(n_183), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_192), .A2(n_188), .B(n_183), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_196), .A2(n_183), .B(n_185), .Y(n_258) );
O2A1O1Ixp5_ASAP7_75t_L g259 ( .A1(n_196), .A2(n_185), .B(n_165), .C(n_182), .Y(n_259) );
CKINVDCx8_ASAP7_75t_R g260 ( .A(n_230), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_225), .B(n_100), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_224), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g263 ( .A(n_226), .B(n_117), .C(n_126), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_198), .A2(n_185), .B(n_171), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_221), .B(n_179), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_221), .Y(n_266) );
INVx3_ASAP7_75t_SL g267 ( .A(n_225), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_197), .B(n_141), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_200), .B(n_141), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_211), .A2(n_141), .B1(n_145), .B2(n_147), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_SL g272 ( .A1(n_220), .A2(n_103), .B(n_182), .C(n_165), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_204), .B(n_147), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_195), .B(n_147), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_202), .Y(n_275) );
INVx5_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_201), .B(n_186), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_198), .A2(n_170), .B(n_171), .C(n_172), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_223), .A2(n_170), .B(n_172), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_219), .B(n_147), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_249), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_267), .B(n_203), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_228), .B(n_218), .C(n_222), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_244), .A2(n_232), .B1(n_209), .B2(n_210), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_244), .A2(n_236), .B1(n_212), .B2(n_207), .Y(n_285) );
AOI21xp33_ASAP7_75t_SL g286 ( .A1(n_238), .A2(n_234), .B(n_10), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_243), .A2(n_236), .B1(n_201), .B2(n_215), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_237), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_245), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_255), .A2(n_223), .B(n_220), .C(n_231), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_246), .A2(n_229), .B(n_216), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_256), .A2(n_229), .B(n_216), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_214), .B(n_235), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_264), .B(n_280), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_250), .A2(n_174), .A3(n_214), .B(n_235), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_242), .A2(n_141), .B(n_145), .C(n_147), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_237), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_261), .B(n_215), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_271), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_276), .B(n_201), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_252), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_278), .A2(n_215), .B(n_202), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_253), .B(n_201), .Y(n_305) );
AOI221xp5_ASAP7_75t_SL g306 ( .A1(n_250), .A2(n_215), .B1(n_202), .B2(n_145), .C(n_141), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_276), .B(n_202), .Y(n_307) );
AO31x2_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_174), .A3(n_145), .B(n_186), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_268), .A2(n_186), .B(n_179), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_270), .A2(n_145), .B(n_11), .C(n_13), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_274), .A2(n_186), .B(n_179), .C(n_14), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_248), .B(n_8), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_272), .A2(n_186), .B(n_179), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_260), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_266), .B(n_11), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_SL g316 ( .A1(n_269), .A2(n_48), .B(n_88), .C(n_87), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_284), .B(n_247), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_284), .B(n_248), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_289), .A2(n_266), .B1(n_262), .B2(n_239), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_283), .A2(n_259), .B(n_263), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_286), .A2(n_273), .B1(n_251), .B2(n_265), .C(n_254), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_281), .B(n_251), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_282), .B(n_262), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_282), .B(n_262), .Y(n_326) );
AO31x2_ASAP7_75t_L g327 ( .A1(n_296), .A2(n_275), .A3(n_279), .B(n_186), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_296), .A2(n_240), .B(n_186), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_299), .B(n_266), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
CKINVDCx9p33_ASAP7_75t_R g335 ( .A(n_312), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_283), .A2(n_277), .B(n_179), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_179), .B(n_45), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_315), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_311), .A2(n_179), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_293), .A2(n_47), .B(n_81), .Y(n_343) );
NOR2x1_ASAP7_75t_SL g344 ( .A(n_285), .B(n_43), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_292), .A2(n_50), .B(n_79), .Y(n_345) );
OA21x2_ASAP7_75t_L g346 ( .A1(n_306), .A2(n_42), .B(n_78), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_338), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_325), .A2(n_311), .B(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_325), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_338), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_329), .B(n_308), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_335), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_318), .B(n_308), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_340), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_331), .A2(n_291), .B(n_305), .Y(n_356) );
OAI33xp33_ASAP7_75t_L g357 ( .A1(n_321), .A2(n_287), .A3(n_310), .B1(n_297), .B2(n_288), .B3(n_290), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_331), .B(n_302), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_334), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_340), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_334), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_317), .B(n_287), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_336), .B(n_314), .Y(n_366) );
AOI21xp33_ASAP7_75t_SL g367 ( .A1(n_342), .A2(n_333), .B(n_324), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_344), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_318), .B(n_302), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_341), .B(n_307), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_320), .A2(n_309), .B(n_316), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
OAI31xp33_ASAP7_75t_L g375 ( .A1(n_326), .A2(n_332), .A3(n_319), .B(n_323), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_355), .Y(n_376) );
INVx4_ASAP7_75t_L g377 ( .A(n_372), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_354), .B(n_327), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_354), .B(n_327), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_362), .B(n_327), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_354), .B(n_328), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_362), .B(n_328), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_328), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
AND2x2_ASAP7_75t_SL g390 ( .A(n_347), .B(n_346), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_362), .B(n_351), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_352), .B(n_344), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_352), .B(n_346), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_352), .B(n_346), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_347), .B(n_346), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_359), .B(n_330), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_359), .B(n_330), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_330), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_350), .B(n_14), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_361), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_350), .B(n_15), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_360), .B(n_18), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_379), .B(n_355), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_406), .B(n_358), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_379), .B(n_360), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_406), .B(n_358), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_407), .B(n_410), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_406), .B(n_374), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_387), .B(n_358), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_410), .B(n_360), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_408), .B(n_409), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_407), .B(n_360), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_408), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_408), .B(n_358), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_409), .B(n_370), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_409), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_377), .B(n_366), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_379), .B(n_364), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_364), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_380), .B(n_364), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_376), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_376), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_363), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_389), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_395), .B(n_396), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_380), .B(n_369), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_396), .B(n_370), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_403), .B(n_371), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_391), .B(n_370), .Y(n_449) );
AND2x4_ASAP7_75t_SL g450 ( .A(n_377), .B(n_353), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_387), .B(n_363), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_383), .B(n_369), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_383), .B(n_363), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_391), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_394), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_404), .B(n_369), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_383), .B(n_371), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_392), .A2(n_375), .B1(n_353), .B2(n_357), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_402), .B(n_365), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_435), .B(n_367), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_450), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_439), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_436), .B(n_437), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_450), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_436), .B(n_402), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_421), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_437), .B(n_392), .Y(n_470) );
NAND2x1_ASAP7_75t_SL g471 ( .A(n_434), .B(n_401), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_438), .B(n_404), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_401), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_430), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_459), .B(n_375), .C(n_367), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_412), .Y(n_476) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_447), .A2(n_367), .B(n_366), .C(n_392), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_442), .B(n_365), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_425), .B(n_398), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_412), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_438), .B(n_393), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_416), .B(n_393), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_425), .B(n_398), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_415), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_458), .B(n_404), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_451), .B(n_405), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_461), .B(n_381), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_454), .B(n_381), .Y(n_488) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_448), .B(n_377), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_416), .B(n_393), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_449), .B(n_385), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_446), .B(n_385), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_446), .B(n_397), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_452), .B(n_397), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_451), .B(n_405), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_452), .B(n_397), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_453), .B(n_405), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_429), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_419), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_417), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_411), .B(n_403), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_419), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_453), .B(n_394), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_411), .B(n_394), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_414), .B(n_378), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_425), .B(n_378), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_420), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_457), .B(n_377), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_422), .Y(n_511) );
NAND4xp25_ASAP7_75t_SL g512 ( .A(n_427), .B(n_399), .C(n_337), .D(n_298), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_378), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_448), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_378), .Y(n_515) );
OAI33xp33_ASAP7_75t_L g516 ( .A1(n_433), .A2(n_19), .A3(n_357), .B1(n_348), .B2(n_368), .B3(n_390), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_418), .B(n_356), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_460), .B(n_368), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_432), .B(n_374), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_460), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_426), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_520), .B(n_443), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_464), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_464), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_514), .B(n_448), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_470), .B(n_413), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_484), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_467), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_484), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_502), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_467), .A2(n_448), .B1(n_423), .B2(n_431), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_466), .B(n_428), .Y(n_534) );
OAI222xp33_ASAP7_75t_L g535 ( .A1(n_489), .A2(n_423), .B1(n_445), .B2(n_440), .C1(n_413), .C2(n_444), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_498), .B(n_423), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_521), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_498), .B(n_413), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_509), .Y(n_539) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_479), .B(n_441), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_492), .B(n_428), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_511), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
NAND2xp33_ASAP7_75t_R g544 ( .A(n_479), .B(n_426), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_465), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_470), .B(n_455), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_478), .B(n_455), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_472), .B(n_424), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_476), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_480), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_478), .B(n_424), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_481), .B(n_399), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_481), .B(n_348), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_482), .B(n_399), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_475), .A2(n_316), .B(n_374), .C(n_372), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_491), .B(n_348), .Y(n_557) );
AOI21xp33_ASAP7_75t_SL g558 ( .A1(n_462), .A2(n_477), .B(n_518), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_494), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_482), .B(n_348), .Y(n_560) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_471), .A2(n_339), .B(n_345), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_490), .B(n_348), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_462), .B(n_374), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_493), .B(n_348), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_479), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_500), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_473), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_499), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_495), .B(n_348), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
INVxp33_ASAP7_75t_L g572 ( .A(n_518), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_483), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_490), .B(n_356), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_544), .A2(n_510), .B1(n_517), .B2(n_474), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_548), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_540), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_574), .B(n_497), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_545), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_535), .A2(n_516), .B(n_483), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_560), .B(n_515), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_560), .A2(n_487), .B1(n_488), .B2(n_515), .C1(n_468), .C2(n_503), .Y(n_584) );
NOR3xp33_ASAP7_75t_SL g585 ( .A(n_544), .B(n_512), .C(n_343), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_523), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_562), .B(n_506), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_542), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_558), .B(n_508), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_550), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_540), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_565), .B(n_508), .Y(n_593) );
AOI32xp33_ASAP7_75t_L g594 ( .A1(n_572), .A2(n_503), .A3(n_483), .B1(n_513), .B2(n_506), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_565), .B(n_519), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_572), .A2(n_507), .B1(n_486), .B2(n_501), .C(n_496), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_525), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_530), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_541), .B(n_504), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_538), .B(n_504), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_562), .B(n_501), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_563), .A2(n_372), .B(n_322), .C(n_373), .Y(n_605) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_563), .A2(n_372), .B(n_373), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_569), .B(n_356), .Y(n_607) );
OAI21xp33_ASAP7_75t_SL g608 ( .A1(n_573), .A2(n_390), .B(n_373), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_571), .B(n_356), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
AOI322xp5_ASAP7_75t_L g611 ( .A1(n_590), .A2(n_553), .A3(n_555), .B1(n_537), .B2(n_567), .C1(n_538), .C2(n_554), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_590), .A2(n_526), .B1(n_533), .B2(n_568), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_591), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_579), .A2(n_573), .B1(n_526), .B2(n_536), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_584), .B(n_527), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_586), .Y(n_616) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_582), .A2(n_573), .B(n_556), .C(n_564), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_575), .A2(n_526), .B(n_522), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_579), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_524), .B(n_547), .C(n_552), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_592), .A2(n_536), .B1(n_570), .B2(n_549), .Y(n_621) );
NOR2xp67_ASAP7_75t_L g622 ( .A(n_581), .B(n_528), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_597), .B(n_553), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_598), .A2(n_546), .A3(n_555), .B1(n_557), .B2(n_531), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_599), .A2(n_561), .B(n_543), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_610), .B(n_543), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_594), .A2(n_531), .B1(n_529), .B2(n_561), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_606), .A2(n_529), .B(n_301), .C(n_561), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
AOI221xp5_ASAP7_75t_SL g630 ( .A1(n_576), .A2(n_20), .B1(n_21), .B2(n_22), .C(n_23), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_576), .A2(n_373), .B(n_356), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_577), .B(n_373), .Y(n_632) );
OAI221xp5_ASAP7_75t_SL g633 ( .A1(n_611), .A2(n_608), .B1(n_581), .B2(n_607), .C(n_609), .Y(n_633) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_616), .B(n_593), .Y(n_634) );
OAI21xp33_ASAP7_75t_SL g635 ( .A1(n_622), .A2(n_596), .B(n_587), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_627), .A2(n_588), .B1(n_589), .B2(n_578), .C(n_602), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_619), .A2(n_585), .B1(n_601), .B2(n_604), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_618), .B(n_605), .C(n_585), .D(n_583), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_615), .B(n_580), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_614), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_620), .A2(n_618), .B(n_621), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_617), .A2(n_603), .B1(n_600), .B2(n_313), .C(n_390), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_625), .A2(n_373), .B(n_356), .C(n_313), .Y(n_643) );
AND4x1_ASAP7_75t_L g644 ( .A(n_612), .B(n_24), .C(n_25), .D(n_29), .Y(n_644) );
AND4x2_ASAP7_75t_L g645 ( .A(n_624), .B(n_30), .C(n_31), .D(n_32), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_633), .A2(n_623), .B(n_628), .C(n_631), .Y(n_646) );
NOR5xp2_ASAP7_75t_L g647 ( .A(n_638), .B(n_629), .C(n_613), .D(n_630), .E(n_626), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_641), .A2(n_637), .B1(n_640), .B2(n_635), .C(n_642), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_636), .B(n_632), .C(n_373), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_639), .A2(n_34), .B(n_35), .C(n_37), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_634), .B(n_38), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_643), .A2(n_39), .B(n_51), .C(n_52), .Y(n_652) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_648), .A2(n_645), .B(n_644), .C(n_59), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_647), .B(n_55), .C(n_56), .D(n_62), .Y(n_654) );
XNOR2x1_ASAP7_75t_L g655 ( .A(n_649), .B(n_356), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_651), .B(n_63), .C(n_64), .D(n_65), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_653), .B(n_646), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g658 ( .A(n_654), .B(n_650), .C(n_652), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_660), .Y(n_662) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_660), .A2(n_658), .B1(n_655), .B2(n_68), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_661), .B(n_67), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_664), .Y(n_665) );
AO221x1_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_662), .B1(n_69), .B2(n_70), .C(n_72), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_66), .B(n_74), .C(n_85), .Y(n_667) );
endmodule