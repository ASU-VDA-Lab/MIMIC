module fake_netlist_6_3504_n_2367 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2367);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2367;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2090;
wire n_2058;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_399),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_439),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_315),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_5),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_253),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_277),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_378),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_128),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_396),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_117),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_145),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_457),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_359),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_63),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_295),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_3),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_35),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_37),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_33),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_145),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_51),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_2),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_257),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_174),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_317),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_412),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_136),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_99),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_49),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_94),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_130),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_205),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_114),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_318),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_135),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_237),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_231),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_99),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_124),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_184),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_417),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_0),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_270),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_60),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_493),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_45),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_224),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_87),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_259),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_346),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_245),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_333),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_319),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_233),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_0),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_254),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_454),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_477),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_490),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_358),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_36),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_226),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_124),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_236),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_498),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_349),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_234),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_106),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_208),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_492),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_310),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_51),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_235),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_324),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_503),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_496),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_456),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_34),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_377),
.Y(n_605)
);

BUFx5_ASAP7_75t_L g606 ( 
.A(n_325),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_240),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_160),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_96),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_313),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_362),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_352),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_488),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_134),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_122),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_211),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g618 ( 
.A(n_302),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_485),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_311),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_138),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_357),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_506),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_244),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_134),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_405),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_200),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_52),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_221),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_102),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_495),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_167),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_502),
.Y(n_633)
);

BUFx5_ASAP7_75t_L g634 ( 
.A(n_176),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_198),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_188),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_105),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_135),
.Y(n_638)
);

BUFx8_ASAP7_75t_SL g639 ( 
.A(n_472),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_480),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_296),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_78),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_314),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_282),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_344),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_432),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_351),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_28),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_165),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_504),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_96),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_334),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_509),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_281),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_510),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_107),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_19),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_491),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_342),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_102),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_94),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_21),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_449),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_243),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_89),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_275),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_445),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_420),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_331),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_410),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_20),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_403),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_223),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_306),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_64),
.Y(n_675)
);

CKINVDCx16_ASAP7_75t_R g676 ( 
.A(n_501),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_184),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_16),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_45),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_252),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_416),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_447),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_430),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_292),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_133),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_210),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_427),
.Y(n_687)
);

CKINVDCx14_ASAP7_75t_R g688 ( 
.A(n_177),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_508),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_75),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_71),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_42),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_77),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_218),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_192),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_8),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_22),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_500),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_379),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_360),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_223),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_286),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_340),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_436),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_441),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_148),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_327),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_497),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_63),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_303),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_40),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_86),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_182),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_345),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_519),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_168),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_213),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_202),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_191),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_494),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_177),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_182),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_47),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_109),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_38),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_185),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_17),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_191),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_297),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_380),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_28),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_24),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_48),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_266),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_507),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_168),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_44),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_196),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_330),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_634),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_634),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_634),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_634),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_543),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_634),
.Y(n_746)
);

CKINVDCx14_ASAP7_75t_R g747 ( 
.A(n_688),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_564),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_581),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_564),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_564),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_606),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_521),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_627),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_564),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_559),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_673),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_580),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_617),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_617),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_617),
.Y(n_762)
);

INVxp33_ASAP7_75t_SL g763 ( 
.A(n_581),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_724),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_724),
.Y(n_766)
);

INVxp33_ASAP7_75t_L g767 ( 
.A(n_616),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_612),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_724),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_717),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_522),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_724),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_614),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_580),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_629),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_632),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_533),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_596),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_688),
.B(n_1),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_539),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_546),
.Y(n_781)
);

INVxp33_ASAP7_75t_SL g782 ( 
.A(n_612),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_557),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_562),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_563),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_523),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_565),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_589),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_534),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_538),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_592),
.Y(n_791)
);

INVxp33_ASAP7_75t_SL g792 ( 
.A(n_525),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_594),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_608),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_625),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_630),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_642),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_649),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_679),
.Y(n_799)
);

INVxp33_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_675),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_686),
.Y(n_802)
);

CKINVDCx14_ASAP7_75t_R g803 ( 
.A(n_540),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_735),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_735),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_718),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_719),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_723),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_550),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_725),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_693),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_524),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_606),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_526),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_551),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_576),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_527),
.Y(n_819)
);

BUFx2_ASAP7_75t_SL g820 ( 
.A(n_530),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_535),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_536),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_529),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_675),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_542),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_548),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_532),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_570),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_622),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_584),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_590),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_537),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_586),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_593),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_599),
.Y(n_835)
);

INVxp33_ASAP7_75t_SL g836 ( 
.A(n_544),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_626),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_748),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_758),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_758),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_758),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_743),
.A2(n_734),
.B(n_668),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_758),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_774),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_832),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_753),
.B(n_583),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_771),
.B(n_591),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_786),
.B(n_610),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_774),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_750),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_789),
.B(n_647),
.Y(n_851)
);

OA21x2_ASAP7_75t_L g852 ( 
.A1(n_740),
.A2(n_603),
.B(n_601),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_756),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_751),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_790),
.B(n_655),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_805),
.B(n_714),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_747),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_747),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_778),
.B(n_640),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_774),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_755),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_759),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_811),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_774),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_761),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_762),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_743),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_817),
.B(n_615),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_806),
.B(n_619),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_620),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_749),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_746),
.Y(n_872)
);

AND2x2_ASAP7_75t_SL g873 ( 
.A(n_779),
.B(n_653),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_764),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_746),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_741),
.A2(n_645),
.B(n_623),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_742),
.A2(n_652),
.B(n_650),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_765),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_782),
.A2(n_676),
.B1(n_658),
.B2(n_633),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_813),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_831),
.B(n_837),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_752),
.A2(n_659),
.B(n_654),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_766),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_752),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_744),
.Y(n_885)
);

BUFx8_ASAP7_75t_SL g886 ( 
.A(n_745),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_769),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_772),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_760),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_760),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_815),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_815),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_814),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_756),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_775),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_776),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

INVx6_ASAP7_75t_L g898 ( 
.A(n_829),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_819),
.Y(n_899)
);

OA21x2_ASAP7_75t_L g900 ( 
.A1(n_821),
.A2(n_666),
.B(n_664),
.Y(n_900)
);

OA21x2_ASAP7_75t_L g901 ( 
.A1(n_822),
.A2(n_674),
.B(n_669),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_825),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_869),
.B(n_768),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_872),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_872),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_873),
.A2(n_782),
.B1(n_791),
.B2(n_779),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_875),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_875),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_839),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_897),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_885),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_839),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_875),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_885),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_881),
.B(n_792),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_890),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_890),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_890),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_880),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_889),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_889),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_842),
.A2(n_828),
.B(n_826),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_889),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_882),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_882),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_867),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_838),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_839),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_868),
.B(n_636),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_867),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_853),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_867),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_899),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_839),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_871),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_839),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_899),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_864),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_864),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_899),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_881),
.B(n_830),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_887),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_886),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_899),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_864),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_891),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_899),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_855),
.B(n_792),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_887),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_881),
.B(n_780),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_895),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_871),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_895),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_891),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_873),
.B(n_823),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_864),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_891),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_891),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_891),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_893),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_892),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_892),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_864),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_892),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_893),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_838),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_902),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_859),
.B(n_823),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_853),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_892),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_850),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_894),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_902),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_892),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_843),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_894),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_841),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_842),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_843),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_883),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_850),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_840),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_840),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_843),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_844),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_860),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_950),
.Y(n_989)
);

BUFx8_ASAP7_75t_SL g990 ( 
.A(n_937),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_919),
.B(n_857),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_971),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_906),
.B(n_845),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_928),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_971),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_920),
.B(n_921),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_903),
.B(n_857),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_952),
.B(n_846),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_L g999 ( 
.A(n_980),
.B(n_847),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_915),
.B(n_827),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_921),
.B(n_923),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_928),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_923),
.B(n_856),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_982),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_968),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_952),
.B(n_848),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_952),
.A2(n_869),
.B1(n_870),
.B2(n_763),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_907),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_980),
.Y(n_1009)
);

HAxp5_ASAP7_75t_SL g1010 ( 
.A(n_957),
.B(n_879),
.CON(n_1010),
.SN(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_932),
.B(n_827),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_903),
.B(n_870),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_984),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_968),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_974),
.B(n_856),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_943),
.B(n_856),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_909),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_978),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_980),
.B(n_851),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_984),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_978),
.B(n_820),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_937),
.B(n_898),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_953),
.Y(n_1023)
);

BUFx4f_ASAP7_75t_L g1024 ( 
.A(n_955),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_910),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_930),
.B(n_858),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_973),
.B(n_858),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_962),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_973),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_930),
.B(n_863),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_970),
.B(n_863),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_907),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_983),
.B(n_767),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_983),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_967),
.B(n_767),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_969),
.Y(n_1036)
);

INVxp67_ASAP7_75t_SL g1037 ( 
.A(n_979),
.Y(n_1037)
);

BUFx10_ASAP7_75t_L g1038 ( 
.A(n_975),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_911),
.B(n_852),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_922),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_980),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_914),
.B(n_979),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_982),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_979),
.B(n_836),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_925),
.B(n_852),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_908),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_922),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_954),
.B(n_770),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_925),
.B(n_836),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_945),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_944),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_944),
.B(n_770),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_951),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_951),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_908),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_985),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_924),
.A2(n_901),
.B1(n_900),
.B2(n_876),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_927),
.B(n_803),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_934),
.B(n_781),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_980),
.B(n_531),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_924),
.B(n_606),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_977),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_931),
.B(n_852),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_926),
.B(n_580),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_939),
.B(n_585),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_988),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_942),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_913),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_988),
.Y(n_1070)
);

INVx4_ASAP7_75t_SL g1071 ( 
.A(n_926),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_933),
.B(n_876),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_905),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_905),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_946),
.B(n_600),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_904),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_933),
.B(n_898),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_904),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_981),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_949),
.A2(n_901),
.B1(n_900),
.B2(n_877),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_913),
.B(n_876),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_916),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_935),
.B(n_876),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_916),
.B(n_777),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_909),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_917),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_935),
.B(n_877),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_956),
.B(n_877),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_917),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_918),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_909),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_918),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_956),
.A2(n_900),
.B1(n_901),
.B2(n_877),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_959),
.B(n_898),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_959),
.B(n_624),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_986),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_948),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_948),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_961),
.A2(n_901),
.B1(n_900),
.B2(n_689),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_961),
.B(n_860),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_987),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_972),
.B(n_844),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_972),
.A2(n_698),
.B1(n_700),
.B2(n_682),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_976),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_976),
.B(n_801),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_909),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_909),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_948),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_960),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_982),
.B(n_528),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_960),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_912),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_960),
.B(n_783),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_963),
.A2(n_703),
.B1(n_618),
.B2(n_606),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_982),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_963),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_912),
.Y(n_1117)
);

AND2x6_ASAP7_75t_L g1118 ( 
.A(n_963),
.B(n_580),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_964),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_982),
.B(n_720),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_912),
.B(n_896),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_964),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1000),
.A2(n_556),
.B1(n_692),
.B2(n_552),
.C(n_541),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1016),
.B(n_964),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1012),
.B(n_896),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1013),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1010),
.B(n_896),
.C(n_824),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1073),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1012),
.B(n_966),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1037),
.B(n_966),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_994),
.B(n_966),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1003),
.A2(n_993),
.B1(n_1001),
.B2(n_996),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1002),
.A2(n_834),
.B(n_835),
.C(n_833),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_990),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1018),
.B(n_561),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1022),
.B(n_898),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_999),
.A2(n_884),
.B(n_912),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1074),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1009),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1018),
.B(n_566),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1005),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1020),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1064),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1064),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1014),
.B(n_958),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_989),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1029),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1033),
.B(n_745),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1023),
.B(n_568),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1023),
.B(n_574),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_L g1156 ( 
.A(n_991),
.B(n_773),
.C(n_716),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1034),
.B(n_938),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_995),
.B(n_784),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1024),
.B(n_575),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1053),
.B(n_941),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1051),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1104),
.B(n_941),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1024),
.B(n_577),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1104),
.B(n_947),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_998),
.A2(n_733),
.B1(n_706),
.B2(n_579),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1084),
.B(n_929),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_997),
.B(n_578),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_989),
.B(n_754),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1052),
.B(n_1035),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1060),
.A2(n_618),
.B1(n_715),
.B2(n_606),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1008),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1011),
.B(n_754),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1015),
.B(n_597),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1054),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1006),
.A2(n_678),
.B(n_677),
.C(n_709),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1101),
.B(n_912),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1105),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_996),
.A2(n_1001),
.B1(n_1059),
.B2(n_1113),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_L g1179 ( 
.A(n_1041),
.B(n_618),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1059),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1015),
.B(n_605),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1048),
.B(n_757),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1101),
.B(n_936),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1032),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_SL g1185 ( 
.A(n_1022),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1025),
.A2(n_757),
.B1(n_800),
.B2(n_777),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1049),
.B(n_940),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1122),
.B(n_940),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1022),
.B(n_785),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1122),
.B(n_941),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1021),
.B(n_800),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1044),
.B(n_639),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1007),
.B(n_607),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1046),
.Y(n_1194)
);

XOR2xp5_ASAP7_75t_L g1195 ( 
.A(n_1050),
.B(n_611),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_992),
.B(n_773),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1113),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1027),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1027),
.B(n_613),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1036),
.B(n_639),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1076),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1031),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1055),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1069),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1028),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1038),
.B(n_697),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1089),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1019),
.A2(n_641),
.B1(n_643),
.B2(n_631),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1056),
.B(n_947),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1041),
.B(n_644),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1038),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1078),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1067),
.B(n_958),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1085),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1079),
.B(n_646),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1058),
.A2(n_602),
.B1(n_683),
.B2(n_540),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_L g1218 ( 
.A(n_1026),
.B(n_788),
.C(n_787),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1068),
.B(n_545),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1082),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1079),
.B(n_663),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_1040),
.B(n_582),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1077),
.B(n_1096),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1062),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1043),
.B(n_670),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1094),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1121),
.B(n_547),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1042),
.B(n_965),
.Y(n_1228)
);

NOR2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1039),
.B(n_549),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1066),
.B(n_554),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1085),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1075),
.B(n_555),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1039),
.A2(n_874),
.B(n_878),
.C(n_866),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1043),
.B(n_672),
.Y(n_1234)
);

INVxp33_ASAP7_75t_L g1235 ( 
.A(n_1030),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1043),
.B(n_680),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1086),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1099),
.B(n_941),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1095),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1085),
.B(n_681),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1070),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1092),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1094),
.B(n_558),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1094),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1111),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1110),
.B(n_560),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1116),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1109),
.B(n_929),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1119),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1120),
.B(n_793),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1004),
.B(n_1115),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1091),
.B(n_687),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1004),
.B(n_936),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1115),
.B(n_936),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1071),
.B(n_794),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1091),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1103),
.A2(n_715),
.B1(n_618),
.B2(n_667),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1091),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1097),
.B(n_938),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1098),
.B(n_938),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1114),
.A2(n_569),
.B1(n_572),
.B2(n_571),
.C(n_567),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1108),
.B(n_965),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1112),
.B(n_699),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1045),
.B(n_929),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1100),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1081),
.B(n_697),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1106),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1112),
.B(n_702),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1102),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1063),
.B(n_938),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1081),
.B(n_795),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1061),
.A2(n_1083),
.B1(n_1087),
.B2(n_1072),
.Y(n_1272)
);

INVx8_ASAP7_75t_L g1273 ( 
.A(n_1112),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1106),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1071),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1107),
.B(n_796),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1088),
.B(n_947),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1093),
.B(n_797),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1107),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1117),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1017),
.B(n_798),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1117),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1057),
.B(n_965),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1017),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1047),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1065),
.B(n_965),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1080),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1065),
.B(n_704),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1065),
.B(n_708),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1065),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1118),
.B(n_573),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1118),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1118),
.B(n_936),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1118),
.B(n_710),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1016),
.B(n_938),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1016),
.B(n_940),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1013),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1073),
.Y(n_1298)
);

OAI22x1_ASAP7_75t_L g1299 ( 
.A1(n_1000),
.A2(n_587),
.B1(n_595),
.B2(n_588),
.Y(n_1299)
);

BUFx5_ASAP7_75t_L g1300 ( 
.A(n_1040),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1073),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1013),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1012),
.B(n_729),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1016),
.B(n_936),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_989),
.B(n_598),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1073),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1016),
.B(n_940),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1012),
.B(n_730),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1073),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_991),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1016),
.B(n_940),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1000),
.A2(n_604),
.B1(n_628),
.B2(n_621),
.C(n_609),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1073),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1009),
.B(n_618),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1012),
.B(n_739),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1016),
.B(n_947),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1016),
.B(n_947),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_991),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1016),
.B(n_958),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1013),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1134),
.B(n_878),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1169),
.B(n_888),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1196),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1266),
.B(n_888),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1153),
.B(n_1310),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1191),
.B(n_799),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1215),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1244),
.B(n_802),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1177),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1172),
.A2(n_861),
.B1(n_862),
.B2(n_854),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1182),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1229),
.A2(n_861),
.B1(n_862),
.B2(n_854),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1138),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1226),
.B(n_958),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1175),
.A2(n_1246),
.B(n_1232),
.C(n_1230),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1198),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1241),
.Y(n_1337)
);

NAND2x1_ASAP7_75t_L g1338 ( 
.A(n_1127),
.B(n_958),
.Y(n_1338)
);

NOR3xp33_ASAP7_75t_SL g1339 ( 
.A(n_1129),
.B(n_637),
.C(n_635),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1178),
.B(n_865),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1165),
.A2(n_638),
.B1(n_656),
.B2(n_648),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1318),
.B(n_804),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1123),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1124),
.A2(n_715),
.B1(n_582),
.B2(n_705),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1197),
.A2(n_715),
.B1(n_582),
.B2(n_705),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1206),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1143),
.B(n_865),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1150),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1271),
.B(n_1223),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1130),
.B(n_1140),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1202),
.A2(n_1168),
.B1(n_1217),
.B2(n_1136),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1298),
.B(n_866),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1226),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1215),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1301),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1149),
.A2(n_661),
.B1(n_662),
.B2(n_657),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1306),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1224),
.B(n_807),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1165),
.B(n_665),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1189),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1205),
.B(n_808),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1189),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1275),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1138),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1219),
.B(n_809),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1309),
.B(n_874),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1313),
.B(n_671),
.Y(n_1367)
);

BUFx4f_ASAP7_75t_L g1368 ( 
.A(n_1189),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1180),
.B(n_810),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1161),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1156),
.B(n_812),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1158),
.Y(n_1372)
);

BUFx4f_ASAP7_75t_SL g1373 ( 
.A(n_1137),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1174),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1128),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1227),
.A2(n_849),
.B(n_844),
.C(n_651),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1255),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1276),
.A2(n_1278),
.B1(n_1308),
.B2(n_1303),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1201),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1265),
.B(n_1176),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1144),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1213),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1185),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1186),
.B(n_602),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1273),
.Y(n_1385)
);

BUFx4f_ASAP7_75t_L g1386 ( 
.A(n_1281),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1211),
.B(n_683),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1183),
.B(n_690),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1305),
.Y(n_1389)
);

NOR3xp33_ASAP7_75t_L g1390 ( 
.A(n_1192),
.B(n_695),
.C(n_691),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1220),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1166),
.B(n_696),
.Y(n_1392)
);

NOR3xp33_ASAP7_75t_SL g1393 ( 
.A(n_1199),
.B(n_1200),
.C(n_1243),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1160),
.B(n_701),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1239),
.A2(n_707),
.B1(n_684),
.B2(n_715),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1145),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1281),
.B(n_1273),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1273),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1276),
.A2(n_582),
.B1(n_705),
.B2(n_667),
.Y(n_1399)
);

AND2x6_ASAP7_75t_L g1400 ( 
.A(n_1287),
.B(n_667),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1237),
.Y(n_1401)
);

INVx5_ASAP7_75t_L g1402 ( 
.A(n_1215),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1269),
.B(n_1131),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1242),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1315),
.A2(n_1167),
.B1(n_1181),
.B2(n_1173),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1195),
.A2(n_712),
.B1(n_713),
.B2(n_711),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1235),
.A2(n_726),
.B1(n_727),
.B2(n_721),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1158),
.B(n_731),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1187),
.B(n_732),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1142),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_SL g1411 ( 
.A(n_1312),
.B(n_737),
.C(n_736),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1320),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1193),
.A2(n_705),
.B1(n_707),
.B2(n_684),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1264),
.A2(n_884),
.B(n_841),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1255),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1250),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1146),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1299),
.A2(n_738),
.B1(n_660),
.B2(n_728),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1238),
.A2(n_1272),
.B(n_1283),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1284),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1171),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1231),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1147),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1297),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1272),
.B(n_553),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1218),
.B(n_1),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1126),
.B(n_238),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1302),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1231),
.B(n_883),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1261),
.B(n_2),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1295),
.B(n_849),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1184),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1194),
.B(n_239),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1203),
.Y(n_1434)
);

OR2x4_ASAP7_75t_L g1435 ( 
.A(n_1291),
.B(n_883),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1204),
.B(n_3),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1207),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1212),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1256),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1296),
.B(n_1304),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1307),
.B(n_1311),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1185),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1256),
.B(n_883),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1316),
.B(n_849),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1256),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1447)
);

INVx5_ASAP7_75t_L g1448 ( 
.A(n_1258),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1285),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_SL g1450 ( 
.A(n_1208),
.B(n_4),
.C(n_5),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1245),
.Y(n_1451)
);

AND2x2_ASAP7_75t_SL g1452 ( 
.A(n_1170),
.B(n_4),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1159),
.B(n_1163),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1125),
.B(n_883),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1247),
.B(n_241),
.Y(n_1455)
);

INVx5_ASAP7_75t_L g1456 ( 
.A(n_1258),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1258),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1208),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1162),
.B(n_6),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1164),
.B(n_7),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1249),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1133),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1148),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1210),
.B(n_8),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_R g1465 ( 
.A(n_1127),
.B(n_242),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1267),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1216),
.B(n_884),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1240),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1221),
.B(n_9),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1279),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1274),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1157),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1270),
.B(n_9),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1252),
.A2(n_884),
.B1(n_12),
.B2(n_10),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1263),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1280),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1268),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1277),
.B(n_11),
.Y(n_1478)
);

BUFx4f_ASAP7_75t_L g1479 ( 
.A(n_1282),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1141),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1209),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1214),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1135),
.B(n_1233),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_SL g1484 ( 
.A(n_1225),
.B(n_13),
.C(n_14),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1141),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_L g1486 ( 
.A(n_1300),
.B(n_246),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1234),
.B(n_13),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1259),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1151),
.B(n_1152),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1151),
.B(n_14),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1152),
.B(n_247),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1188),
.B(n_15),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1236),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1190),
.B(n_15),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1260),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1262),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1222),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1497)
);

BUFx4f_ASAP7_75t_L g1498 ( 
.A(n_1292),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1248),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1251),
.B(n_18),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1222),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1132),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1288),
.A2(n_1289),
.B1(n_1314),
.B2(n_1179),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1300),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1294),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1228),
.B(n_19),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1290),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1507)
);

AOI21xp33_ASAP7_75t_L g1508 ( 
.A1(n_1286),
.A2(n_23),
.B(n_24),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1293),
.B(n_23),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1300),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1300),
.B(n_25),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1257),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1300),
.B(n_251),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1253),
.B(n_25),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1222),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1254),
.B(n_255),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1222),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1139),
.B(n_26),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1169),
.B(n_256),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1134),
.B(n_27),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1143),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1241),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1198),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1359),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1524)
);

BUFx2_ASAP7_75t_SL g1525 ( 
.A(n_1398),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1491),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1348),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1491),
.Y(n_1528)
);

AOI21xp33_ASAP7_75t_L g1529 ( 
.A1(n_1335),
.A2(n_30),
.B(n_31),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1458),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1355),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1357),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1521),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1389),
.B(n_32),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1349),
.B(n_35),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1419),
.A2(n_260),
.B(n_258),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1350),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1331),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1370),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1449),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1398),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1374),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1379),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1326),
.B(n_39),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1403),
.B(n_39),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1325),
.B(n_1365),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1416),
.B(n_40),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1410),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1380),
.B(n_41),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1441),
.A2(n_262),
.B(n_261),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1327),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1386),
.B(n_43),
.Y(n_1552)
);

AND2x4_ASAP7_75t_SL g1553 ( 
.A(n_1385),
.B(n_263),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1411),
.A2(n_47),
.B1(n_44),
.B2(n_46),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1364),
.B(n_520),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1382),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1469),
.A2(n_49),
.B(n_46),
.C(n_48),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1391),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1502),
.B(n_50),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1329),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1430),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1336),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1327),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1401),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1404),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1337),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1452),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1512),
.B(n_54),
.Y(n_1569)
);

BUFx8_ASAP7_75t_L g1570 ( 
.A(n_1360),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1408),
.B(n_55),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1327),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1432),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1398),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1523),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1434),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1436),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1439),
.B(n_1322),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1372),
.B(n_1493),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1453),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1394),
.B(n_59),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1347),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1352),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1402),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1451),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1341),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1324),
.B(n_61),
.Y(n_1587)
);

AND3x1_ASAP7_75t_SL g1588 ( 
.A(n_1406),
.B(n_62),
.C(n_64),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1366),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1477),
.B(n_62),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1390),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1591)
);

XNOR2xp5_ASAP7_75t_L g1592 ( 
.A(n_1351),
.B(n_264),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1427),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1388),
.B(n_68),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1354),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1471),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1520),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1476),
.Y(n_1598)
);

OAI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1373),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1462),
.B(n_72),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1461),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1343),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1409),
.B(n_72),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1412),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1363),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1375),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1463),
.B(n_73),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1472),
.B(n_73),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1381),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1354),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1321),
.A2(n_1425),
.B(n_1442),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1420),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1402),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1377),
.B(n_265),
.Y(n_1614)
);

AND2x6_ASAP7_75t_L g1615 ( 
.A(n_1504),
.B(n_267),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1354),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1450),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1342),
.B(n_74),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1418),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1333),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1323),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1371),
.B(n_79),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1397),
.B(n_268),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1346),
.B(n_79),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1519),
.B(n_80),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1519),
.B(n_80),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1397),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1468),
.B(n_81),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1328),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_L g1630 ( 
.A(n_1415),
.B(n_269),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1362),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1447),
.B(n_1460),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1392),
.B(n_81),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1402),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1481),
.B(n_82),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1428),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1384),
.A2(n_82),
.B(n_83),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1482),
.B(n_83),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1368),
.B(n_84),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1328),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1494),
.B(n_84),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1448),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1446),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1506),
.B(n_85),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1396),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1427),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1417),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1385),
.B(n_271),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1423),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1488),
.B(n_88),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1369),
.B(n_518),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1495),
.B(n_88),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1499),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1358),
.B(n_89),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1383),
.B(n_1443),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1424),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1466),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1358),
.B(n_90),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1361),
.B(n_1369),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1339),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1361),
.B(n_90),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1470),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1393),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1405),
.B(n_91),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1421),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1448),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1422),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1499),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1496),
.B(n_91),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1426),
.B(n_92),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1499),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1433),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1448),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1500),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1438),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1353),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1490),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1378),
.A2(n_97),
.B(n_93),
.C(n_95),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1480),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1464),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1455),
.B(n_272),
.Y(n_1681)
);

CKINVDCx11_ASAP7_75t_R g1682 ( 
.A(n_1455),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1456),
.B(n_273),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1437),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1459),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1367),
.B(n_97),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1492),
.B(n_98),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1465),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1433),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1489),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1456),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1479),
.Y(n_1692)
);

AND2x6_ASAP7_75t_SL g1693 ( 
.A(n_1489),
.B(n_98),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1440),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1514),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1456),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1334),
.B(n_274),
.Y(n_1697)
);

BUFx12f_ASAP7_75t_L g1698 ( 
.A(n_1487),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1484),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1440),
.B(n_276),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1457),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1457),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1475),
.A2(n_103),
.B1(n_100),
.B2(n_101),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1485),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1473),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1478),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1498),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1330),
.B(n_1340),
.Y(n_1708)
);

AND3x1_ASAP7_75t_SL g1709 ( 
.A(n_1497),
.B(n_100),
.C(n_101),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1413),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.C(n_107),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1429),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1509),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1511),
.Y(n_1713)
);

AOI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1687),
.A2(n_1454),
.B(n_1445),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1536),
.A2(n_1431),
.B(n_1510),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1531),
.Y(n_1716)
);

AOI211x1_ASAP7_75t_L g1717 ( 
.A1(n_1599),
.A2(n_1508),
.B(n_1387),
.C(n_1518),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1707),
.B(n_1516),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_SL g1719 ( 
.A(n_1525),
.B(n_1513),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1550),
.A2(n_1414),
.B(n_1713),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1632),
.A2(n_1486),
.B(n_1467),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1672),
.A2(n_1338),
.B(n_1483),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1611),
.A2(n_1503),
.B(n_1435),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1672),
.A2(n_1444),
.B(n_1700),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1546),
.B(n_1395),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1708),
.A2(n_1516),
.B(n_1501),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1582),
.B(n_1332),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1583),
.B(n_1474),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1532),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1533),
.Y(n_1730)
);

AOI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1664),
.A2(n_1344),
.B(n_1376),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1644),
.A2(n_1400),
.B(n_1345),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1589),
.B(n_1407),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1537),
.B(n_1356),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1578),
.B(n_1705),
.Y(n_1735)
);

BUFx4f_ASAP7_75t_L g1736 ( 
.A(n_1634),
.Y(n_1736)
);

AOI22x1_ASAP7_75t_L g1737 ( 
.A1(n_1706),
.A2(n_1517),
.B1(n_1400),
.B2(n_1515),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1695),
.A2(n_1501),
.B(n_1429),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1641),
.A2(n_1400),
.B(n_1505),
.Y(n_1739)
);

NAND2xp33_ASAP7_75t_L g1740 ( 
.A(n_1634),
.B(n_1400),
.Y(n_1740)
);

NOR2xp67_ASAP7_75t_L g1741 ( 
.A(n_1560),
.B(n_1501),
.Y(n_1741)
);

AO31x2_ASAP7_75t_L g1742 ( 
.A1(n_1678),
.A2(n_1507),
.A3(n_1399),
.B(n_109),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1544),
.B(n_104),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1663),
.A2(n_111),
.B1(n_108),
.B2(n_110),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1685),
.A2(n_108),
.B(n_110),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1526),
.A2(n_279),
.B(n_278),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1541),
.B(n_280),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1526),
.A2(n_284),
.B(n_283),
.Y(n_1748)
);

AND2x2_ASAP7_75t_SL g1749 ( 
.A(n_1567),
.B(n_1617),
.Y(n_1749)
);

AO21x1_ASAP7_75t_L g1750 ( 
.A1(n_1529),
.A2(n_111),
.B(n_112),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_SL g1751 ( 
.A1(n_1559),
.A2(n_112),
.B(n_113),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1623),
.B(n_1681),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1528),
.A2(n_1689),
.B(n_1681),
.Y(n_1753)
);

AO32x2_ASAP7_75t_L g1754 ( 
.A1(n_1530),
.A2(n_115),
.A3(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1528),
.A2(n_287),
.B(n_285),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1712),
.B(n_115),
.Y(n_1756)
);

AOI21xp33_ASAP7_75t_L g1757 ( 
.A1(n_1686),
.A2(n_116),
.B(n_117),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1541),
.B(n_288),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1684),
.B(n_118),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1659),
.B(n_118),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1543),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1634),
.Y(n_1762)
);

BUFx4f_ASAP7_75t_SL g1763 ( 
.A(n_1698),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1569),
.B(n_289),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1604),
.A2(n_291),
.B(n_290),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1562),
.Y(n_1766)
);

OAI21x1_ASAP7_75t_L g1767 ( 
.A1(n_1636),
.A2(n_1576),
.B(n_1573),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1603),
.A2(n_294),
.B(n_293),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1633),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_1769)
);

NAND2x1_ASAP7_75t_L g1770 ( 
.A(n_1574),
.B(n_298),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1601),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1545),
.A2(n_300),
.B(n_299),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1621),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1581),
.A2(n_304),
.B(n_301),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1535),
.B(n_119),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1565),
.Y(n_1776)
);

AOI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1594),
.A2(n_307),
.B(n_305),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1527),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1680),
.B(n_120),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1587),
.B(n_121),
.Y(n_1780)
);

AOI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1549),
.A2(n_309),
.B(n_308),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1579),
.B(n_122),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1625),
.B(n_312),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1539),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1622),
.B(n_123),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1618),
.B(n_123),
.Y(n_1786)
);

AO31x2_ASAP7_75t_L g1787 ( 
.A1(n_1597),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1542),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1703),
.A2(n_125),
.B(n_126),
.Y(n_1789)
);

NOR2x1_ASAP7_75t_SL g1790 ( 
.A(n_1697),
.B(n_316),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1677),
.B(n_127),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1600),
.B(n_128),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1697),
.A2(n_517),
.B(n_321),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1626),
.A2(n_516),
.B(n_322),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1540),
.Y(n_1795)
);

OAI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1556),
.A2(n_1564),
.B(n_1558),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1699),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1554),
.A2(n_132),
.B(n_129),
.C(n_131),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1660),
.A2(n_136),
.B1(n_132),
.B2(n_133),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1607),
.B(n_137),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1608),
.A2(n_515),
.B(n_323),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1637),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1683),
.A2(n_514),
.B(n_326),
.Y(n_1803)
);

INVxp67_ASAP7_75t_SL g1804 ( 
.A(n_1575),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1557),
.A2(n_139),
.B(n_140),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1635),
.B(n_140),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1638),
.B(n_141),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1653),
.B(n_320),
.Y(n_1808)
);

NOR2xp67_ASAP7_75t_SL g1809 ( 
.A(n_1710),
.B(n_141),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1670),
.B(n_142),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1612),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_SL g1812 ( 
.A1(n_1650),
.A2(n_142),
.B(n_143),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1596),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1652),
.B(n_143),
.Y(n_1814)
);

NAND2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1574),
.B(n_1584),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1645),
.A2(n_329),
.B(n_328),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1683),
.A2(n_513),
.B(n_335),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1586),
.A2(n_144),
.B(n_146),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1669),
.A2(n_512),
.B(n_336),
.Y(n_1819)
);

OAI21x1_ASAP7_75t_SL g1820 ( 
.A1(n_1593),
.A2(n_144),
.B(n_146),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1688),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1821)
);

NAND2x1_ASAP7_75t_L g1822 ( 
.A(n_1584),
.B(n_1613),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1591),
.A2(n_150),
.B(n_147),
.C(n_149),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1651),
.A2(n_337),
.B(n_332),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1585),
.B(n_150),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1629),
.B(n_1640),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1566),
.B(n_151),
.Y(n_1827)
);

INVx3_ASAP7_75t_SL g1828 ( 
.A(n_1605),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1631),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1653),
.B(n_338),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1568),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1570),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_SL g1833 ( 
.A1(n_1577),
.A2(n_151),
.B(n_152),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1647),
.A2(n_341),
.B(n_339),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1646),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1668),
.B(n_153),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1666),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1619),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1667),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1674),
.A2(n_155),
.B(n_156),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1668),
.B(n_157),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1665),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1842)
);

AOI21x1_ASAP7_75t_SL g1843 ( 
.A1(n_1571),
.A2(n_158),
.B(n_159),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1643),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1666),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1590),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1656),
.A2(n_347),
.B(n_343),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1657),
.A2(n_350),
.B(n_348),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1598),
.A2(n_354),
.B(n_353),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1580),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_SL g1851 ( 
.A1(n_1711),
.A2(n_163),
.B(n_164),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1524),
.A2(n_1561),
.B(n_1624),
.Y(n_1852)
);

OAI21x1_ASAP7_75t_SL g1853 ( 
.A1(n_1690),
.A2(n_164),
.B(n_165),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1602),
.A2(n_356),
.B(n_355),
.Y(n_1854)
);

O2A1O1Ixp5_ASAP7_75t_L g1855 ( 
.A1(n_1534),
.A2(n_169),
.B(n_166),
.C(n_167),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1675),
.A2(n_166),
.B(n_169),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1671),
.B(n_170),
.Y(n_1857)
);

AOI22x1_ASAP7_75t_L g1858 ( 
.A1(n_1592),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1858)
);

AO21x1_ASAP7_75t_L g1859 ( 
.A1(n_1538),
.A2(n_171),
.B(n_172),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1654),
.B(n_173),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1606),
.A2(n_363),
.B(n_361),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1627),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1570),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1671),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1682),
.A2(n_178),
.B1(n_175),
.B2(n_176),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1694),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1651),
.A2(n_511),
.B(n_365),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1609),
.A2(n_366),
.B(n_364),
.Y(n_1868)
);

AO31x2_ASAP7_75t_L g1869 ( 
.A1(n_1649),
.A2(n_180),
.A3(n_178),
.B(n_179),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1639),
.B(n_367),
.Y(n_1870)
);

AOI221x1_ASAP7_75t_L g1871 ( 
.A1(n_1628),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.C(n_183),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1548),
.A2(n_185),
.B(n_181),
.C(n_183),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1692),
.B(n_186),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_L g1874 ( 
.A1(n_1662),
.A2(n_369),
.B(n_368),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1679),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1630),
.A2(n_371),
.B(n_370),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1729),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1735),
.B(n_1658),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1721),
.A2(n_1648),
.B(n_1623),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1725),
.B(n_1661),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1804),
.B(n_1676),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1749),
.A2(n_1547),
.B1(n_1552),
.B2(n_1620),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1805),
.B(n_1555),
.C(n_1614),
.Y(n_1883)
);

AND2x2_ASAP7_75t_SL g1884 ( 
.A(n_1740),
.B(n_1648),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1764),
.A2(n_1709),
.B1(n_1588),
.B2(n_1555),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1723),
.A2(n_1614),
.B(n_1610),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1727),
.B(n_1813),
.Y(n_1887)
);

CKINVDCx11_ASAP7_75t_R g1888 ( 
.A(n_1828),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1839),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1734),
.B(n_1693),
.Y(n_1890)
);

NOR2xp67_ASAP7_75t_SL g1891 ( 
.A(n_1726),
.B(n_1666),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_SL g1892 ( 
.A(n_1872),
.B(n_1655),
.C(n_1704),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1736),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1844),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1840),
.A2(n_1553),
.B(n_1696),
.C(n_1702),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1778),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1785),
.B(n_1701),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1733),
.A2(n_1613),
.B1(n_1642),
.B2(n_1696),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1766),
.B(n_1551),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1757),
.A2(n_1691),
.B1(n_1673),
.B2(n_1551),
.C(n_1616),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1752),
.B(n_1610),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_SL g1902 ( 
.A1(n_1798),
.A2(n_1615),
.B(n_1610),
.C(n_1642),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1739),
.A2(n_1691),
.B(n_1673),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1863),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1736),
.Y(n_1905)
);

CKINVDCx8_ASAP7_75t_R g1906 ( 
.A(n_1762),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1760),
.B(n_1551),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1773),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1732),
.A2(n_1691),
.B(n_1673),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1775),
.B(n_1615),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1808),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1716),
.B(n_1615),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1796),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1810),
.B(n_1563),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1762),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1795),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1730),
.B(n_1615),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1866),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1870),
.A2(n_1783),
.B1(n_1752),
.B2(n_1809),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1767),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1860),
.B(n_1563),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1808),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1771),
.Y(n_1923)
);

BUFx12f_ASAP7_75t_L g1924 ( 
.A(n_1832),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1811),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1829),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1864),
.B(n_1563),
.Y(n_1927)
);

OR2x6_ASAP7_75t_L g1928 ( 
.A(n_1753),
.B(n_1616),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1761),
.B(n_1572),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1776),
.B(n_1572),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1858),
.A2(n_1818),
.B1(n_1789),
.B2(n_1859),
.Y(n_1931)
);

NAND2x1p5_ASAP7_75t_L g1932 ( 
.A(n_1762),
.B(n_1572),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1718),
.B(n_1595),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1830),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1728),
.B(n_1595),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1784),
.Y(n_1936)
);

OA22x2_ASAP7_75t_L g1937 ( 
.A1(n_1799),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1875),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1772),
.A2(n_1616),
.B(n_1595),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1837),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1830),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1792),
.B(n_1800),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_L g1943 ( 
.A(n_1823),
.B(n_187),
.C(n_189),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1806),
.B(n_189),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1788),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1717),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1837),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1763),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1852),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1869),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1831),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1837),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1845),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1845),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1869),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1869),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1718),
.B(n_372),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1845),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1827),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1815),
.Y(n_1960)
);

INVx5_ASAP7_75t_L g1961 ( 
.A(n_1790),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1787),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1807),
.B(n_194),
.Y(n_1963)
);

CKINVDCx16_ASAP7_75t_R g1964 ( 
.A(n_1826),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1814),
.B(n_195),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1822),
.Y(n_1966)
);

O2A1O1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1846),
.A2(n_195),
.B(n_196),
.C(n_197),
.Y(n_1967)
);

O2A1O1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1850),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1741),
.B(n_373),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1786),
.B(n_374),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1720),
.A2(n_376),
.B(n_375),
.Y(n_1971)
);

O2A1O1Ixp33_ASAP7_75t_SL g1972 ( 
.A1(n_1802),
.A2(n_199),
.B(n_200),
.C(n_201),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1780),
.B(n_381),
.Y(n_1973)
);

BUFx12f_ASAP7_75t_L g1974 ( 
.A(n_1747),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1865),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1836),
.Y(n_1976)
);

NAND3xp33_ASAP7_75t_L g1977 ( 
.A(n_1769),
.B(n_203),
.C(n_204),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1838),
.A2(n_1745),
.B1(n_1856),
.B2(n_1750),
.Y(n_1978)
);

BUFx2_ASAP7_75t_L g1979 ( 
.A(n_1841),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1758),
.B(n_382),
.Y(n_1980)
);

AOI21x1_ASAP7_75t_SL g1981 ( 
.A1(n_1910),
.A2(n_1782),
.B(n_1779),
.Y(n_1981)
);

AOI21x1_ASAP7_75t_SL g1982 ( 
.A1(n_1944),
.A2(n_1791),
.B(n_1756),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1962),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1938),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1914),
.B(n_1907),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1923),
.B(n_1959),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1950),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_SL g1988 ( 
.A1(n_1895),
.A2(n_1790),
.B(n_1871),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1896),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1936),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1919),
.B(n_1743),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1921),
.B(n_1979),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1897),
.B(n_1787),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1936),
.Y(n_1994)
);

INVx4_ASAP7_75t_L g1995 ( 
.A(n_1974),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1945),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1964),
.B(n_1787),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1918),
.B(n_1722),
.Y(n_1998)
);

OR2x6_ASAP7_75t_SL g1999 ( 
.A(n_1904),
.B(n_1744),
.Y(n_1999)
);

NOR2xp67_ASAP7_75t_L g2000 ( 
.A(n_1889),
.B(n_1774),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_SL g2001 ( 
.A1(n_1891),
.A2(n_1793),
.B(n_1835),
.C(n_1794),
.Y(n_2001)
);

INVx4_ASAP7_75t_L g2002 ( 
.A(n_1901),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1883),
.A2(n_1855),
.B(n_1867),
.C(n_1824),
.Y(n_2003)
);

NOR2xp67_ASAP7_75t_L g2004 ( 
.A(n_1926),
.B(n_1801),
.Y(n_2004)
);

AND2x2_ASAP7_75t_SL g2005 ( 
.A(n_1884),
.B(n_1931),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1879),
.A2(n_1886),
.B(n_1902),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1887),
.B(n_1759),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1968),
.A2(n_1719),
.B(n_1854),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1951),
.B(n_1857),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1976),
.B(n_1873),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1950),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1980),
.A2(n_1731),
.B(n_1738),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1945),
.B(n_1825),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1966),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1920),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1901),
.B(n_1724),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1913),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1878),
.B(n_1821),
.Y(n_2018)
);

A2O1A1Ixp33_ASAP7_75t_SL g2019 ( 
.A1(n_1967),
.A2(n_1819),
.B(n_1803),
.C(n_1817),
.Y(n_2019)
);

OR2x6_ASAP7_75t_SL g2020 ( 
.A(n_1948),
.B(n_1882),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1955),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1956),
.Y(n_2022)
);

A2O1A1Ixp33_ASAP7_75t_L g2023 ( 
.A1(n_1943),
.A2(n_1876),
.B(n_1797),
.C(n_1862),
.Y(n_2023)
);

A2O1A1Ixp33_ASAP7_75t_SL g2024 ( 
.A1(n_1978),
.A2(n_1949),
.B(n_1890),
.C(n_1939),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1877),
.Y(n_2025)
);

INVx2_ASAP7_75t_SL g2026 ( 
.A(n_1908),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1916),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1928),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1894),
.B(n_1768),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1942),
.B(n_1714),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1888),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1881),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1880),
.B(n_1751),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1924),
.Y(n_2034)
);

INVxp67_ASAP7_75t_SL g2035 ( 
.A(n_1935),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1954),
.B(n_1754),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1925),
.B(n_1742),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1912),
.B(n_1742),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1892),
.B(n_1777),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1885),
.A2(n_1977),
.B1(n_1937),
.B2(n_1975),
.Y(n_2040)
);

INVxp33_ASAP7_75t_L g2041 ( 
.A(n_1992),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1996),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1983),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_2005),
.B(n_1961),
.Y(n_2045)
);

NOR2x1_ASAP7_75t_R g2046 ( 
.A(n_2031),
.B(n_1961),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1990),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_2016),
.Y(n_2048)
);

AOI21x1_ASAP7_75t_L g2049 ( 
.A1(n_2006),
.A2(n_1971),
.B(n_1903),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1994),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_2017),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1987),
.Y(n_2052)
);

OA21x2_ASAP7_75t_L g2053 ( 
.A1(n_2021),
.A2(n_1909),
.B(n_1765),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1993),
.B(n_1961),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1987),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1997),
.B(n_1754),
.Y(n_2056)
);

AOI21x1_ASAP7_75t_L g2057 ( 
.A1(n_2012),
.A2(n_1781),
.B(n_1946),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2011),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2011),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2015),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2022),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1983),
.Y(n_2062)
);

OA21x2_ASAP7_75t_L g2063 ( 
.A1(n_2039),
.A2(n_1715),
.B(n_1816),
.Y(n_2063)
);

OA21x2_ASAP7_75t_L g2064 ( 
.A1(n_2039),
.A2(n_1847),
.B(n_1834),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2035),
.B(n_1917),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_2037),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_2030),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2035),
.Y(n_2068)
);

INVx2_ASAP7_75t_SL g2069 ( 
.A(n_2016),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2015),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2005),
.A2(n_1833),
.B1(n_1820),
.B2(n_1812),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1989),
.B(n_1927),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1984),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2028),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2040),
.A2(n_1999),
.B1(n_1991),
.B2(n_2020),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2022),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2042),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2047),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2067),
.B(n_2065),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2042),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2062),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2075),
.A2(n_2023),
.B1(n_1988),
.B2(n_1991),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2047),
.Y(n_2083)
);

INVx5_ASAP7_75t_L g2084 ( 
.A(n_2076),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2041),
.B(n_2032),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2068),
.B(n_2038),
.Y(n_2086)
);

NOR2xp67_ASAP7_75t_R g2087 ( 
.A(n_2046),
.B(n_1995),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_2062),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2050),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2048),
.B(n_2036),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2050),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2042),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2043),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2066),
.B(n_1986),
.Y(n_2094)
);

AND2x4_ASAP7_75t_SL g2095 ( 
.A(n_2054),
.B(n_2014),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_2075),
.A2(n_2018),
.B1(n_1842),
.B2(n_2033),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2043),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2043),
.Y(n_2098)
);

OR2x6_ASAP7_75t_L g2099 ( 
.A(n_2082),
.B(n_2008),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2077),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2078),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2077),
.Y(n_2102)
);

AOI222xp33_ASAP7_75t_L g2103 ( 
.A1(n_2096),
.A2(n_2024),
.B1(n_1963),
.B2(n_1965),
.C1(n_2056),
.C2(n_2023),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2090),
.B(n_2048),
.Y(n_2104)
);

OA21x2_ASAP7_75t_L g2105 ( 
.A1(n_2080),
.A2(n_2044),
.B(n_2076),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2086),
.Y(n_2106)
);

AOI21xp33_ASAP7_75t_L g2107 ( 
.A1(n_2096),
.A2(n_2024),
.B(n_2067),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2101),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_2106),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2105),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2104),
.B(n_2079),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2100),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2104),
.B(n_2095),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2109),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2111),
.B(n_2108),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2113),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2112),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2113),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2110),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2110),
.B(n_2095),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_2109),
.Y(n_2121)
);

NAND2x1_ASAP7_75t_L g2122 ( 
.A(n_2109),
.B(n_2105),
.Y(n_2122)
);

NAND3xp33_ASAP7_75t_L g2123 ( 
.A(n_2109),
.B(n_2103),
.C(n_2107),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2117),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_2121),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2114),
.B(n_2099),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2123),
.B(n_1985),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2116),
.B(n_1995),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2117),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2115),
.B(n_2099),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_2118),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_2120),
.B(n_2099),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2119),
.B(n_2085),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2119),
.Y(n_2134)
);

NOR2xp67_ASAP7_75t_L g2135 ( 
.A(n_2125),
.B(n_2084),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_2131),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2134),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2124),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2128),
.A2(n_2045),
.B1(n_2122),
.B2(n_2004),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2129),
.Y(n_2140)
);

AOI32xp33_ASAP7_75t_L g2141 ( 
.A1(n_2127),
.A2(n_2056),
.A3(n_2071),
.B1(n_2054),
.B2(n_2090),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2132),
.B(n_2034),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2136),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2138),
.B(n_2126),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2142),
.B(n_2132),
.Y(n_2145)
);

NAND2x1p5_ASAP7_75t_L g2146 ( 
.A(n_2135),
.B(n_2130),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2146),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_SL g2148 ( 
.A(n_2143),
.B(n_2144),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2145),
.A2(n_2141),
.B1(n_2139),
.B2(n_2133),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2143),
.Y(n_2150)
);

NOR2xp67_ASAP7_75t_L g2151 ( 
.A(n_2147),
.B(n_2150),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2149),
.A2(n_2140),
.B1(n_2137),
.B2(n_2084),
.Y(n_2152)
);

NAND2x1p5_ASAP7_75t_L g2153 ( 
.A(n_2148),
.B(n_1969),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2150),
.B(n_2094),
.Y(n_2154)
);

OAI31xp33_ASAP7_75t_L g2155 ( 
.A1(n_2148),
.A2(n_1972),
.A3(n_2019),
.B(n_2003),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_2151),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2152),
.A2(n_2026),
.B(n_2000),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2154),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_L g2159 ( 
.A(n_2153),
.B(n_2087),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2155),
.B(n_2100),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2153),
.B(n_2102),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2154),
.B(n_2102),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_2153),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_2074),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_2153),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_2163),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2158),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2156),
.B(n_2165),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_2165),
.B(n_1973),
.C(n_1970),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2160),
.B(n_2081),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2164),
.B(n_2161),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2162),
.B(n_2081),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_R g2173 ( 
.A(n_2159),
.B(n_204),
.Y(n_2173)
);

CKINVDCx14_ASAP7_75t_R g2174 ( 
.A(n_2157),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_2156),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2165),
.A2(n_2084),
.B1(n_2105),
.B2(n_2088),
.Y(n_2176)
);

AOI211xp5_ASAP7_75t_SL g2177 ( 
.A1(n_2156),
.A2(n_1969),
.B(n_1957),
.C(n_1899),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2158),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2168),
.Y(n_2179)
);

NOR2x1_ASAP7_75t_L g2180 ( 
.A(n_2167),
.B(n_205),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2166),
.B(n_2084),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2175),
.B(n_2178),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2171),
.B(n_2088),
.Y(n_2183)
);

AOI211x1_ASAP7_75t_L g2184 ( 
.A1(n_2170),
.A2(n_2010),
.B(n_1898),
.C(n_2007),
.Y(n_2184)
);

NOR2x1_ASAP7_75t_L g2185 ( 
.A(n_2169),
.B(n_206),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2172),
.Y(n_2186)
);

NAND4xp25_ASAP7_75t_L g2187 ( 
.A(n_2177),
.B(n_1900),
.C(n_2019),
.D(n_2001),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2173),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2174),
.A2(n_2046),
.B(n_1853),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2176),
.Y(n_2190)
);

NAND3xp33_ASAP7_75t_SL g2191 ( 
.A(n_2173),
.B(n_1906),
.C(n_1770),
.Y(n_2191)
);

NAND4xp25_ASAP7_75t_L g2192 ( 
.A(n_2182),
.B(n_2002),
.C(n_2014),
.D(n_2001),
.Y(n_2192)
);

O2A1O1Ixp33_ASAP7_75t_L g2193 ( 
.A1(n_2190),
.A2(n_1851),
.B(n_1905),
.C(n_1893),
.Y(n_2193)
);

NAND4xp25_ASAP7_75t_SL g2194 ( 
.A(n_2189),
.B(n_2003),
.C(n_2013),
.D(n_2029),
.Y(n_2194)
);

NAND3xp33_ASAP7_75t_L g2195 ( 
.A(n_2180),
.B(n_206),
.C(n_207),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2188),
.B(n_2083),
.Y(n_2196)
);

NOR2x1_ASAP7_75t_L g2197 ( 
.A(n_2179),
.B(n_207),
.Y(n_2197)
);

NOR2x1_ASAP7_75t_SL g2198 ( 
.A(n_2191),
.B(n_1915),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2185),
.B(n_2048),
.Y(n_2199)
);

NOR5xp2_ASAP7_75t_L g2200 ( 
.A(n_2186),
.B(n_208),
.C(n_209),
.D(n_210),
.E(n_211),
.Y(n_2200)
);

OAI211xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2183),
.A2(n_213),
.B(n_209),
.C(n_212),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2181),
.Y(n_2202)
);

NOR3x1_ASAP7_75t_L g2203 ( 
.A(n_2187),
.B(n_1952),
.C(n_212),
.Y(n_2203)
);

AOI211xp5_ASAP7_75t_L g2204 ( 
.A1(n_2201),
.A2(n_2184),
.B(n_216),
.C(n_214),
.Y(n_2204)
);

AOI211xp5_ASAP7_75t_L g2205 ( 
.A1(n_2202),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2205)
);

NAND4xp75_ASAP7_75t_L g2206 ( 
.A(n_2197),
.B(n_218),
.C(n_215),
.D(n_217),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_2195),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2193),
.A2(n_1930),
.B(n_1929),
.Y(n_2208)
);

NOR2x1_ASAP7_75t_L g2209 ( 
.A(n_2199),
.B(n_217),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2203),
.B(n_219),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2198),
.B(n_2196),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2192),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2194),
.Y(n_2213)
);

NAND3xp33_ASAP7_75t_L g2214 ( 
.A(n_2200),
.B(n_219),
.C(n_220),
.Y(n_2214)
);

NAND2x1p5_ASAP7_75t_L g2215 ( 
.A(n_2197),
.B(n_1947),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2197),
.B(n_1958),
.Y(n_2216)
);

OAI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2195),
.A2(n_1748),
.B(n_1746),
.Y(n_2217)
);

NOR3xp33_ASAP7_75t_L g2218 ( 
.A(n_2195),
.B(n_220),
.C(n_221),
.Y(n_2218)
);

NOR3xp33_ASAP7_75t_L g2219 ( 
.A(n_2195),
.B(n_222),
.C(n_224),
.Y(n_2219)
);

NAND4xp75_ASAP7_75t_L g2220 ( 
.A(n_2209),
.B(n_2210),
.C(n_2211),
.D(n_2212),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2216),
.B(n_2205),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2216),
.B(n_222),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2214),
.A2(n_1953),
.B1(n_1940),
.B2(n_1915),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2206),
.B(n_225),
.Y(n_2224)
);

NOR2x1_ASAP7_75t_L g2225 ( 
.A(n_2213),
.B(n_225),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2215),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2218),
.B(n_226),
.Y(n_2227)
);

INVxp33_ASAP7_75t_SL g2228 ( 
.A(n_2219),
.Y(n_2228)
);

XOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2207),
.B(n_227),
.Y(n_2229)
);

NOR4xp25_ASAP7_75t_L g2230 ( 
.A(n_2204),
.B(n_229),
.C(n_227),
.D(n_228),
.Y(n_2230)
);

NOR3xp33_ASAP7_75t_L g2231 ( 
.A(n_2208),
.B(n_228),
.C(n_229),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2217),
.B(n_230),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2215),
.B(n_230),
.Y(n_2233)
);

NOR3x1_ASAP7_75t_L g2234 ( 
.A(n_2214),
.B(n_231),
.C(n_232),
.Y(n_2234)
);

NAND3xp33_ASAP7_75t_L g2235 ( 
.A(n_2209),
.B(n_232),
.C(n_1915),
.Y(n_2235)
);

OA21x2_ASAP7_75t_L g2236 ( 
.A1(n_2210),
.A2(n_1755),
.B(n_1848),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2207),
.B(n_1953),
.C(n_2002),
.Y(n_2237)
);

NOR2x1_ASAP7_75t_L g2238 ( 
.A(n_2206),
.B(n_1940),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2209),
.Y(n_2239)
);

NOR2x1_ASAP7_75t_L g2240 ( 
.A(n_2206),
.B(n_1940),
.Y(n_2240)
);

NAND4xp75_ASAP7_75t_L g2241 ( 
.A(n_2209),
.B(n_1854),
.C(n_2009),
.D(n_2065),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2209),
.Y(n_2242)
);

NOR2xp67_ASAP7_75t_L g2243 ( 
.A(n_2214),
.B(n_383),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2216),
.B(n_2089),
.Y(n_2244)
);

NAND4xp75_ASAP7_75t_L g2245 ( 
.A(n_2209),
.B(n_1982),
.C(n_2091),
.D(n_2061),
.Y(n_2245)
);

AOI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2230),
.A2(n_2098),
.B1(n_2097),
.B2(n_2093),
.C(n_2092),
.Y(n_2246)
);

NAND2x1p5_ASAP7_75t_L g2247 ( 
.A(n_2239),
.B(n_1960),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2234),
.B(n_2069),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2224),
.B(n_2028),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2243),
.A2(n_2044),
.B1(n_1932),
.B2(n_1960),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_2221),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2229),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2222),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2238),
.B(n_2069),
.Y(n_2254)
);

NOR2xp67_ASAP7_75t_L g2255 ( 
.A(n_2235),
.B(n_384),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2242),
.B(n_2080),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_SL g2257 ( 
.A1(n_2233),
.A2(n_1933),
.B(n_1927),
.C(n_1843),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2225),
.B(n_1933),
.Y(n_2258)
);

NAND4xp75_ASAP7_75t_L g2259 ( 
.A(n_2226),
.B(n_385),
.C(n_386),
.D(n_387),
.Y(n_2259)
);

XNOR2xp5_ASAP7_75t_L g2260 ( 
.A(n_2220),
.B(n_388),
.Y(n_2260)
);

OAI211xp5_ASAP7_75t_SL g2261 ( 
.A1(n_2232),
.A2(n_1981),
.B(n_390),
.C(n_391),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2228),
.B(n_389),
.Y(n_2262)
);

NAND4xp75_ASAP7_75t_L g2263 ( 
.A(n_2240),
.B(n_392),
.C(n_393),
.D(n_394),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2231),
.B(n_2061),
.C(n_2063),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2237),
.B(n_2027),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2252),
.B(n_2227),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2248),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2255),
.B(n_2244),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2254),
.B(n_2223),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2258),
.B(n_2245),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2259),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2263),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_2247),
.Y(n_2273)
);

XNOR2xp5_ASAP7_75t_L g2274 ( 
.A(n_2260),
.B(n_2251),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2250),
.B(n_2241),
.Y(n_2275)
);

NOR2x1_ASAP7_75t_L g2276 ( 
.A(n_2262),
.B(n_2236),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2249),
.B(n_2236),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_2256),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2253),
.B(n_2063),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2261),
.A2(n_2069),
.B1(n_2058),
.B2(n_2059),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2265),
.B(n_2063),
.Y(n_2281)
);

XNOR2x1_ASAP7_75t_L g2282 ( 
.A(n_2264),
.B(n_395),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2257),
.Y(n_2283)
);

XOR2x1_ASAP7_75t_L g2284 ( 
.A(n_2246),
.B(n_397),
.Y(n_2284)
);

XOR2xp5_ASAP7_75t_L g2285 ( 
.A(n_2251),
.B(n_398),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2259),
.Y(n_2286)
);

HB1xp67_ASAP7_75t_L g2287 ( 
.A(n_2252),
.Y(n_2287)
);

NAND2x1_ASAP7_75t_SL g2288 ( 
.A(n_2273),
.B(n_2287),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2267),
.B(n_400),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2274),
.A2(n_2052),
.B1(n_2055),
.B2(n_2058),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2268),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2272),
.B(n_2072),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_SL g2293 ( 
.A1(n_2285),
.A2(n_401),
.B(n_402),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2271),
.B(n_2072),
.Y(n_2294)
);

NAND2x1p5_ASAP7_75t_L g2295 ( 
.A(n_2286),
.B(n_2278),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2284),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2280),
.A2(n_2052),
.B1(n_2055),
.B2(n_2059),
.Y(n_2297)
);

AOI21xp33_ASAP7_75t_SL g2298 ( 
.A1(n_2274),
.A2(n_404),
.B(n_406),
.Y(n_2298)
);

AOI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_2270),
.A2(n_407),
.B(n_409),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2282),
.Y(n_2300)
);

OAI22x1_ASAP7_75t_L g2301 ( 
.A1(n_2283),
.A2(n_2057),
.B1(n_2049),
.B2(n_1737),
.Y(n_2301)
);

NAND2x1_ASAP7_75t_SL g2302 ( 
.A(n_2276),
.B(n_2277),
.Y(n_2302)
);

AO22x2_ASAP7_75t_L g2303 ( 
.A1(n_2266),
.A2(n_2076),
.B1(n_414),
.B2(n_415),
.Y(n_2303)
);

XOR2xp5_ASAP7_75t_L g2304 ( 
.A(n_2269),
.B(n_411),
.Y(n_2304)
);

NAND4xp75_ASAP7_75t_L g2305 ( 
.A(n_2275),
.B(n_418),
.C(n_419),
.D(n_421),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2279),
.B(n_422),
.Y(n_2306)
);

A2O1A1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2288),
.A2(n_2281),
.B(n_1849),
.C(n_1868),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2302),
.Y(n_2308)
);

AND3x2_ASAP7_75t_L g2309 ( 
.A(n_2296),
.B(n_423),
.C(n_424),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2303),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2292),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2294),
.B(n_425),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2291),
.B(n_426),
.C(n_428),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2295),
.Y(n_2314)
);

AOI211xp5_ASAP7_75t_L g2315 ( 
.A1(n_2293),
.A2(n_429),
.B(n_431),
.C(n_433),
.Y(n_2315)
);

OAI21xp33_ASAP7_75t_L g2316 ( 
.A1(n_2300),
.A2(n_2049),
.B(n_1998),
.Y(n_2316)
);

AOI221x1_ASAP7_75t_L g2317 ( 
.A1(n_2289),
.A2(n_2306),
.B1(n_2303),
.B2(n_2298),
.C(n_2299),
.Y(n_2317)
);

OAI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2290),
.A2(n_2057),
.B1(n_2064),
.B2(n_1911),
.C(n_1941),
.Y(n_2318)
);

NAND4xp25_ASAP7_75t_L g2319 ( 
.A(n_2297),
.B(n_434),
.C(n_435),
.D(n_437),
.Y(n_2319)
);

OAI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2305),
.A2(n_1861),
.B(n_1874),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_SL g2321 ( 
.A1(n_2304),
.A2(n_1941),
.B1(n_1922),
.B2(n_1934),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2301),
.A2(n_2073),
.B1(n_1911),
.B2(n_1922),
.Y(n_2322)
);

AOI221xp5_ASAP7_75t_L g2323 ( 
.A1(n_2303),
.A2(n_2073),
.B1(n_1998),
.B2(n_2025),
.C(n_2051),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2288),
.B(n_438),
.Y(n_2324)
);

NAND3xp33_ASAP7_75t_SL g2325 ( 
.A(n_2308),
.B(n_440),
.C(n_442),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_L g2326 ( 
.A(n_2314),
.B(n_443),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_SL g2327 ( 
.A1(n_2310),
.A2(n_1934),
.B1(n_2064),
.B2(n_2063),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2324),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2311),
.Y(n_2329)
);

OAI322xp33_ASAP7_75t_L g2330 ( 
.A1(n_2312),
.A2(n_444),
.A3(n_446),
.B1(n_448),
.B2(n_450),
.C1(n_451),
.C2(n_452),
.Y(n_2330)
);

NOR3xp33_ASAP7_75t_L g2331 ( 
.A(n_2315),
.B(n_2319),
.C(n_2313),
.Y(n_2331)
);

NAND4xp25_ASAP7_75t_L g2332 ( 
.A(n_2317),
.B(n_2309),
.C(n_2322),
.D(n_2307),
.Y(n_2332)
);

NAND4xp25_ASAP7_75t_L g2333 ( 
.A(n_2320),
.B(n_453),
.C(n_455),
.D(n_458),
.Y(n_2333)
);

NAND4xp25_ASAP7_75t_L g2334 ( 
.A(n_2318),
.B(n_2316),
.C(n_2323),
.D(n_2321),
.Y(n_2334)
);

NOR2x1p5_ASAP7_75t_L g2335 ( 
.A(n_2324),
.B(n_459),
.Y(n_2335)
);

AO21x2_ASAP7_75t_L g2336 ( 
.A1(n_2329),
.A2(n_460),
.B(n_461),
.Y(n_2336)
);

OA21x2_ASAP7_75t_L g2337 ( 
.A1(n_2328),
.A2(n_462),
.B(n_463),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2326),
.Y(n_2338)
);

AOI221x1_ASAP7_75t_L g2339 ( 
.A1(n_2332),
.A2(n_464),
.B1(n_465),
.B2(n_467),
.C(n_468),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2331),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2333),
.A2(n_2073),
.B1(n_2064),
.B2(n_2070),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2334),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2325),
.A2(n_2064),
.B1(n_2070),
.B2(n_2060),
.Y(n_2343)
);

OAI22xp33_ASAP7_75t_SL g2344 ( 
.A1(n_2330),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2327),
.B(n_473),
.Y(n_2345)
);

NAND4xp75_ASAP7_75t_L g2346 ( 
.A(n_2329),
.B(n_474),
.C(n_476),
.D(n_478),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2335),
.B(n_479),
.Y(n_2347)
);

AO22x2_ASAP7_75t_L g2348 ( 
.A1(n_2338),
.A2(n_481),
.B1(n_482),
.B2(n_483),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2344),
.B(n_2342),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2340),
.B(n_484),
.C(n_486),
.Y(n_2350)
);

XNOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2347),
.B(n_487),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2345),
.A2(n_2053),
.B1(n_2060),
.B2(n_2070),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_2336),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2337),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2339),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2353),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2351),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2354),
.Y(n_2358)
);

AOI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2358),
.A2(n_2349),
.B(n_2355),
.Y(n_2359)
);

NAND3xp33_ASAP7_75t_L g2360 ( 
.A(n_2356),
.B(n_2350),
.C(n_2341),
.Y(n_2360)
);

NAND2xp33_ASAP7_75t_SL g2361 ( 
.A(n_2359),
.B(n_2357),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2361),
.Y(n_2362)
);

BUFx2_ASAP7_75t_L g2363 ( 
.A(n_2361),
.Y(n_2363)
);

AND2x2_ASAP7_75t_SL g2364 ( 
.A(n_2363),
.B(n_2360),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2362),
.B(n_2343),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2364),
.A2(n_2348),
.B(n_2352),
.Y(n_2366)
);

AOI211xp5_ASAP7_75t_L g2367 ( 
.A1(n_2366),
.A2(n_2365),
.B(n_2346),
.C(n_2348),
.Y(n_2367)
);


endmodule