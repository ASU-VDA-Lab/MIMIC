module fake_jpeg_4922_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_31),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_21),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.C(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_50),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_66),
.B1(n_69),
.B2(n_17),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_29),
.B1(n_19),
.B2(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_56),
.B1(n_59),
.B2(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_62),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_62),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_19),
.B2(n_3),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_61),
.Y(n_93)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_14),
.B1(n_27),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_34),
.Y(n_72)
);

OAI22x1_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_29),
.B1(n_19),
.B2(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_32),
.A2(n_23),
.B1(n_17),
.B2(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_87),
.B1(n_59),
.B2(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_88),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_44),
.B1(n_42),
.B2(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_47),
.B1(n_59),
.B2(n_46),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_100),
.B1(n_107),
.B2(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_59),
.B1(n_70),
.B2(n_71),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_108),
.C(n_80),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_79),
.B(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_68),
.B1(n_65),
.B2(n_47),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_51),
.C(n_61),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_57),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_51),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_96),
.B(n_79),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_101),
.B(n_113),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_87),
.B1(n_77),
.B2(n_94),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_119),
.B(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_83),
.B1(n_81),
.B2(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_83),
.B1(n_95),
.B2(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_89),
.B1(n_57),
.B2(n_49),
.Y(n_127)
);

OR2x6_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_49),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_106),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_108),
.C(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_137),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_138),
.B(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_106),
.C(n_98),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_140),
.C(n_117),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_147),
.B(n_138),
.Y(n_154)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_129),
.A3(n_128),
.B1(n_117),
.B2(n_120),
.C1(n_125),
.C2(n_118),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_133),
.B1(n_136),
.B2(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_146),
.B1(n_137),
.B2(n_128),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_117),
.B1(n_100),
.B2(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_154),
.C(n_141),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_135),
.B1(n_143),
.B2(n_132),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_148),
.B1(n_119),
.B2(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_149),
.A3(n_154),
.B1(n_152),
.B2(n_101),
.C1(n_122),
.C2(n_86),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_153),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_158),
.B1(n_86),
.B2(n_60),
.C(n_13),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_163),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C(n_12),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_11),
.A3(n_12),
.B1(n_60),
.B2(n_159),
.C1(n_40),
.C2(n_52),
.Y(n_165)
);


endmodule