module fake_netlist_5_2422_n_1062 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1062);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1062;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_947;
wire n_757;
wire n_820;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_723;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_952;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_80),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_62),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_52),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_42),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_16),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_13),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_27),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_99),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_51),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_33),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_113),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_61),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_22),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_141),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_118),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_144),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_90),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_95),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_47),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_29),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_54),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_195),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_101),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_167),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_139),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_77),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_111),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_177),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_49),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_87),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_166),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_67),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_217),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_202),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_203),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_227),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_204),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_217),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_213),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_206),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_208),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_230),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_215),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_223),
.Y(n_295)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_0),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_242),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_233),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_221),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_234),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_226),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_257),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_213),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_228),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_213),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_256),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_268),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_257),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_275),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_270),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_272),
.A2(n_265),
.B1(n_250),
.B2(n_236),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_300),
.B(n_265),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_267),
.A2(n_207),
.B1(n_258),
.B2(n_259),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_207),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx11_ASAP7_75t_R g348 ( 
.A(n_267),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_282),
.B(n_231),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_309),
.A2(n_235),
.B(n_232),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_311),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_278),
.A2(n_258),
.B1(n_259),
.B2(n_248),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_L g359 ( 
.A(n_294),
.B(n_241),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_240),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_254),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_279),
.B(n_244),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_255),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_285),
.B(n_260),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_360),
.B(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_261),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

NOR2x1p5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_246),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_263),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

BUFx6f_ASAP7_75t_SL g382 ( 
.A(n_367),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_347),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_347),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_264),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_348),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_352),
.B(n_251),
.Y(n_398)
);

AND3x2_ASAP7_75t_L g399 ( 
.A(n_316),
.B(n_0),
.C(n_1),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_334),
.A2(n_247),
.B1(n_249),
.B2(n_253),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_358),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_343),
.B(n_291),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_353),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

NOR2x1p5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_262),
.Y(n_417)
);

AND3x2_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_1),
.C(n_2),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_345),
.B(n_291),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

BUFx6f_ASAP7_75t_SL g433 ( 
.A(n_367),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_333),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_332),
.B(n_34),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_357),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_432),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_378),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_315),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

OR2x2_ASAP7_75t_SL g445 ( 
.A(n_438),
.B(n_340),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_386),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_397),
.B(n_325),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_368),
.B(n_324),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_428),
.A2(n_363),
.B(n_362),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_439),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_325),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_386),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_375),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_429),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_319),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_375),
.Y(n_462)
);

XNOR2x2_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_329),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_315),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_361),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_368),
.B(n_355),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_400),
.B(n_304),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_390),
.Y(n_471)
);

INVx4_ASAP7_75t_SL g472 ( 
.A(n_436),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_390),
.B(n_367),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_403),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_374),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_388),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_341),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_304),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_366),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_391),
.B(n_359),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

XNOR2x2_ASAP7_75t_L g492 ( 
.A(n_399),
.B(n_338),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_371),
.B(n_364),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_387),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

OR2x2_ASAP7_75t_SL g500 ( 
.A(n_398),
.B(n_366),
.Y(n_500)
);

INVx4_ASAP7_75t_SL g501 ( 
.A(n_382),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_428),
.A2(n_322),
.B(n_359),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_382),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_392),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_382),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_371),
.B(n_364),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_393),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_341),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_391),
.B(n_312),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_384),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_454),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_464),
.A2(n_338),
.B1(n_377),
.B2(n_391),
.Y(n_518)
);

O2A1O1Ixp33_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_345),
.B(n_377),
.C(n_344),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_459),
.B(n_278),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_464),
.B(n_391),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_443),
.B(n_417),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_460),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_466),
.B(n_414),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_440),
.B(n_416),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_411),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_444),
.B(n_416),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_401),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g532 ( 
.A(n_448),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_419),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_421),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_470),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_421),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_449),
.B(n_332),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_468),
.B(n_382),
.Y(n_538)
);

BUFx5_ASAP7_75t_L g539 ( 
.A(n_498),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_451),
.B(n_446),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_461),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_494),
.B(n_415),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_424),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_477),
.B(n_424),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_468),
.B(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_425),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_425),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_458),
.A2(n_430),
.B1(n_433),
.B2(n_337),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_480),
.B(n_420),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_465),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_473),
.B(n_346),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_441),
.B(n_433),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_483),
.B(n_422),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_489),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_433),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_514),
.B(n_418),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_489),
.B(n_354),
.Y(n_559)
);

NAND2x1_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_402),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_452),
.B(n_422),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_486),
.B(n_423),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_476),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_488),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_504),
.B(n_426),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_472),
.B(n_426),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_426),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_508),
.B(n_427),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_471),
.A2(n_372),
.B(n_370),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_442),
.B(n_427),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_472),
.B(n_384),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_485),
.B(n_402),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_487),
.B(n_384),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_499),
.B(n_402),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_SL g576 ( 
.A(n_520),
.B(n_462),
.C(n_456),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_527),
.B(n_463),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_SL g578 ( 
.A(n_538),
.B(n_469),
.C(n_471),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_491),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_571),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_532),
.A2(n_453),
.B1(n_500),
.B2(n_445),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_535),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_569),
.B(n_501),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_535),
.B(n_501),
.Y(n_586)
);

NOR3xp33_ASAP7_75t_SL g587 ( 
.A(n_558),
.B(n_492),
.C(n_510),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_559),
.Y(n_588)
);

NOR2x1_ASAP7_75t_R g589 ( 
.A(n_535),
.B(n_566),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_556),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_541),
.B(n_493),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_521),
.B(n_534),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_551),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_521),
.B(n_496),
.Y(n_596)
);

CKINVDCx14_ASAP7_75t_R g597 ( 
.A(n_574),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_540),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_522),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_553),
.B(n_497),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_518),
.B(n_502),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_557),
.B(n_501),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_525),
.Y(n_605)
);

CKINVDCx6p67_ASAP7_75t_R g606 ( 
.A(n_529),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_SL g607 ( 
.A(n_549),
.B(n_512),
.C(n_511),
.Y(n_607)
);

OR2x2_ASAP7_75t_SL g608 ( 
.A(n_524),
.B(n_515),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_531),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_548),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_552),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_549),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_543),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_564),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_554),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_528),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_560),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_544),
.B(n_505),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_548),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_575),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_536),
.B(n_506),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_519),
.B(n_507),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_447),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_572),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_567),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_545),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_539),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_539),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_617),
.Y(n_638)
);

BUFx2_ASAP7_75t_SL g639 ( 
.A(n_583),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_581),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_577),
.B(n_618),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_594),
.A2(n_526),
.B(n_546),
.Y(n_642)
);

NAND2x1p5_ASAP7_75t_L g643 ( 
.A(n_628),
.B(n_478),
.Y(n_643)
);

AOI21xp33_ASAP7_75t_L g644 ( 
.A1(n_577),
.A2(n_547),
.B(n_550),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_594),
.A2(n_555),
.B(n_562),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_580),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_586),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_621),
.B(n_563),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_628),
.A2(n_570),
.B(n_484),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_588),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_597),
.B(n_475),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_628),
.B(n_478),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_583),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_584),
.B(n_481),
.Y(n_654)
);

AND3x4_ASAP7_75t_L g655 ( 
.A(n_587),
.B(n_408),
.C(n_513),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_478),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_636),
.A2(n_495),
.B(n_482),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_607),
.A2(n_632),
.B(n_614),
.C(n_622),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_582),
.A2(n_539),
.B1(n_370),
.B2(n_373),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_610),
.B(n_408),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_634),
.A2(n_478),
.B(n_330),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_591),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_584),
.B(n_395),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_601),
.B(n_395),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_627),
.A2(n_435),
.A3(n_431),
.B(n_374),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_606),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_609),
.A2(n_619),
.B(n_627),
.Y(n_668)
);

OAI22x1_ASAP7_75t_L g669 ( 
.A1(n_590),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_619),
.A2(n_592),
.B(n_579),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_600),
.A2(n_407),
.B1(n_396),
.B2(n_395),
.Y(n_671)
);

AO31x2_ASAP7_75t_L g672 ( 
.A1(n_603),
.A2(n_435),
.A3(n_431),
.B(n_407),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_623),
.B(n_395),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_596),
.A2(n_407),
.B(n_396),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_586),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_596),
.A2(n_407),
.B(n_396),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_396),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_595),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_600),
.A2(n_435),
.B1(n_431),
.B2(n_5),
.Y(n_679)
);

AOI21x1_ASAP7_75t_SL g680 ( 
.A1(n_579),
.A2(n_3),
.B(n_4),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_620),
.A2(n_615),
.B(n_578),
.C(n_605),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_625),
.B(n_5),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_626),
.B(n_6),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_592),
.A2(n_37),
.B(n_36),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_624),
.A2(n_629),
.B(n_633),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_586),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_631),
.B(n_41),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_578),
.B(n_7),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_629),
.A2(n_114),
.A3(n_199),
.B(n_197),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_668),
.A2(n_604),
.B(n_613),
.Y(n_690)
);

OA21x2_ASAP7_75t_L g691 ( 
.A1(n_670),
.A2(n_616),
.B(n_612),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_641),
.B(n_599),
.Y(n_692)
);

AOI221xp5_ASAP7_75t_SL g693 ( 
.A1(n_669),
.A2(n_608),
.B1(n_602),
.B2(n_591),
.C(n_593),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_651),
.A2(n_576),
.B1(n_593),
.B2(n_611),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_685),
.A2(n_631),
.B(n_635),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_658),
.A2(n_630),
.B(n_601),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_638),
.B(n_593),
.Y(n_700)
);

OAI22x1_ASAP7_75t_L g701 ( 
.A1(n_660),
.A2(n_601),
.B1(n_589),
.B2(n_611),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_649),
.A2(n_591),
.B(n_44),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_645),
.A2(n_45),
.B(n_43),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_647),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_648),
.B(n_585),
.Y(n_705)
);

AO21x1_ASAP7_75t_L g706 ( 
.A1(n_684),
.A2(n_8),
.B(n_9),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_659),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_707)
);

CKINVDCx6p67_ASAP7_75t_R g708 ( 
.A(n_647),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_678),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_SL g710 ( 
.A1(n_681),
.A2(n_53),
.B(n_50),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_646),
.B(n_10),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_682),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_683),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_673),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_675),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_667),
.A2(n_687),
.B1(n_688),
.B2(n_677),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_674),
.A2(n_56),
.B(n_55),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_644),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_661),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_676),
.A2(n_123),
.B(n_196),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_646),
.B(n_14),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_679),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_654),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_642),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_654),
.B(n_17),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_666),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_675),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_671),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_663),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_662),
.A2(n_127),
.B(n_193),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_23),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_664),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_664),
.B(n_26),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_637),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_643),
.A2(n_200),
.B(n_129),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_57),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_652),
.A2(n_131),
.B(n_189),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_656),
.A2(n_128),
.B(n_188),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_672),
.A2(n_28),
.A3(n_30),
.B(n_31),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_SL g741 ( 
.A1(n_657),
.A2(n_31),
.B(n_58),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_653),
.B(n_60),
.Y(n_742)
);

AO31x2_ASAP7_75t_L g743 ( 
.A1(n_672),
.A2(n_191),
.A3(n_64),
.B(n_65),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_639),
.A2(n_63),
.B(n_66),
.C(n_68),
.Y(n_744)
);

AO21x1_ASAP7_75t_L g745 ( 
.A1(n_680),
.A2(n_69),
.B(n_70),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_657),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_665),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_746),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_716),
.A2(n_655),
.B1(n_689),
.B2(n_74),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_707),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_706),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_694),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_730),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_709),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

CKINVDCx11_ASAP7_75t_R g756 ( 
.A(n_746),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_705),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_712),
.A2(n_97),
.B1(n_100),
.B2(n_103),
.Y(n_759)
);

INVx8_ASAP7_75t_L g760 ( 
.A(n_704),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_713),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_691),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_703),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_704),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_692),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_765)
);

AOI22x1_ASAP7_75t_L g766 ( 
.A1(n_701),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_725),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_741),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_699),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_724),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_714),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_740),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_698),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_711),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_740),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_698),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_704),
.Y(n_778)
);

CKINVDCx8_ASAP7_75t_R g779 ( 
.A(n_737),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_726),
.A2(n_137),
.B1(n_140),
.B2(n_143),
.Y(n_780)
);

BUFx2_ASAP7_75t_SL g781 ( 
.A(n_728),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_720),
.Y(n_782)
);

CKINVDCx11_ASAP7_75t_R g783 ( 
.A(n_747),
.Y(n_783)
);

BUFx8_ASAP7_75t_L g784 ( 
.A(n_732),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_728),
.Y(n_785)
);

BUFx4f_ASAP7_75t_SL g786 ( 
.A(n_715),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_745),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_787)
);

BUFx8_ASAP7_75t_SL g788 ( 
.A(n_717),
.Y(n_788)
);

INVx6_ASAP7_75t_L g789 ( 
.A(n_700),
.Y(n_789)
);

CKINVDCx11_ASAP7_75t_R g790 ( 
.A(n_722),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_717),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_742),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_693),
.B(n_153),
.Y(n_794)
);

INVx6_ASAP7_75t_L g795 ( 
.A(n_734),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_735),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_723),
.A2(n_733),
.B1(n_710),
.B2(n_719),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_727),
.Y(n_799)
);

INVx4_ASAP7_75t_SL g800 ( 
.A(n_729),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_702),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_757),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_743),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_800),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_801),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_801),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_762),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_773),
.A2(n_690),
.B(n_776),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_800),
.Y(n_809)
);

BUFx4f_ASAP7_75t_SL g810 ( 
.A(n_764),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_801),
.B(n_743),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_798),
.A2(n_718),
.B(n_731),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_755),
.B(n_743),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_782),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_772),
.Y(n_815)
);

CKINVDCx6p67_ASAP7_75t_R g816 ( 
.A(n_760),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_796),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_799),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_799),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_749),
.A2(n_721),
.B(n_697),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_774),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_754),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_796),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_777),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_791),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_791),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_791),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_766),
.A2(n_738),
.B(n_736),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_794),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_781),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_785),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_775),
.B(n_744),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_785),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_770),
.Y(n_834)
);

OA21x2_ASAP7_75t_L g835 ( 
.A1(n_787),
.A2(n_739),
.B(n_158),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_778),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_778),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_795),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_771),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_795),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_786),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_802),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_814),
.Y(n_843)
);

INVx4_ASAP7_75t_SL g844 ( 
.A(n_817),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_802),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_821),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_817),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_807),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_807),
.B(n_751),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_809),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_813),
.B(n_779),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_834),
.B(n_784),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_819),
.B(n_752),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_813),
.B(n_790),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_814),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_815),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_834),
.B(n_784),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_808),
.A2(n_797),
.B(n_769),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_815),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_804),
.B(n_809),
.Y(n_860)
);

INVx4_ASAP7_75t_SL g861 ( 
.A(n_817),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_822),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_803),
.B(n_760),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_808),
.A2(n_761),
.B(n_759),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_817),
.B(n_748),
.Y(n_866)
);

OR2x6_ASAP7_75t_L g867 ( 
.A(n_804),
.B(n_789),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_821),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_816),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_SL g870 ( 
.A1(n_849),
.A2(n_832),
.B1(n_753),
.B2(n_750),
.C(n_829),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_842),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_846),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_842),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_846),
.B(n_818),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_868),
.B(n_829),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_845),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_860),
.B(n_819),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_845),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_848),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_860),
.B(n_818),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_856),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_860),
.B(n_818),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_860),
.B(n_803),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_859),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_856),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_850),
.B(n_840),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_850),
.B(n_840),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_859),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_854),
.B(n_840),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_872),
.Y(n_891)
);

AO21x2_ASAP7_75t_L g892 ( 
.A1(n_885),
.A2(n_858),
.B(n_830),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_884),
.B(n_854),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_876),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_884),
.B(n_851),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_871),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_878),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_878),
.B(n_844),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_878),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_881),
.B(n_851),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_890),
.B(n_862),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_890),
.B(n_862),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_881),
.B(n_844),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_883),
.B(n_867),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_894),
.B(n_887),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_891),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_891),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_900),
.B(n_888),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_901),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_900),
.B(n_888),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_902),
.B(n_849),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_896),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_892),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_895),
.B(n_883),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_898),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_893),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_896),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_892),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_SL g920 ( 
.A1(n_917),
.A2(n_893),
.B(n_895),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_SL g921 ( 
.A1(n_915),
.A2(n_904),
.B(n_905),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_907),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_916),
.B(n_903),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_916),
.B(n_898),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_908),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_909),
.B(n_903),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_910),
.B(n_897),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_918),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_927),
.B(n_911),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_923),
.B(n_897),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_924),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_927),
.B(n_912),
.Y(n_932)
);

NOR4xp25_ASAP7_75t_SL g933 ( 
.A(n_928),
.B(n_899),
.C(n_925),
.D(n_922),
.Y(n_933)
);

AO221x2_ASAP7_75t_L g934 ( 
.A1(n_921),
.A2(n_920),
.B1(n_852),
.B2(n_857),
.C(n_841),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_926),
.B(n_906),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_931),
.B(n_924),
.Y(n_936)
);

OAI33xp33_ASAP7_75t_L g937 ( 
.A1(n_932),
.A2(n_929),
.A3(n_935),
.B1(n_933),
.B2(n_919),
.B3(n_913),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_934),
.B(n_924),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_930),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_931),
.B(n_903),
.Y(n_940)
);

AOI32xp33_ASAP7_75t_L g941 ( 
.A1(n_930),
.A2(n_914),
.A3(n_832),
.B1(n_919),
.B2(n_853),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_931),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_931),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_903),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_931),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_942),
.B(n_918),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_937),
.A2(n_858),
.B1(n_892),
.B2(n_898),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_943),
.A2(n_914),
.B(n_899),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_945),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_936),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_939),
.B(n_904),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_940),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_938),
.A2(n_867),
.B1(n_869),
.B2(n_873),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_944),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_947),
.A2(n_941),
.B(n_870),
.C(n_898),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_948),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_946),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_949),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_948),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_941),
.Y(n_960)
);

OAI32xp33_ASAP7_75t_L g961 ( 
.A1(n_951),
.A2(n_952),
.A3(n_954),
.B1(n_953),
.B2(n_873),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_947),
.A2(n_869),
.B1(n_867),
.B2(n_841),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_948),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_960),
.B(n_839),
.Y(n_964)
);

AOI221x1_ASAP7_75t_L g965 ( 
.A1(n_959),
.A2(n_768),
.B1(n_758),
.B2(n_830),
.C(n_765),
.Y(n_965)
);

OAI31xp33_ASAP7_75t_L g966 ( 
.A1(n_955),
.A2(n_963),
.A3(n_962),
.B(n_956),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_957),
.B(n_756),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_963),
.A2(n_866),
.B1(n_838),
.B2(n_789),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_961),
.B(n_783),
.C(n_763),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_958),
.A2(n_867),
.B1(n_810),
.B2(n_816),
.Y(n_970)
);

BUFx12f_ASAP7_75t_L g971 ( 
.A(n_967),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_788),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_968),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_970),
.B(n_838),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_966),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_969),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_965),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_964),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_966),
.B(n_875),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_964),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_966),
.B(n_872),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_971),
.B(n_838),
.Y(n_982)
);

AOI211xp5_ASAP7_75t_L g983 ( 
.A1(n_975),
.A2(n_847),
.B(n_853),
.C(n_817),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_972),
.B(n_875),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_977),
.B(n_847),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_979),
.A2(n_828),
.B(n_823),
.Y(n_986)
);

OA22x2_ASAP7_75t_L g987 ( 
.A1(n_976),
.A2(n_836),
.B1(n_837),
.B2(n_831),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_973),
.B(n_816),
.Y(n_988)
);

XOR2x2_ASAP7_75t_L g989 ( 
.A(n_978),
.B(n_853),
.Y(n_989)
);

NOR2xp67_ASAP7_75t_L g990 ( 
.A(n_980),
.B(n_157),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_981),
.B(n_847),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_SL g992 ( 
.A1(n_981),
.A2(n_847),
.B1(n_817),
.B2(n_823),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_988),
.B(n_985),
.C(n_990),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_982),
.B(n_974),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_989),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_991),
.B(n_831),
.Y(n_996)
);

NAND5xp2_ASAP7_75t_L g997 ( 
.A(n_983),
.B(n_780),
.C(n_792),
.D(n_767),
.E(n_833),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_889),
.Y(n_998)
);

AOI211xp5_ASAP7_75t_L g999 ( 
.A1(n_986),
.A2(n_847),
.B(n_836),
.C(n_837),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_992),
.A2(n_987),
.B1(n_833),
.B2(n_835),
.C(n_827),
.Y(n_1000)
);

OR5x1_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_844),
.C(n_861),
.D(n_827),
.E(n_826),
.Y(n_1001)
);

AOI211xp5_ASAP7_75t_L g1002 ( 
.A1(n_995),
.A2(n_828),
.B(n_825),
.C(n_826),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_889),
.Y(n_1003)
);

NAND4xp25_ASAP7_75t_L g1004 ( 
.A(n_996),
.B(n_999),
.C(n_1000),
.D(n_998),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_997),
.A2(n_885),
.B1(n_877),
.B2(n_874),
.C(n_879),
.Y(n_1005)
);

NAND4xp25_ASAP7_75t_SL g1006 ( 
.A(n_993),
.B(n_825),
.C(n_826),
.D(n_864),
.Y(n_1006)
);

AOI221x1_ASAP7_75t_L g1007 ( 
.A1(n_993),
.A2(n_877),
.B1(n_874),
.B2(n_879),
.C(n_880),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_994),
.B(n_844),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_994),
.B(n_886),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1001),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_1008),
.B(n_825),
.Y(n_1011)
);

NAND4xp75_ASAP7_75t_L g1012 ( 
.A(n_1009),
.B(n_835),
.C(n_865),
.D(n_880),
.Y(n_1012)
);

NAND5xp2_ASAP7_75t_L g1013 ( 
.A(n_1002),
.B(n_1003),
.C(n_1006),
.D(n_1004),
.E(n_1005),
.Y(n_1013)
);

AOI211xp5_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_828),
.B(n_824),
.C(n_864),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1003),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_L g1016 ( 
.A(n_1008),
.B(n_159),
.Y(n_1016)
);

NOR2x1p5_ASAP7_75t_L g1017 ( 
.A(n_1004),
.B(n_806),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_1008),
.B(n_812),
.C(n_806),
.Y(n_1018)
);

AND3x4_ASAP7_75t_L g1019 ( 
.A(n_1016),
.B(n_861),
.C(n_811),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_812),
.C(n_806),
.Y(n_1020)
);

NOR2x1p5_ASAP7_75t_L g1021 ( 
.A(n_1010),
.B(n_806),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_1013),
.B(n_805),
.C(n_820),
.Y(n_1022)
);

XNOR2xp5_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_160),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_1011),
.B(n_861),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_1012),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1014),
.B(n_861),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_161),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_1017),
.B(n_886),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1013),
.B(n_824),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_1016),
.B(n_162),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1017),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1023),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_1031),
.A2(n_858),
.B(n_835),
.C(n_165),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1027),
.A2(n_163),
.B(n_164),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1024),
.B(n_882),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1019),
.Y(n_1037)
);

XNOR2x1_ASAP7_75t_L g1038 ( 
.A(n_1021),
.B(n_168),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1028),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_1022),
.B(n_863),
.C(n_855),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1037),
.A2(n_1025),
.B1(n_1029),
.B2(n_1026),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1039),
.B(n_1020),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_1033),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1032),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1038),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1036),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1043),
.A2(n_1040),
.B1(n_1035),
.B2(n_1034),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1044),
.Y(n_1048)
);

INVx3_ASAP7_75t_SL g1049 ( 
.A(n_1045),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1048),
.A2(n_1041),
.B1(n_1042),
.B2(n_1046),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

AOI222xp33_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_1049),
.B1(n_1047),
.B2(n_805),
.C1(n_843),
.C2(n_863),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1052),
.A2(n_882),
.B1(n_805),
.B2(n_871),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1052),
.A2(n_805),
.B1(n_835),
.B2(n_811),
.Y(n_1054)
);

OAI22xp33_ASAP7_75t_SL g1055 ( 
.A1(n_1052),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_1055),
.B(n_173),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_174),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1053),
.A2(n_175),
.B(n_178),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_1058),
.A2(n_179),
.B(n_182),
.Y(n_1059)
);

OR2x2_ASAP7_75t_SL g1060 ( 
.A(n_1057),
.B(n_183),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_1056),
.B1(n_185),
.B2(n_184),
.C(n_811),
.Y(n_1061)
);

AOI211xp5_ASAP7_75t_L g1062 ( 
.A1(n_1061),
.A2(n_1059),
.B(n_811),
.C(n_820),
.Y(n_1062)
);


endmodule