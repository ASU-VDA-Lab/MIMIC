module real_jpeg_28337_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_5),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_23),
.B1(n_49),
.B2(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_6),
.B(n_49),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_5),
.A2(n_8),
.B(n_32),
.C(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_49),
.B1(n_54),
.B2(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_49),
.B1(n_54),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_9),
.Y(n_72)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_10),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_95),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_94),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_87),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_15),
.B(n_87),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_76),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_66),
.B1(n_74),
.B2(n_75),
.Y(n_16)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_46),
.B2(n_65),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_18),
.A2(n_19),
.B1(n_78),
.B2(n_79),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_34),
.B2(n_45),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_20),
.A2(n_21),
.B1(n_131),
.B2(n_132),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI211xp5_ASAP7_75t_L g92 ( 
.A1(n_21),
.A2(n_57),
.B(n_86),
.C(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_23),
.A2(n_24),
.B(n_30),
.C(n_82),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_23),
.A2(n_40),
.B(n_60),
.C(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_23),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_119),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_23),
.A2(n_39),
.B(n_41),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_34),
.A2(n_45),
.B1(n_57),
.B2(n_73),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_34),
.A2(n_45),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_34),
.B(n_83),
.C(n_143),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_40),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_73),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_45),
.A2(n_73),
.B(n_133),
.C(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_57),
.B1(n_73),
.B2(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_55),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_54),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_73),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_73),
.B1(n_104),
.B2(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_83),
.C(n_108),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_73),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_139),
.C(n_148),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_86),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_84),
.B1(n_107),
.B2(n_111),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_84),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_83),
.A2(n_84),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_89),
.Y(n_167)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_168),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_163),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_151),
.B(n_162),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_135),
.B(n_150),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_124),
.B(n_134),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_112),
.B(n_123),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);


endmodule