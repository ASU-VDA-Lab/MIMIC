module fake_jpeg_17858_n_342 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_42),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_47),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_23),
.A2(n_13),
.B(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_23),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_7),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_48),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_67),
.B(n_71),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_25),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_106),
.B1(n_10),
.B2(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_38),
.A2(n_52),
.B1(n_57),
.B2(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_74),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_27),
.B1(n_14),
.B2(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_39),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_60),
.B1(n_26),
.B2(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_26),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_24),
.B1(n_34),
.B2(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_41),
.B(n_22),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_81),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_0),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_41),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_18),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_18),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_45),
.A2(n_34),
.B(n_21),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_36),
.B(n_9),
.C(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_18),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_38),
.A2(n_34),
.B1(n_21),
.B2(n_19),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_83),
.B1(n_70),
.B2(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_44),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_0),
.Y(n_126)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_36),
.B1(n_0),
.B2(n_4),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_128),
.B1(n_153),
.B2(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_150),
.B1(n_84),
.B2(n_102),
.Y(n_172)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_10),
.B1(n_5),
.B2(n_7),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_123),
.A2(n_124),
.B1(n_155),
.B2(n_157),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_36),
.B1(n_5),
.B2(n_9),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_137),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_5),
.B(n_9),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_135),
.B(n_149),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_84),
.B1(n_102),
.B2(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_11),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_133),
.B(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_72),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_143),
.Y(n_168)
);

NAND2x1p5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_0),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_12),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_104),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_75),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_147),
.Y(n_187)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_74),
.B(n_85),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_85),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_84),
.C(n_102),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_105),
.B(n_89),
.C(n_81),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_161),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_76),
.A2(n_98),
.B1(n_83),
.B2(n_113),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_92),
.B1(n_88),
.B2(n_69),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_69),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_115),
.Y(n_189)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_75),
.B(n_77),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_77),
.A2(n_110),
.B1(n_33),
.B2(n_28),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_155),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_77),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_166),
.C(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_205),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_175),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_169),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_173),
.B1(n_198),
.B2(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_121),
.B1(n_151),
.B2(n_123),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_131),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_178),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_178),
.Y(n_209)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_163),
.B1(n_125),
.B2(n_126),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_193),
.B1(n_182),
.B2(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_122),
.B1(n_117),
.B2(n_147),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_197),
.B(n_202),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_194),
.B(n_179),
.Y(n_220)
);

BUFx24_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_119),
.A2(n_162),
.B1(n_159),
.B2(n_148),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_142),
.A2(n_163),
.B1(n_133),
.B2(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_120),
.B(n_154),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_119),
.B1(n_124),
.B2(n_138),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_171),
.B1(n_179),
.B2(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_119),
.B1(n_135),
.B2(n_140),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_116),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_213),
.C(n_233),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_217),
.B(n_220),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_210),
.B(n_211),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_180),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_221),
.B(n_174),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_217),
.B1(n_209),
.B2(n_206),
.C(n_210),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_199),
.C(n_171),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_216),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_188),
.B(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_188),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_167),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_201),
.B1(n_165),
.B2(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_182),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_177),
.B(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_239),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_170),
.C(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_213),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_174),
.A2(n_205),
.B1(n_170),
.B2(n_183),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_215),
.B1(n_261),
.B2(n_242),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_248),
.B1(n_259),
.B2(n_263),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_165),
.B1(n_196),
.B2(n_229),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_260),
.C(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_209),
.B1(n_228),
.B2(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_221),
.C(n_212),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_262),
.B(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_207),
.B1(n_234),
.B2(n_214),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_223),
.C(n_214),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_227),
.C(n_232),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_264),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_275),
.C(n_279),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_215),
.C(n_241),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_285),
.B1(n_263),
.B2(n_266),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_215),
.C(n_258),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_215),
.CI(n_260),
.CON(n_281),
.SN(n_281)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_265),
.C(n_253),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_287),
.C(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_259),
.A2(n_248),
.B1(n_255),
.B2(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_255),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_242),
.B(n_250),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_288),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_281),
.B1(n_280),
.B2(n_288),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_296),
.B1(n_298),
.B2(n_300),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_245),
.B1(n_247),
.B2(n_252),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_245),
.B1(n_252),
.B2(n_271),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_285),
.B1(n_268),
.B2(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_306),
.C(n_282),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_279),
.C(n_270),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_298),
.B1(n_290),
.B2(n_299),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_278),
.B(n_274),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_316),
.B(n_299),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_287),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_310),
.C(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_280),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_286),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_274),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_283),
.C(n_284),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_318),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_322),
.B(n_301),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_303),
.B1(n_305),
.B2(n_301),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_296),
.B1(n_313),
.B2(n_316),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_303),
.B1(n_305),
.B2(n_304),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_314),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_291),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_332),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_333),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_315),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_327),
.B(n_320),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_334),
.A2(n_333),
.B(n_328),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_338),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_321),
.C(n_325),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_335),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_326),
.Y(n_342)
);


endmodule