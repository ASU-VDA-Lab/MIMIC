module fake_jpeg_11609_n_524 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_524);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_524;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_54),
.A2(n_28),
.B(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_8),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_65),
.Y(n_143)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_26),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_34),
.Y(n_105)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_29),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_100),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_34),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_105),
.B(n_29),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_52),
.A2(n_45),
.B1(n_41),
.B2(n_19),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_110),
.A2(n_41),
.B1(n_45),
.B2(n_19),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_30),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_114),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_30),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_113),
.B(n_61),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_54),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_27),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_49),
.B1(n_42),
.B2(n_43),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_120),
.A2(n_124),
.B1(n_38),
.B2(n_22),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_69),
.A2(n_49),
.B1(n_42),
.B2(n_43),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_126),
.A2(n_141),
.B1(n_22),
.B2(n_31),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_SL g144 ( 
.A(n_67),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_144),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_29),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_153),
.B(n_134),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_70),
.B(n_49),
.C(n_43),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_27),
.Y(n_197)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_143),
.B1(n_110),
.B2(n_80),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_174),
.Y(n_245)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_169),
.Y(n_268)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

OR2x2_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_71),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_172),
.A2(n_184),
.B(n_193),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_173),
.A2(n_194),
.B1(n_203),
.B2(n_209),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_99),
.B1(n_98),
.B2(n_97),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_116),
.A2(n_58),
.B1(n_50),
.B2(n_81),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_204),
.B1(n_206),
.B2(n_213),
.Y(n_248)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_78),
.B1(n_75),
.B2(n_76),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_182),
.A2(n_156),
.B1(n_127),
.B2(n_139),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_103),
.B(n_34),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_103),
.B(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_198),
.Y(n_224)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_192),
.B(n_196),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_112),
.A2(n_38),
.B(n_47),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_121),
.A2(n_88),
.B1(n_92),
.B2(n_91),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_27),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_200),
.B(n_211),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_106),
.B(n_68),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_210),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_145),
.A2(n_73),
.B1(n_72),
.B2(n_93),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_96),
.B1(n_59),
.B2(n_47),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_31),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_22),
.Y(n_221)
);

AOI32xp33_ASAP7_75t_L g215 ( 
.A1(n_147),
.A2(n_62),
.A3(n_85),
.B1(n_95),
.B2(n_42),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_128),
.A2(n_41),
.B1(n_45),
.B2(n_19),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_47),
.B1(n_196),
.B2(n_188),
.Y(n_256)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_251),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_179),
.A2(n_162),
.B(n_180),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_227),
.A2(n_44),
.B(n_10),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_166),
.B(n_150),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_238),
.B(n_239),
.C(n_17),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_142),
.C(n_140),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_240),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_156),
.B1(n_139),
.B2(n_130),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_241),
.A2(n_188),
.B1(n_174),
.B2(n_217),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_130),
.B1(n_148),
.B2(n_31),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_172),
.A2(n_101),
.B1(n_148),
.B2(n_104),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_193),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_267),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_173),
.A2(n_101),
.B1(n_23),
.B2(n_64),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_174),
.A2(n_23),
.B1(n_44),
.B2(n_2),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_178),
.B1(n_175),
.B2(n_167),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_0),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_171),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_272),
.A2(n_276),
.B1(n_242),
.B2(n_246),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_213),
.B1(n_209),
.B2(n_212),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_287),
.B1(n_288),
.B2(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_211),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_279),
.C(n_292),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_161),
.B1(n_165),
.B2(n_170),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_206),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_278),
.B(n_282),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_239),
.C(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_302),
.Y(n_318)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_230),
.A2(n_204),
.B1(n_201),
.B2(n_195),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_283),
.A2(n_297),
.B1(n_306),
.B2(n_316),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_245),
.A2(n_44),
.B1(n_167),
.B2(n_4),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_289),
.A2(n_300),
.B(n_242),
.C(n_220),
.Y(n_345)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_222),
.B(n_0),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_314),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_44),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_293),
.B(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_10),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_296),
.Y(n_352)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_10),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_298),
.B(n_303),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_237),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_312),
.Y(n_336)
);

AO21x2_ASAP7_75t_SL g300 ( 
.A1(n_262),
.A2(n_1),
.B(n_4),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_245),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_221),
.B(n_1),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_223),
.B(n_224),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_304),
.A2(n_310),
.B1(n_315),
.B2(n_300),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_243),
.A2(n_253),
.B(n_257),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_279),
.B(n_275),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_248),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_253),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_234),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_223),
.B(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_231),
.Y(n_313)
);

INVx11_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_240),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_229),
.A2(n_1),
.B1(n_7),
.B2(n_12),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_317),
.A2(n_326),
.B(n_310),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_285),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_323),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_281),
.A2(n_224),
.B1(n_243),
.B2(n_247),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_328),
.B1(n_329),
.B2(n_342),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_254),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_237),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_330),
.C(n_353),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_286),
.A2(n_268),
.B1(n_263),
.B2(n_265),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_286),
.A2(n_268),
.B1(n_265),
.B2(n_233),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_252),
.C(n_259),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_249),
.B(n_267),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_331),
.A2(n_332),
.B(n_309),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_249),
.B(n_252),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_340),
.B1(n_350),
.B2(n_313),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_283),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_300),
.A2(n_233),
.B1(n_246),
.B2(n_259),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_284),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_348),
.Y(n_370)
);

AO21x2_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_272),
.B(n_294),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_300),
.A2(n_246),
.B1(n_269),
.B2(n_266),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_347),
.B1(n_351),
.B2(n_354),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_300),
.A2(n_308),
.B1(n_314),
.B2(n_280),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_277),
.B(n_269),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_306),
.A2(n_232),
.B1(n_220),
.B2(n_250),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_287),
.A2(n_228),
.B1(n_250),
.B2(n_232),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_284),
.A2(n_228),
.B1(n_232),
.B2(n_231),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_7),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_356),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_360),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_372),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_291),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_363),
.C(n_371),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_291),
.Y(n_363)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_327),
.B(n_316),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_368),
.B(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_321),
.B(n_303),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_380),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_278),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_357),
.B(n_274),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_383),
.B1(n_322),
.B2(n_347),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_334),
.B(n_278),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_375),
.A2(n_340),
.B1(n_345),
.B2(n_346),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_296),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_378),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_334),
.B(n_301),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_377),
.B(n_352),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_293),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_331),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_341),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_307),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_382),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_326),
.A2(n_297),
.B1(n_315),
.B2(n_304),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_282),
.Y(n_384)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_356),
.Y(n_397)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_271),
.Y(n_388)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_311),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_389),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_290),
.Y(n_390)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_356),
.A2(n_7),
.B(n_14),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_335),
.B(n_339),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_336),
.B(n_16),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_392),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_345),
.Y(n_446)
);

AOI22x1_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_328),
.B1(n_329),
.B2(n_342),
.Y(n_399)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_400),
.A2(n_375),
.B1(n_358),
.B2(n_365),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_405),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_348),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_407),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_408),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_375),
.A2(n_337),
.B1(n_343),
.B2(n_318),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_418),
.B1(n_420),
.B2(n_359),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_411),
.B(n_387),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_421),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_343),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_413),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_379),
.A2(n_345),
.B(n_337),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_385),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_375),
.A2(n_365),
.B1(n_358),
.B2(n_366),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_381),
.B(n_319),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_378),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_376),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_444),
.Y(n_452)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_398),
.B(n_360),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_428),
.B(n_442),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_415),
.B1(n_405),
.B2(n_421),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_414),
.B(n_425),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_382),
.C(n_374),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_433),
.C(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_393),
.C(n_362),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_434),
.A2(n_435),
.B1(n_440),
.B2(n_443),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_420),
.A2(n_409),
.B1(n_418),
.B2(n_404),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_371),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_437),
.B(n_439),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_393),
.B(n_363),
.C(n_377),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_368),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_404),
.A2(n_383),
.B1(n_375),
.B2(n_323),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_446),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_398),
.B(n_419),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_351),
.B1(n_345),
.B2(n_354),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_355),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_319),
.C(n_333),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_422),
.C(n_408),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_425),
.Y(n_450)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_416),
.B1(n_412),
.B2(n_397),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_440),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_458),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_397),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_462),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_435),
.A2(n_400),
.B1(n_396),
.B2(n_401),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_447),
.A2(n_416),
.B1(n_394),
.B2(n_395),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_434),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_394),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_396),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_463),
.B(n_466),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_417),
.B(n_413),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_467),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_431),
.B(n_401),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_437),
.B(n_395),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_444),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_455),
.A2(n_447),
.B1(n_454),
.B2(n_423),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_470),
.A2(n_448),
.B1(n_453),
.B2(n_443),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_438),
.C(n_426),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_472),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_427),
.C(n_439),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_457),
.C(n_452),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_461),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_432),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_478),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_407),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_480),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_451),
.A2(n_446),
.B1(n_441),
.B2(n_399),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_482),
.B1(n_483),
.B2(n_475),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_490),
.B1(n_476),
.B2(n_386),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_484),
.A2(n_451),
.B1(n_460),
.B2(n_465),
.Y(n_490)
);

OAI321xp33_ASAP7_75t_L g492 ( 
.A1(n_470),
.A2(n_459),
.A3(n_399),
.B1(n_406),
.B2(n_460),
.C(n_333),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_452),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_495),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_471),
.A2(n_456),
.B(n_464),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_464),
.C(n_406),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_349),
.C(n_16),
.Y(n_506)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_491),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_499),
.B(n_485),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_497),
.A2(n_479),
.B1(n_481),
.B2(n_473),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_501),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_391),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_504),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_339),
.B(n_349),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_16),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_496),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_511),
.B(n_512),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_507),
.B(n_490),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_513),
.B(n_508),
.Y(n_515)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_510),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_514),
.A2(n_517),
.B(n_506),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_515),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_498),
.C(n_502),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_500),
.B(n_503),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_520),
.A2(n_516),
.B(n_518),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_493),
.B(n_16),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_493),
.C(n_17),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_523),
.Y(n_524)
);


endmodule