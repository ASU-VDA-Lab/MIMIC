module fake_jpeg_27560_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_34),
.Y(n_55)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_50),
.B1(n_59),
.B2(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_33),
.B1(n_22),
.B2(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_33),
.B1(n_18),
.B2(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_33),
.B1(n_24),
.B2(n_34),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_45),
.B1(n_44),
.B2(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_47),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_17),
.B(n_30),
.C(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_77),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_45),
.B1(n_55),
.B2(n_65),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_47),
.C(n_20),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_68),
.C(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_82),
.Y(n_99)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_113),
.Y(n_122)
);

OA22x2_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_82),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_84),
.B1(n_52),
.B2(n_72),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_51),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_17),
.B1(n_45),
.B2(n_58),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_49),
.B1(n_60),
.B2(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_49),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_57),
.B1(n_42),
.B2(n_66),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_20),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_121),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_68),
.C(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_131),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_68),
.B(n_73),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_127),
.B(n_133),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_39),
.B(n_68),
.C(n_77),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_93),
.B1(n_87),
.B2(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_142),
.B1(n_103),
.B2(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_71),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_16),
.B(n_2),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_20),
.C(n_35),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_34),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_111),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_141),
.B(n_117),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_25),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_52),
.B1(n_42),
.B2(n_32),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_147),
.B(n_151),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_114),
.B1(n_103),
.B2(n_107),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_165),
.B1(n_110),
.B2(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_104),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_160),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_155),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_139),
.B(n_125),
.Y(n_168)
);

AO22x2_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_117),
.B1(n_114),
.B2(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_34),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_35),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_42),
.B1(n_75),
.B2(n_110),
.Y(n_165)
);

OAI322xp33_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_141),
.A3(n_120),
.B1(n_121),
.B2(n_137),
.C1(n_140),
.C2(n_139),
.Y(n_166)
);

OAI322xp33_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_150),
.A3(n_161),
.B1(n_162),
.B2(n_156),
.C1(n_145),
.C2(n_158),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_180),
.B(n_3),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_144),
.B1(n_158),
.B2(n_145),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_136),
.C(n_41),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_152),
.C(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_178),
.Y(n_193)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_35),
.B(n_28),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_191),
.Y(n_203)
);

OA21x2_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_168),
.B(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_151),
.B1(n_147),
.B2(n_144),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_194),
.B1(n_171),
.B2(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_41),
.B1(n_28),
.B2(n_25),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_201),
.B1(n_174),
.B2(n_173),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_25),
.C(n_37),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_37),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_1),
.B(n_2),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_5),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_178),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_200),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_207),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_185),
.B(n_179),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_209),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_171),
.B1(n_176),
.B2(n_173),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_167),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_215),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_183),
.C(n_172),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_196),
.C(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_213),
.B(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_192),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_183),
.B(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_224),
.B(n_6),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_203),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_225),
.B(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_195),
.B1(n_211),
.B2(n_9),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_6),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_236),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_212),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_229),
.A2(n_8),
.B(n_9),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_8),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_240),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_228),
.B1(n_10),
.B2(n_11),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_8),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_10),
.B(n_12),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_10),
.B(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_41),
.C(n_37),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_12),
.C(n_246),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_12),
.Y(n_248)
);


endmodule