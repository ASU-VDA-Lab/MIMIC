module fake_jpeg_14172_n_558 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_558);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_558;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_62),
.B(n_66),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_69),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_94),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_71),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_82),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_83),
.B(n_104),
.Y(n_175)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_84),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_59),
.B1(n_57),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_27),
.B1(n_56),
.B2(n_53),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_87),
.Y(n_165)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_93),
.B(n_36),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_16),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_106),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_58),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_1),
.C(n_2),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_2),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_124),
.Y(n_153)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_28),
.Y(n_120)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_41),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_16),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_46),
.B1(n_55),
.B2(n_54),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_127),
.A2(n_129),
.B1(n_142),
.B2(n_169),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_55),
.B1(n_46),
.B2(n_42),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_84),
.A2(n_42),
.B1(n_37),
.B2(n_55),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_131),
.A2(n_134),
.B1(n_141),
.B2(n_145),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_37),
.B1(n_28),
.B2(n_38),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_41),
.CON(n_135),
.SN(n_135)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_135),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_136),
.B(n_148),
.Y(n_254)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_36),
.CON(n_139),
.SN(n_139)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_120),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_91),
.A2(n_75),
.B1(n_63),
.B2(n_68),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_64),
.A2(n_45),
.B1(n_39),
.B2(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_27),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_45),
.B1(n_39),
.B2(n_40),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_154),
.A2(n_160),
.B1(n_168),
.B2(n_174),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_64),
.A2(n_48),
.B1(n_44),
.B2(n_56),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_53),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_199),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_74),
.A2(n_48),
.B1(n_44),
.B2(n_47),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_109),
.A2(n_47),
.B1(n_30),
.B2(n_26),
.Y(n_169)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_71),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_203),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_72),
.A2(n_30),
.B1(n_4),
.B2(n_7),
.Y(n_174)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_72),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_188),
.B1(n_78),
.B2(n_119),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_77),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_188)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_80),
.B(n_3),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_77),
.B(n_88),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_205),
.A2(n_226),
.B(n_248),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_211),
.Y(n_275)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_140),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_129),
.A2(n_92),
.B1(n_101),
.B2(n_113),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_213),
.A2(n_268),
.B1(n_128),
.B2(n_183),
.Y(n_281)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_214),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_153),
.B1(n_143),
.B2(n_168),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_215),
.A2(n_240),
.B1(n_252),
.B2(n_257),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_217),
.A2(n_218),
.B1(n_249),
.B2(n_255),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_125),
.A2(n_154),
.B1(n_180),
.B2(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_161),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_231),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_123),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_222),
.B(n_223),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_117),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_114),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_102),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_67),
.C(n_100),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_232),
.C(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_156),
.B(n_103),
.C(n_71),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_237),
.Y(n_276)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_12),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_250),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_134),
.A2(n_121),
.B1(n_118),
.B2(n_87),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_160),
.B(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_258),
.Y(n_282)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_245),
.Y(n_287)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_189),
.B(n_98),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_150),
.A2(n_138),
.B1(n_157),
.B2(n_147),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_193),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_131),
.A2(n_58),
.B1(n_14),
.B2(n_16),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_182),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_171),
.A2(n_176),
.B1(n_192),
.B2(n_137),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_162),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_141),
.A2(n_188),
.B1(n_177),
.B2(n_145),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_159),
.Y(n_259)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_193),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_150),
.B(n_144),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_128),
.C(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_130),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_130),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_155),
.A2(n_137),
.B1(n_170),
.B2(n_190),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_266),
.A2(n_252),
.B1(n_230),
.B2(n_246),
.Y(n_317)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_170),
.A2(n_190),
.B1(n_155),
.B2(n_139),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_147),
.B(n_157),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_138),
.Y(n_292)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_151),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_200),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_277),
.B(n_291),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_281),
.A2(n_298),
.B1(n_266),
.B2(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_225),
.A2(n_215),
.B1(n_240),
.B2(n_257),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_288),
.A2(n_317),
.B1(n_315),
.B2(n_301),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_204),
.B(n_151),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_292),
.B(n_310),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_231),
.B(n_184),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_309),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_184),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_297),
.B(n_316),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_305),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_208),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_239),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_244),
.A2(n_261),
.B(n_205),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_324),
.B(n_326),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_205),
.B(n_226),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_237),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_219),
.C(n_232),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_258),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_311),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_216),
.B(n_219),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_253),
.B(n_248),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_228),
.B(n_207),
.C(n_220),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_323),
.B(n_305),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_271),
.A2(n_262),
.B(n_207),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_262),
.A2(n_235),
.B(n_270),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_317),
.B1(n_324),
.B2(n_323),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_330),
.B1(n_336),
.B2(n_347),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_328),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_247),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_340),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_213),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_333),
.A2(n_358),
.B(n_273),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_334),
.A2(n_335),
.B1(n_341),
.B2(n_333),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_282),
.A2(n_212),
.B1(n_214),
.B2(n_227),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_282),
.A2(n_227),
.B1(n_210),
.B2(n_269),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_275),
.B(n_236),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_281),
.A2(n_210),
.B1(n_269),
.B2(n_272),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_294),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_239),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_351),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_283),
.A2(n_241),
.B1(n_265),
.B2(n_267),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_293),
.A2(n_251),
.B1(n_260),
.B2(n_245),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_352),
.B1(n_364),
.B2(n_365),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_319),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_283),
.A2(n_245),
.B1(n_274),
.B2(n_310),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_279),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_359),
.Y(n_398)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_299),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_276),
.B(n_309),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_289),
.B(n_303),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_287),
.C(n_320),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_279),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_303),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_274),
.A2(n_292),
.B1(n_276),
.B2(n_285),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_291),
.A2(n_290),
.B1(n_326),
.B2(n_311),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_318),
.B(n_290),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

OAI22x1_ASAP7_75t_SL g367 ( 
.A1(n_306),
.A2(n_305),
.B1(n_321),
.B2(n_277),
.Y(n_367)
);

AO21x2_ASAP7_75t_L g396 ( 
.A1(n_367),
.A2(n_342),
.B(n_352),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_337),
.A2(n_312),
.B(n_321),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_365),
.A2(n_336),
.B1(n_327),
.B2(n_334),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_335),
.B1(n_341),
.B2(n_329),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_361),
.B(n_313),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_335),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_334),
.A2(n_312),
.B1(n_296),
.B2(n_313),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_378),
.B1(n_380),
.B2(n_383),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_322),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_384),
.C(n_387),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_330),
.A2(n_296),
.B1(n_322),
.B2(n_304),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_327),
.A2(n_304),
.B1(n_320),
.B2(n_307),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_365),
.A2(n_284),
.B1(n_307),
.B2(n_302),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_284),
.C(n_273),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_337),
.A2(n_302),
.B1(n_280),
.B2(n_325),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_388),
.A2(n_395),
.B1(n_399),
.B2(n_347),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_389),
.A2(n_392),
.B(n_393),
.Y(n_403)
);

A2O1A1O1Ixp25_ASAP7_75t_L g392 ( 
.A1(n_338),
.A2(n_280),
.B(n_286),
.C(n_325),
.D(n_364),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_358),
.A2(n_332),
.B(n_353),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_356),
.A2(n_342),
.B1(n_359),
.B2(n_333),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_367),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_356),
.A2(n_358),
.B1(n_338),
.B2(n_341),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_372),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_417),
.C(n_418),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_350),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_406),
.A2(n_398),
.B(n_392),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_394),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_407),
.B(n_410),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_362),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_374),
.B(n_343),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_394),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_413),
.A2(n_425),
.B1(n_370),
.B2(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_374),
.B(n_366),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_379),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_416),
.A2(n_378),
.B1(n_375),
.B2(n_380),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_349),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_349),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_349),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_419),
.B(n_422),
.Y(n_459)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_349),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_388),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_347),
.B1(n_367),
.B2(n_350),
.Y(n_425)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_401),
.B(n_340),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_427),
.B(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_387),
.C(n_393),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_396),
.Y(n_452)
);

XNOR2x1_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_385),
.Y(n_446)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_434),
.B(n_435),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_437),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_439),
.A2(n_440),
.B1(n_442),
.B2(n_444),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_430),
.A2(n_399),
.B1(n_389),
.B2(n_397),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_430),
.A2(n_397),
.B1(n_370),
.B2(n_391),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_390),
.B1(n_396),
.B2(n_381),
.Y(n_444)
);

XOR2x2_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_331),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_448),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_403),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_449),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_396),
.B1(n_392),
.B2(n_381),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_415),
.C(n_418),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_425),
.A2(n_406),
.B1(n_411),
.B2(n_426),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_411),
.A2(n_402),
.B1(n_400),
.B2(n_386),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_346),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_456),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_405),
.B(n_348),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_445),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_466),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_442),
.A2(n_423),
.B1(n_412),
.B2(n_431),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_478),
.B1(n_451),
.B2(n_453),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_470),
.Y(n_488)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_412),
.B(n_422),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_471),
.A2(n_473),
.B(n_479),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_415),
.C(n_417),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_477),
.C(n_481),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_SL g473 ( 
.A(n_444),
.B(n_408),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_480),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_432),
.C(n_408),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_439),
.A2(n_429),
.B1(n_424),
.B2(n_421),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_328),
.B(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_428),
.C(n_351),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_482),
.B(n_457),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_477),
.C(n_472),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_443),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g510 ( 
.A(n_486),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_489),
.B1(n_491),
.B2(n_495),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_437),
.B1(n_454),
.B2(n_443),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_467),
.B(n_455),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_476),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_447),
.B1(n_448),
.B2(n_459),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_473),
.A2(n_435),
.B(n_446),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_492),
.A2(n_493),
.B(n_482),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_440),
.B(n_441),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_461),
.A2(n_441),
.B1(n_450),
.B2(n_386),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_494),
.A2(n_465),
.B1(n_469),
.B2(n_460),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_464),
.A2(n_450),
.B1(n_344),
.B2(n_373),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_468),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_500),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_466),
.B(n_331),
.C(n_360),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_461),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_501),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_505),
.Y(n_523)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_504),
.Y(n_527)
);

FAx1_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_460),
.CI(n_465),
.CON(n_506),
.SN(n_506)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_506),
.A2(n_514),
.B1(n_486),
.B2(n_493),
.Y(n_517)
);

OAI221xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_476),
.B1(n_463),
.B2(n_479),
.C(n_481),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_497),
.B1(n_489),
.B2(n_488),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_462),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_511),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_486),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_509),
.B(n_515),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_482),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_496),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_363),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_480),
.B1(n_470),
.B2(n_474),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_498),
.C(n_500),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_519),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_498),
.C(n_495),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_512),
.A2(n_501),
.B1(n_494),
.B2(n_497),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_522),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_487),
.C(n_491),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_528),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_502),
.A2(n_510),
.B1(n_469),
.B2(n_488),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_525),
.A2(n_514),
.B1(n_506),
.B2(n_510),
.Y(n_532)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_373),
.Y(n_533)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_533),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_527),
.B(n_519),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_536),
.B(n_537),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_523),
.A2(n_506),
.B(n_483),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_518),
.B(n_373),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_523),
.B(n_503),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_526),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_534),
.A2(n_517),
.B(n_520),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_539),
.A2(n_534),
.B(n_531),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_522),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_541),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_526),
.Y(n_545)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_545),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_547),
.Y(n_551)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_544),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_550),
.B(n_548),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_552),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_549),
.B(n_543),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_553),
.B(n_542),
.C(n_539),
.Y(n_555)
);

NAND4xp25_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_551),
.C(n_546),
.D(n_531),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_556),
.A2(n_554),
.B(n_538),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_355),
.C(n_554),
.Y(n_558)
);


endmodule