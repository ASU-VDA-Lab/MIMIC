module fake_jpeg_20139_n_343 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_42),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_31),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_31),
.C(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_54),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_50),
.B1(n_39),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_84),
.B1(n_100),
.B2(n_59),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_51),
.B(n_43),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_77),
.Y(n_132)
);

CKINVDCx9p33_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_53),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_59),
.B1(n_68),
.B2(n_64),
.Y(n_116)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_96),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_21),
.B1(n_25),
.B2(n_35),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_59),
.B1(n_60),
.B2(n_38),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_99),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_21),
.B1(n_38),
.B2(n_35),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_112),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_129),
.B(n_92),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_43),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_124),
.B(n_91),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_33),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_111),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_93),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_33),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_28),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_58),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_24),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_26),
.Y(n_160)
);

AOI22x1_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_34),
.B1(n_19),
.B2(n_33),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_138),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_137),
.B(n_34),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_81),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_140),
.B(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_153),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_122),
.B1(n_91),
.B2(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_90),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_104),
.Y(n_166)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_159),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_109),
.C(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_176),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_124),
.B1(n_118),
.B2(n_132),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_169),
.B1(n_180),
.B2(n_155),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_115),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_127),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_118),
.B1(n_98),
.B2(n_89),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_143),
.B1(n_159),
.B2(n_151),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_82),
.B1(n_119),
.B2(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_187),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_30),
.B(n_34),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_19),
.B(n_34),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_158),
.C(n_103),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_114),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_203),
.B1(n_184),
.B2(n_163),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_148),
.B1(n_144),
.B2(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_215),
.B1(n_163),
.B2(n_182),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_135),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_208),
.Y(n_232)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_201),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_142),
.B(n_140),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_197),
.B(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_144),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_140),
.B1(n_155),
.B2(n_119),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_207),
.B(n_167),
.Y(n_233)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_211),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_168),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_17),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_217),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_157),
.B(n_158),
.Y(n_210)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_157),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_216),
.Y(n_240)
);

NOR2x1p5_ASAP7_75t_SL g213 ( 
.A(n_162),
.B(n_117),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_200),
.B1(n_199),
.B2(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_82),
.B1(n_117),
.B2(n_86),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_134),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_134),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_79),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_231),
.B1(n_215),
.B2(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_161),
.C(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_206),
.C(n_194),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_210),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_244),
.B1(n_0),
.B2(n_1),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_167),
.B(n_184),
.C(n_83),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_207),
.B1(n_197),
.B2(n_203),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_239),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_34),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_20),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_20),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_245),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_20),
.B1(n_18),
.B2(n_63),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_20),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_196),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_256),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_259),
.B1(n_239),
.B2(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_201),
.C(n_205),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_236),
.C(n_220),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_201),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_211),
.B(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_17),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_63),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_18),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_2),
.B(n_3),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_238),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_267),
.B1(n_231),
.B2(n_245),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_223),
.Y(n_273)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_256),
.C(n_262),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_224),
.C(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_285),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_227),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_287),
.B(n_290),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_253),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_264),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_257),
.C(n_227),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_224),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_230),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_3),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_246),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_260),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_260),
.B1(n_231),
.B2(n_241),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_271),
.B1(n_269),
.B2(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_309),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_304),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_283),
.B(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_283),
.C(n_18),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_18),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_4),
.C(n_5),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_289),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_291),
.C(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_321),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_288),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_288),
.C(n_6),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_7),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_4),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_6),
.B(n_7),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_305),
.B(n_308),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_331),
.B(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_319),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_308),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_334),
.B(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_7),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_330),
.B(n_9),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_8),
.B(n_9),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_337),
.C(n_11),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_13),
.B(n_10),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_10),
.B(n_12),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_12),
.C(n_339),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);


endmodule