module fake_jpeg_18569_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_20),
.B1(n_34),
.B2(n_32),
.Y(n_59)
);

NAND2x1_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_34),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_34),
.B(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_38),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_36),
.Y(n_65)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_59),
.B1(n_76),
.B2(n_82),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_61),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_39),
.B(n_23),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_67),
.B(n_79),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_36),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_32),
.Y(n_67)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_33),
.CI(n_39),
.CON(n_69),
.SN(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_18),
.B1(n_24),
.B2(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_23),
.B(n_24),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_35),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_37),
.B(n_17),
.C(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_69),
.Y(n_97)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_88),
.B(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_32),
.B(n_35),
.C(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_35),
.B1(n_20),
.B2(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_103),
.B1(n_52),
.B2(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_35),
.B1(n_20),
.B2(n_28),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_79),
.B1(n_82),
.B2(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_73),
.B1(n_85),
.B2(n_77),
.Y(n_117)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_67),
.B1(n_79),
.B2(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_63),
.B1(n_80),
.B2(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_25),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_26),
.C(n_46),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_119),
.B1(n_129),
.B2(n_132),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_68),
.B1(n_72),
.B2(n_56),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_89),
.C(n_112),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_70),
.B1(n_68),
.B2(n_46),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_99),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_28),
.B1(n_19),
.B2(n_15),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_99),
.B1(n_100),
.B2(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_113),
.C(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_21),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_87),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_52),
.B1(n_46),
.B2(n_28),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_139),
.B(n_93),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_90),
.A2(n_15),
.B1(n_27),
.B2(n_16),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_15),
.B1(n_27),
.B2(n_16),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_133),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_19),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_104),
.C(n_12),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_104),
.B1(n_14),
.B2(n_13),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_102),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_29),
.B(n_31),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_89),
.B(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_88),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_111),
.B1(n_92),
.B2(n_108),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_159),
.B1(n_122),
.B2(n_138),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_158),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_155),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_152),
.B1(n_156),
.B2(n_167),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_168),
.C(n_124),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_157),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_95),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_108),
.B1(n_91),
.B2(n_112),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_114),
.B1(n_105),
.B2(n_86),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_86),
.B1(n_105),
.B2(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_26),
.B1(n_14),
.B2(n_13),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_164),
.B(n_161),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_0),
.B(n_1),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_54),
.B1(n_26),
.B2(n_104),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_104),
.C(n_26),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_11),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_195),
.C(n_199),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_180),
.B(n_145),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_187),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_116),
.B(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_194),
.Y(n_219)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_146),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_167),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_135),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_200),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_119),
.C(n_132),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_145),
.A2(n_129),
.B1(n_123),
.B2(n_141),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_153),
.B1(n_152),
.B2(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_137),
.C(n_12),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_11),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_163),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_206),
.B1(n_173),
.B2(n_147),
.Y(n_222)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_172),
.C(n_154),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_221),
.C(n_199),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_180),
.B(n_192),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_164),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_169),
.B1(n_152),
.B2(n_166),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_193),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_247),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_177),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_235),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_233),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_224),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_182),
.B1(n_195),
.B2(n_203),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_196),
.B1(n_227),
.B2(n_214),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_178),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_200),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_239),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_223),
.C(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_202),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_204),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_248),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_191),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_191),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_258),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_218),
.B1(n_226),
.B2(n_229),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_260),
.B1(n_264),
.B2(n_245),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_225),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_261),
.C(n_236),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_229),
.B1(n_228),
.B2(n_220),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_225),
.C(n_198),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_183),
.B1(n_197),
.B2(n_190),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_185),
.B1(n_206),
.B2(n_197),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_235),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_272),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_219),
.B(n_190),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_276),
.B(n_7),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_250),
.C(n_262),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_253),
.B(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_248),
.B1(n_181),
.B2(n_230),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_181),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_279),
.Y(n_282)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_249),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_4),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_278),
.B1(n_266),
.B2(n_6),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_4),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_256),
.C(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_286),
.Y(n_291)
);

NAND4xp25_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_268),
.C(n_276),
.D(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_268),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_10),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_7),
.C(n_9),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_279),
.C(n_277),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_9),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_9),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_287),
.B1(n_289),
.B2(n_10),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_282),
.C(n_281),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_291),
.B(n_299),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_307),
.B(n_303),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_308),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_305),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_10),
.Y(n_314)
);


endmodule