module fake_jpeg_19865_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_22),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_52),
.B1(n_50),
.B2(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_55),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_50),
.B1(n_61),
.B2(n_65),
.Y(n_82)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_86),
.B1(n_51),
.B2(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_66),
.B1(n_76),
.B2(n_68),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_41),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_1),
.B(n_2),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_54),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_99),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_40),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_98),
.B(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_42),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_100),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_44),
.C(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_54),
.B(n_6),
.C(n_7),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_103),
.A3(n_102),
.B1(n_96),
.B2(n_90),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_109),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_112),
.B1(n_113),
.B2(n_105),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_105),
.B1(n_108),
.B2(n_104),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_5),
.C(n_8),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_9),
.A3(n_10),
.B1(n_14),
.B2(n_18),
.C1(n_19),
.C2(n_21),
.Y(n_118)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_24),
.A3(n_25),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_32),
.B(n_33),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_36),
.Y(n_121)
);


endmodule