module real_aes_9200_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g252 ( .A1(n_0), .A2(n_253), .B(n_254), .C(n_257), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_1), .B(n_241), .Y(n_258) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_3), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_4), .A2(n_130), .B(n_133), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_5), .A2(n_125), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_6), .A2(n_125), .B(n_235), .Y(n_234) );
AOI222xp33_ASAP7_75t_SL g113 ( .A1(n_7), .A2(n_61), .B1(n_114), .B2(n_720), .C1(n_721), .C2(n_725), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_8), .B(n_241), .Y(n_543) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_9), .A2(n_160), .B(n_197), .Y(n_196) );
AND2x6_ASAP7_75t_L g130 ( .A(n_10), .B(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_11), .A2(n_130), .B(n_133), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g481 ( .A(n_12), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_13), .B(n_39), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_14), .B(n_217), .Y(n_515) );
INVx1_ASAP7_75t_L g151 ( .A(n_15), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_16), .B(n_169), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_17), .A2(n_170), .B(n_499), .C(n_501), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_18), .B(n_241), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_19), .B(n_145), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_20), .A2(n_133), .B(n_136), .C(n_144), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_21), .A2(n_205), .B(n_256), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_22), .B(n_217), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_23), .B(n_217), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_24), .Y(n_528) );
INVx1_ASAP7_75t_L g453 ( .A(n_25), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_26), .A2(n_133), .B(n_144), .C(n_200), .Y(n_199) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_27), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_28), .Y(n_511) );
INVx1_ASAP7_75t_L g469 ( .A(n_29), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_30), .A2(n_125), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_32), .A2(n_173), .B(n_182), .C(n_184), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_33), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_34), .A2(n_256), .B(n_540), .C(n_542), .Y(n_539) );
INVxp67_ASAP7_75t_L g470 ( .A(n_35), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_36), .B(n_202), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_37), .A2(n_133), .B(n_144), .C(n_452), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g538 ( .A(n_38), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_40), .A2(n_257), .B(n_479), .C(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_41), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_42), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_43), .B(n_169), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_44), .B(n_125), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_45), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_46), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_47), .A2(n_173), .B(n_182), .C(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g255 ( .A(n_48), .Y(n_255) );
AOI222xp33_ASAP7_75t_SL g98 ( .A1(n_49), .A2(n_99), .B1(n_112), .B2(n_728), .C1(n_733), .C2(n_741), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_49), .A2(n_115), .B1(n_723), .B2(n_736), .Y(n_735) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_49), .Y(n_736) );
INVx1_ASAP7_75t_L g227 ( .A(n_50), .Y(n_227) );
INVx1_ASAP7_75t_L g487 ( .A(n_51), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_52), .B(n_125), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_53), .Y(n_153) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_54), .Y(n_477) );
INVx1_ASAP7_75t_L g131 ( .A(n_55), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_56), .B(n_125), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_57), .B(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_58), .A2(n_143), .B(n_166), .C(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_59), .Y(n_740) );
INVx1_ASAP7_75t_L g150 ( .A(n_60), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_61), .Y(n_720) );
INVx1_ASAP7_75t_SL g541 ( .A(n_62), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_63), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_64), .B(n_169), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_65), .B(n_241), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_66), .B(n_170), .Y(n_215) );
INVx1_ASAP7_75t_L g531 ( .A(n_67), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_68), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_69), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_70), .A2(n_133), .B(n_164), .C(n_173), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_71), .Y(n_236) );
INVx1_ASAP7_75t_L g103 ( .A(n_72), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_73), .A2(n_125), .B(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_74), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_75), .A2(n_125), .B(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_76), .A2(n_124), .B(n_465), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_77), .Y(n_450) );
INVx1_ASAP7_75t_L g497 ( .A(n_78), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_79), .B(n_141), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_80), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_81), .A2(n_125), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g500 ( .A(n_82), .Y(n_500) );
INVx2_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
INVx1_ASAP7_75t_L g514 ( .A(n_84), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_85), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_86), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_109), .Y(n_442) );
INVx2_ASAP7_75t_L g719 ( .A(n_87), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_88), .A2(n_133), .B(n_173), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_89), .B(n_125), .Y(n_180) );
INVx1_ASAP7_75t_L g185 ( .A(n_90), .Y(n_185) );
INVxp67_ASAP7_75t_L g239 ( .A(n_91), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_92), .B(n_160), .Y(n_482) );
INVx2_ASAP7_75t_L g490 ( .A(n_93), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_94), .B(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
INVx1_ASAP7_75t_L g211 ( .A(n_96), .Y(n_211) );
AND2x2_ASAP7_75t_L g229 ( .A(n_97), .B(n_147), .Y(n_229) );
INVx1_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_105), .Y(n_100) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g732 ( .A(n_102), .Y(n_732) );
INVx1_ASAP7_75t_L g731 ( .A(n_104), .Y(n_731) );
OA21x2_ASAP7_75t_L g742 ( .A1(n_104), .A2(n_732), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_107), .A2(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_SL g739 ( .A(n_107), .Y(n_739) );
BUFx2_ASAP7_75t_L g743 ( .A(n_107), .Y(n_743) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_108), .B(n_719), .Y(n_727) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g718 ( .A(n_109), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_440), .B1(n_443), .B2(n_716), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g723 ( .A(n_116), .Y(n_723) );
AND3x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_344), .C(n_401), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_289), .C(n_325), .Y(n_117) );
OAI211xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_191), .B(n_243), .C(n_276), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_155), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g246 ( .A(n_121), .B(n_247), .Y(n_246) );
INVx5_ASAP7_75t_L g275 ( .A(n_121), .Y(n_275) );
AND2x2_ASAP7_75t_L g348 ( .A(n_121), .B(n_264), .Y(n_348) );
AND2x2_ASAP7_75t_L g386 ( .A(n_121), .B(n_292), .Y(n_386) );
AND2x2_ASAP7_75t_L g406 ( .A(n_121), .B(n_248), .Y(n_406) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_152), .Y(n_121) );
AOI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_132), .B(n_145), .Y(n_122) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_126), .B(n_130), .Y(n_212) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g143 ( .A(n_127), .Y(n_143) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
INVx1_ASAP7_75t_L g206 ( .A(n_128), .Y(n_206) );
INVx1_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
INVx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx1_ASAP7_75t_L g202 ( .A(n_129), .Y(n_202) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_129), .Y(n_217) );
BUFx3_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
INVx4_ASAP7_75t_SL g174 ( .A(n_130), .Y(n_174) );
INVx5_ASAP7_75t_L g183 ( .A(n_133), .Y(n_183) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
BUFx3_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B(n_142), .Y(n_136) );
INVx2_ASAP7_75t_L g141 ( .A(n_138), .Y(n_141) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx4_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_141), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_141), .A2(n_187), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_141), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_141), .A2(n_516), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_142), .A2(n_169), .B(n_453), .C(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_143), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_146), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_147), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_147), .A2(n_224), .B(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_147), .A2(n_212), .B(n_450), .C(n_451), .Y(n_449) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_147), .A2(n_475), .B(n_482), .Y(n_474) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_L g161 ( .A(n_148), .B(n_149), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_154), .A2(n_510), .B(n_517), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_155), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_178), .Y(n_155) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_156), .Y(n_287) );
AND2x2_ASAP7_75t_L g301 ( .A(n_156), .B(n_247), .Y(n_301) );
INVx1_ASAP7_75t_L g324 ( .A(n_156), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_156), .B(n_275), .Y(n_363) );
OR2x2_ASAP7_75t_L g400 ( .A(n_156), .B(n_245), .Y(n_400) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_157), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_157), .B(n_248), .Y(n_343) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g264 ( .A(n_158), .B(n_248), .Y(n_264) );
BUFx2_ASAP7_75t_L g292 ( .A(n_158), .Y(n_292) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_176), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_159), .B(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_159), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_218), .Y(n_209) );
INVx3_ASAP7_75t_L g241 ( .A(n_159), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_159), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_159), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_159), .A2(n_527), .B(n_533), .Y(n_526) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_160), .A2(n_198), .B(n_199), .Y(n_197) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_175), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_168), .C(n_171), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_167), .A2(n_169), .B1(n_469), .B2(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_167), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_167), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_169), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g253 ( .A(n_169), .Y(n_253) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_170), .B(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g542 ( .A(n_172), .Y(n_542) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_174), .A2(n_183), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_174), .A2(n_183), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_174), .A2(n_183), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_174), .A2(n_183), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_174), .A2(n_183), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_174), .A2(n_183), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_174), .A2(n_183), .B(n_538), .C(n_539), .Y(n_537) );
INVx5_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
BUFx2_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
AND2x2_ASAP7_75t_L g425 ( .A(n_178), .B(n_279), .Y(n_425) );
OR2x6_ASAP7_75t_L g178 ( .A(n_179), .B(n_189), .Y(n_178) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g257 ( .A(n_188), .Y(n_257) );
INVx1_ASAP7_75t_L g501 ( .A(n_188), .Y(n_501) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_230), .Y(n_192) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_193), .A2(n_326), .B1(n_333), .B2(n_334), .C(n_337), .Y(n_325) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_207), .Y(n_193) );
AND2x2_ASAP7_75t_L g231 ( .A(n_194), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_194), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g260 ( .A(n_195), .B(n_208), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_195), .B(n_209), .Y(n_270) );
OR2x2_ASAP7_75t_L g281 ( .A(n_195), .B(n_232), .Y(n_281) );
AND2x2_ASAP7_75t_L g284 ( .A(n_195), .B(n_272), .Y(n_284) );
AND2x2_ASAP7_75t_L g300 ( .A(n_195), .B(n_221), .Y(n_300) );
OR2x2_ASAP7_75t_L g316 ( .A(n_195), .B(n_209), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_195), .B(n_232), .Y(n_378) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_196), .B(n_221), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_196), .B(n_209), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_203), .B(n_204), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g294 ( .A(n_207), .B(n_281), .Y(n_294) );
INVx2_ASAP7_75t_L g320 ( .A(n_207), .Y(n_320) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_221), .Y(n_207) );
AND2x2_ASAP7_75t_L g242 ( .A(n_208), .B(n_222), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_208), .B(n_232), .Y(n_299) );
OR2x2_ASAP7_75t_L g310 ( .A(n_208), .B(n_222), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_208), .B(n_272), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_208), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_402) );
INVx5_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_209), .B(n_232), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_212), .A2(n_511), .B(n_512), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_212), .A2(n_528), .B(n_529), .Y(n_527) );
INVx4_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
INVx2_ASAP7_75t_L g479 ( .A(n_217), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g462 ( .A(n_220), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_221), .B(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_221), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g288 ( .A(n_221), .B(n_260), .Y(n_288) );
OR2x2_ASAP7_75t_L g332 ( .A(n_221), .B(n_232), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_221), .B(n_284), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_221), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_221), .B(n_398), .Y(n_397) );
INVx5_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_222), .B(n_231), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_222), .A2(n_266), .B(n_269), .C(n_273), .Y(n_265) );
OR2x2_ASAP7_75t_L g303 ( .A(n_222), .B(n_299), .Y(n_303) );
OR2x2_ASAP7_75t_L g339 ( .A(n_222), .B(n_281), .Y(n_339) );
OAI311xp33_ASAP7_75t_L g345 ( .A1(n_222), .A2(n_284), .A3(n_346), .B1(n_349), .C1(n_356), .Y(n_345) );
AND2x2_ASAP7_75t_L g396 ( .A(n_222), .B(n_232), .Y(n_396) );
AND2x2_ASAP7_75t_L g404 ( .A(n_222), .B(n_259), .Y(n_404) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_222), .Y(n_422) );
AND2x2_ASAP7_75t_L g439 ( .A(n_222), .B(n_260), .Y(n_439) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_242), .Y(n_230) );
AND2x2_ASAP7_75t_L g267 ( .A(n_231), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g423 ( .A(n_231), .Y(n_423) );
AND2x2_ASAP7_75t_L g259 ( .A(n_232), .B(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g272 ( .A(n_232), .Y(n_272) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
INVxp67_ASAP7_75t_L g354 ( .A(n_232), .Y(n_354) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_240), .Y(n_232) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_233), .A2(n_485), .B(n_491), .Y(n_484) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_233), .A2(n_495), .B(n_502), .Y(n_494) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_233), .A2(n_536), .B(n_543), .Y(n_535) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_241), .A2(n_249), .B(n_258), .Y(n_248) );
AND2x2_ASAP7_75t_L g432 ( .A(n_242), .B(n_280), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_259), .B1(n_261), .B2(n_262), .C(n_265), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_245), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g285 ( .A(n_245), .B(n_275), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_245), .B(n_247), .Y(n_293) );
OR2x2_ASAP7_75t_L g305 ( .A(n_245), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g347 ( .A(n_245), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_245), .Y(n_367) );
AND2x2_ASAP7_75t_L g419 ( .A(n_245), .B(n_343), .Y(n_419) );
OAI31xp33_ASAP7_75t_L g427 ( .A1(n_245), .A2(n_296), .A3(n_395), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_246), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g391 ( .A(n_246), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_246), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g279 ( .A(n_247), .B(n_275), .Y(n_279) );
INVx1_ASAP7_75t_L g366 ( .A(n_247), .Y(n_366) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g416 ( .A(n_248), .B(n_275), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_256), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g516 ( .A(n_257), .Y(n_516) );
INVx1_ASAP7_75t_SL g426 ( .A(n_259), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_260), .B(n_331), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_261), .A2(n_373), .B1(n_411), .B2(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g274 ( .A(n_264), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g333 ( .A(n_264), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_264), .B(n_285), .Y(n_438) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g408 ( .A(n_267), .B(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_268), .A2(n_327), .B(n_329), .Y(n_326) );
OR2x2_ASAP7_75t_L g334 ( .A(n_268), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g355 ( .A(n_268), .B(n_343), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_268), .B(n_366), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_268), .B(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g382 ( .A1(n_269), .A2(n_383), .B1(n_388), .B2(n_391), .C(n_392), .Y(n_382) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OR2x2_ASAP7_75t_L g359 ( .A(n_270), .B(n_332), .Y(n_359) );
INVx1_ASAP7_75t_L g398 ( .A(n_270), .Y(n_398) );
INVx2_ASAP7_75t_L g374 ( .A(n_271), .Y(n_374) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_275), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g342 ( .A(n_275), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g430 ( .A(n_275), .B(n_400), .Y(n_430) );
AOI222xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B1(n_282), .B2(n_285), .C1(n_286), .C2(n_288), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_279), .B(n_287), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_279), .A2(n_329), .B1(n_357), .B2(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_279), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OAI21xp33_ASAP7_75t_SL g317 ( .A1(n_288), .A2(n_318), .B(n_321), .Y(n_317) );
OAI211xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_294), .B(n_295), .C(n_317), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_293), .A2(n_296), .B1(n_301), .B2(n_302), .C(n_304), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_293), .B(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g387 ( .A(n_293), .Y(n_387) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x2_ASAP7_75t_L g389 ( .A(n_298), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g306 ( .A(n_301), .Y(n_306) );
AND2x2_ASAP7_75t_L g312 ( .A(n_301), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_311), .B2(n_314), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_308), .B(n_320), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_309), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g409 ( .A(n_313), .Y(n_409) );
AND2x2_ASAP7_75t_L g428 ( .A(n_313), .B(n_343), .Y(n_428) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_320), .B(n_377), .Y(n_436) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_323), .B(n_391), .Y(n_434) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g357 ( .A(n_335), .Y(n_357) );
BUFx2_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
OAI21xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR3xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_360), .C(n_382), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_364), .B(n_368), .C(n_371), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_361), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp67_ASAP7_75t_SL g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_SL g390 ( .A(n_370), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B(n_379), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g395 ( .A(n_373), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B1(n_397), .B2(n_399), .Y(n_392) );
INVx2_ASAP7_75t_SL g413 ( .A(n_400), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_417), .C(n_429), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_413), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_418), .A2(n_430), .B(n_431), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_439), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g722 ( .A(n_441), .Y(n_722) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g724 ( .A(n_443), .Y(n_724) );
OR5x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_610), .C(n_674), .D(n_690), .E(n_705), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_544), .C(n_571), .D(n_594), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_492), .B(n_503), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_457), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_SL g523 ( .A(n_448), .Y(n_523) );
AND2x4_ASAP7_75t_L g557 ( .A(n_448), .B(n_546), .Y(n_557) );
OR2x2_ASAP7_75t_L g567 ( .A(n_448), .B(n_525), .Y(n_567) );
OR2x2_ASAP7_75t_L g613 ( .A(n_448), .B(n_460), .Y(n_613) );
AND2x2_ASAP7_75t_L g627 ( .A(n_448), .B(n_524), .Y(n_627) );
AND2x2_ASAP7_75t_L g670 ( .A(n_448), .B(n_560), .Y(n_670) );
AND2x2_ASAP7_75t_L g677 ( .A(n_448), .B(n_535), .Y(n_677) );
AND2x2_ASAP7_75t_L g696 ( .A(n_448), .B(n_586), .Y(n_696) );
AND2x2_ASAP7_75t_L g714 ( .A(n_448), .B(n_556), .Y(n_714) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
INVx1_ASAP7_75t_L g679 ( .A(n_457), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_473), .Y(n_457) );
AND2x2_ASAP7_75t_L g589 ( .A(n_458), .B(n_524), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_458), .B(n_609), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g622 ( .A1(n_458), .A2(n_623), .A3(n_626), .B1(n_628), .B2(n_632), .Y(n_622) );
AND2x2_ASAP7_75t_L g692 ( .A(n_458), .B(n_586), .Y(n_692) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g556 ( .A(n_460), .B(n_525), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_460), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g598 ( .A(n_460), .B(n_545), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_460), .B(n_677), .Y(n_676) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_471), .Y(n_460) );
INVx1_ASAP7_75t_L g561 ( .A(n_461), .Y(n_561) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_464), .A2(n_472), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_507), .Y(n_563) );
AND2x2_ASAP7_75t_L g639 ( .A(n_473), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g711 ( .A(n_473), .Y(n_711) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
OR2x2_ASAP7_75t_L g506 ( .A(n_474), .B(n_484), .Y(n_506) );
AND2x2_ASAP7_75t_L g520 ( .A(n_474), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_474), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g570 ( .A(n_474), .Y(n_570) );
AND2x2_ASAP7_75t_L g597 ( .A(n_474), .B(n_484), .Y(n_597) );
BUFx3_ASAP7_75t_L g600 ( .A(n_474), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_474), .B(n_575), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_474), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g551 ( .A(n_483), .Y(n_551) );
AND2x2_ASAP7_75t_L g569 ( .A(n_483), .B(n_549), .Y(n_569) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g580 ( .A(n_484), .B(n_494), .Y(n_580) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_484), .Y(n_593) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_493), .B(n_600), .Y(n_650) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g521 ( .A(n_494), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_494), .B(n_569), .C(n_570), .Y(n_568) );
OR2x2_ASAP7_75t_L g576 ( .A(n_494), .B(n_549), .Y(n_576) );
AND2x2_ASAP7_75t_L g596 ( .A(n_494), .B(n_549), .Y(n_596) );
AND2x2_ASAP7_75t_L g640 ( .A(n_494), .B(n_509), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_519), .B(n_522), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g715 ( .A(n_505), .B(n_640), .Y(n_715) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_506), .A2(n_613), .B1(n_655), .B2(n_657), .Y(n_654) );
OR2x2_ASAP7_75t_L g661 ( .A(n_506), .B(n_576), .Y(n_661) );
OR2x2_ASAP7_75t_L g685 ( .A(n_506), .B(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_506), .B(n_605), .Y(n_698) );
AND2x2_ASAP7_75t_L g591 ( .A(n_507), .B(n_592), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_507), .A2(n_664), .B(n_679), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g699 ( .A1(n_507), .A2(n_589), .A3(n_700), .B1(n_702), .B2(n_703), .Y(n_699) );
OR2x2_ASAP7_75t_L g710 ( .A(n_507), .B(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_508), .B(n_592), .Y(n_657) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
AND2x2_ASAP7_75t_L g615 ( .A(n_509), .B(n_580), .Y(n_615) );
AND3x2_ASAP7_75t_L g624 ( .A(n_509), .B(n_520), .C(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_521), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_521), .B(n_549), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g545 ( .A(n_523), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_523), .B(n_535), .Y(n_603) );
AND2x2_ASAP7_75t_L g621 ( .A(n_523), .B(n_525), .Y(n_621) );
OR2x2_ASAP7_75t_L g635 ( .A(n_523), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g681 ( .A(n_523), .B(n_609), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_524), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
AND2x2_ASAP7_75t_L g582 ( .A(n_525), .B(n_560), .Y(n_582) );
OR2x2_ASAP7_75t_L g636 ( .A(n_525), .B(n_560), .Y(n_636) );
AND2x2_ASAP7_75t_L g689 ( .A(n_525), .B(n_546), .Y(n_689) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g587 ( .A(n_526), .Y(n_587) );
AND2x2_ASAP7_75t_L g609 ( .A(n_526), .B(n_535), .Y(n_609) );
INVx2_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
INVx1_ASAP7_75t_L g566 ( .A(n_535), .Y(n_566) );
AOI211xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_552), .C(n_564), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_545), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g708 ( .A(n_545), .Y(n_708) );
AND2x2_ASAP7_75t_L g586 ( .A(n_546), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_549), .B(n_550), .Y(n_558) );
INVx1_ASAP7_75t_L g643 ( .A(n_549), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_549), .B(n_570), .Y(n_667) );
AND2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_597), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_550), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_558), .B1(n_559), .B2(n_562), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_555), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_556), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g581 ( .A(n_557), .B(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_SL g646 ( .A1(n_557), .A2(n_599), .B1(n_647), .B2(n_652), .C(n_654), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_557), .B(n_620), .Y(n_653) );
INVx1_ASAP7_75t_L g713 ( .A(n_559), .Y(n_713) );
BUFx3_ASAP7_75t_L g620 ( .A(n_560), .Y(n_620) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI21xp33_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_567), .B(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_566), .B(n_620), .Y(n_673) );
INVx1_ASAP7_75t_L g630 ( .A(n_567), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_567), .B(n_620), .Y(n_631) );
INVxp67_ASAP7_75t_L g651 ( .A(n_569), .Y(n_651) );
AND2x2_ASAP7_75t_L g592 ( .A(n_570), .B(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B(n_581), .C(n_583), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_SL g606 ( .A(n_574), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_606), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_575), .B(n_597), .Y(n_648) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_578), .A2(n_584), .B1(n_588), .B2(n_590), .Y(n_583) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g644 ( .A(n_580), .B(n_645), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_582), .A2(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_586), .A2(n_595), .B1(n_598), .B2(n_599), .C(n_601), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_586), .B(n_620), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_586), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g702 ( .A(n_592), .Y(n_702) );
INVxp67_ASAP7_75t_L g625 ( .A(n_593), .Y(n_625) );
INVx1_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g671 ( .A(n_596), .B(n_600), .Y(n_671) );
INVx1_ASAP7_75t_L g645 ( .A(n_600), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_600), .B(n_615), .Y(n_675) );
OAI32xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .A3(n_606), .B1(n_607), .B2(n_608), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g614 ( .A(n_609), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_609), .B(n_641), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_609), .B(n_670), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g709 ( .A(n_609), .B(n_620), .Y(n_709) );
NAND5xp2_ASAP7_75t_L g610 ( .A(n_611), .B(n_633), .C(n_646), .D(n_658), .E(n_659), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B1(n_616), .B2(n_618), .C(n_622), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp33_ASAP7_75t_SL g637 ( .A(n_617), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_620), .B(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_621), .A2(n_634), .B1(n_637), .B2(n_641), .Y(n_633) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI211xp5_ASAP7_75t_SL g628 ( .A1(n_624), .A2(n_629), .B(n_630), .C(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g656 ( .A(n_636), .Y(n_656) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_645), .B(n_694), .Y(n_704) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B1(n_664), .B2(n_668), .C1(n_671), .C2(n_672), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_678), .B2(n_680), .C(n_682), .Y(n_674) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_687), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g694 ( .A(n_686), .Y(n_694) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_695), .B2(n_697), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_710), .C(n_712), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_715), .Y(n_712) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_718), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
endmodule