module fake_netlist_6_3494_n_781 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_781);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_781;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_575;
wire n_368;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_772;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx3_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_42),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_26),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_53),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_30),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_71),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_46),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_35),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_65),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_44),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_75),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_22),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_24),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_110),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_28),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_7),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_74),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx4_ASAP7_75t_R g177 ( 
.A(n_68),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_92),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_27),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_50),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_80),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_14),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_51),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_45),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_34),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_66),
.Y(n_196)
);

BUFx8_ASAP7_75t_SL g197 ( 
.A(n_195),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_0),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_162),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_0),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_1),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_2),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_2),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_144),
.B(n_23),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_149),
.B(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_3),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_4),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_29),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_4),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_31),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_145),
.B(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_162),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_150),
.B(n_5),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

AOI22x1_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_192),
.B1(n_153),
.B2(n_189),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_155),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_190),
.B1(n_187),
.B2(n_154),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_175),
.B1(n_159),
.B2(n_186),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_173),
.B1(n_165),
.B2(n_183),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_158),
.Y(n_247)
);

BUFx6f_ASAP7_75t_SL g248 ( 
.A(n_214),
.Y(n_248)
);

AO22x2_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_178),
.B1(n_168),
.B2(n_182),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_190),
.B1(n_187),
.B2(n_181),
.Y(n_252)
);

OR2x6_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_9),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_224),
.B1(n_228),
.B2(n_215),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

NAND3x1_ASAP7_75t_L g259 ( 
.A(n_202),
.B(n_10),
.C(n_11),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_202),
.B(n_11),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_225),
.B(n_167),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_170),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_12),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_172),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_232),
.B1(n_235),
.B2(n_218),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_180),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_12),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_216),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_216),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_16),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_32),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_218),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_221),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_218),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_216),
.A2(n_21),
.B1(n_33),
.B2(n_36),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_38),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_47),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_198),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_231),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_219),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_231),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_219),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_245),
.B(n_219),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_219),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_226),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_242),
.A2(n_199),
.B(n_198),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_246),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_219),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_222),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_230),
.B(n_229),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_222),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_260),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_278),
.B(n_222),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_248),
.B(n_222),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_247),
.B(n_233),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_222),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_261),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_229),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_275),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_251),
.B(n_211),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_253),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_249),
.B(n_203),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_333),
.A2(n_261),
.B(n_277),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_334),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_287),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_293),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_233),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_249),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_317),
.A2(n_259),
.B(n_229),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_337),
.A2(n_259),
.B(n_253),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_327),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_249),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_301),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_233),
.Y(n_368)
);

OR2x6_ASAP7_75t_L g369 ( 
.A(n_320),
.B(n_250),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_250),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_250),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_320),
.B(n_253),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

BUFx4_ASAP7_75t_SL g378 ( 
.A(n_345),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_212),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_269),
.B1(n_201),
.B2(n_233),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_319),
.B(n_301),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_291),
.B(n_201),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_337),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_300),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_307),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_291),
.B(n_201),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_286),
.B(n_339),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_343),
.B(n_233),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_309),
.B(n_201),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_340),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_290),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_201),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_313),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_312),
.B(n_322),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_316),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_346),
.B(n_203),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_312),
.B(n_199),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_288),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_295),
.B(n_48),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_295),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_354),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_323),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_285),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_306),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_324),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_289),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_380),
.Y(n_423)
);

BUFx4f_ASAP7_75t_L g424 ( 
.A(n_413),
.Y(n_424)
);

CKINVDCx8_ASAP7_75t_R g425 ( 
.A(n_369),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_367),
.B(n_373),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_323),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_325),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_356),
.A2(n_390),
.B(n_382),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_373),
.B(n_325),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_349),
.B(n_347),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_373),
.B(n_292),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

OR2x6_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_294),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_378),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_350),
.B(n_197),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_296),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_197),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_299),
.Y(n_439)
);

OR2x6_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_299),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_353),
.B(n_302),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

CKINVDCx8_ASAP7_75t_R g444 ( 
.A(n_413),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_355),
.B(n_49),
.Y(n_445)
);

NAND2x1_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_52),
.Y(n_446)
);

NAND2x1p5_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_199),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_54),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_376),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_376),
.B(n_199),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_55),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_372),
.B(n_199),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_357),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_372),
.B(n_56),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_58),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_374),
.B(n_59),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_351),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_60),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_351),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_375),
.B(n_62),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_351),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_63),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_374),
.B(n_64),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_404),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

INVx8_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

BUFx12f_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_443),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_351),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_459),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

BUFx2_ASAP7_75t_SL g493 ( 
.A(n_465),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_468),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_357),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_468),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_419),
.Y(n_497)
);

INVx3_ASAP7_75t_SL g498 ( 
.A(n_467),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_422),
.Y(n_500)
);

BUFx24_ASAP7_75t_L g501 ( 
.A(n_460),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_424),
.B(n_462),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_351),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_460),
.B(n_375),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_441),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_429),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_449),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_426),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_426),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

CKINVDCx6p67_ASAP7_75t_R g521 ( 
.A(n_474),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_498),
.A2(n_358),
.B1(n_467),
.B2(n_360),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_498),
.A2(n_358),
.B1(n_467),
.B2(n_360),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_489),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_475),
.A2(n_418),
.B1(n_413),
.B2(n_423),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

BUFx2_ASAP7_75t_SL g530 ( 
.A(n_483),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_490),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_510),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_475),
.A2(n_413),
.B1(n_461),
.B2(n_452),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_501),
.A2(n_464),
.B1(n_363),
.B2(n_445),
.Y(n_537)
);

INVx8_ASAP7_75t_L g538 ( 
.A(n_499),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_498),
.A2(n_381),
.B1(n_444),
.B2(n_439),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_476),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_491),
.A2(n_381),
.B1(n_500),
.B2(n_512),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_500),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_512),
.A2(n_470),
.B1(n_458),
.B2(n_427),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_518),
.A2(n_445),
.B1(n_383),
.B2(n_464),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_483),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_499),
.B(n_359),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_509),
.A2(n_518),
.B1(n_484),
.B2(n_478),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_495),
.B(n_430),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_480),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_478),
.A2(n_484),
.B1(n_495),
.B2(n_480),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_516),
.A2(n_425),
.B1(n_469),
.B2(n_448),
.Y(n_551)
);

BUFx4_ASAP7_75t_SL g552 ( 
.A(n_497),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_478),
.A2(n_484),
.B1(n_480),
.B2(n_515),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_511),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_508),
.A2(n_402),
.B1(n_428),
.B2(n_427),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_481),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_505),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_499),
.B(n_359),
.Y(n_563)
);

CKINVDCx11_ASAP7_75t_R g564 ( 
.A(n_476),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_535),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_537),
.A2(n_431),
.B1(n_484),
.B2(n_478),
.Y(n_566)
);

AOI211xp5_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_409),
.B(n_352),
.C(n_416),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_549),
.A2(n_503),
.B1(n_479),
.B2(n_484),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_520),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_533),
.A2(n_430),
.B1(n_478),
.B2(n_448),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_551),
.A2(n_503),
.B1(n_479),
.B2(n_507),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_537),
.A2(n_352),
.B1(n_416),
.B2(n_480),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_544),
.A2(n_528),
.B1(n_525),
.B2(n_523),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_562),
.B(n_505),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_525),
.A2(n_432),
.B1(n_427),
.B2(n_428),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_L g577 ( 
.A1(n_542),
.A2(n_437),
.B(n_363),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_552),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_555),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_539),
.A2(n_432),
.B1(n_428),
.B2(n_437),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_507),
.B1(n_519),
.B2(n_434),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_552),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_559),
.A2(n_507),
.B1(n_469),
.B2(n_517),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_507),
.B1(n_519),
.B2(n_434),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_536),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_543),
.A2(n_507),
.B1(n_434),
.B2(n_397),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_560),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_556),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_561),
.A2(n_507),
.B1(n_527),
.B2(n_530),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_548),
.A2(n_507),
.B1(n_517),
.B2(n_485),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_524),
.A2(n_517),
.B1(n_485),
.B2(n_502),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_558),
.A2(n_359),
.B1(n_421),
.B2(n_410),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_550),
.B(n_486),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_532),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_541),
.A2(n_359),
.B1(n_421),
.B2(n_410),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_486),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_553),
.B(n_477),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_538),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_545),
.B(n_404),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_553),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_SL g605 ( 
.A1(n_522),
.A2(n_485),
.B1(n_502),
.B2(n_421),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_547),
.B(n_407),
.C(n_446),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_538),
.A2(n_502),
.B1(n_526),
.B2(n_534),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_521),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_553),
.A2(n_359),
.B1(n_361),
.B2(n_348),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_546),
.B(n_477),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_540),
.Y(n_612)
);

BUFx4f_ASAP7_75t_SL g613 ( 
.A(n_526),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_566),
.A2(n_494),
.B1(n_496),
.B2(n_504),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_600),
.B(n_506),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_574),
.A2(n_564),
.B1(n_450),
.B2(n_348),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_575),
.B(n_482),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_570),
.A2(n_534),
.B1(n_493),
.B2(n_563),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_573),
.A2(n_392),
.B1(n_389),
.B2(n_405),
.Y(n_619)
);

AO22x1_ASAP7_75t_L g620 ( 
.A1(n_578),
.A2(n_482),
.B1(n_492),
.B2(n_487),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_581),
.A2(n_504),
.B1(n_546),
.B2(n_563),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_571),
.A2(n_577),
.B1(n_567),
.B2(n_576),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_608),
.A2(n_392),
.B1(n_395),
.B2(n_405),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_608),
.A2(n_389),
.B1(n_395),
.B2(n_412),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_575),
.B(n_506),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_595),
.A2(n_493),
.B1(n_514),
.B2(n_442),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_594),
.A2(n_412),
.B1(n_406),
.B2(n_408),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_582),
.B(n_408),
.C(n_406),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_606),
.A2(n_412),
.B1(n_391),
.B2(n_400),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_591),
.A2(n_504),
.B1(n_487),
.B2(n_492),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_585),
.A2(n_492),
.B1(n_499),
.B2(n_506),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_595),
.A2(n_391),
.B1(n_393),
.B2(n_400),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_598),
.A2(n_391),
.B1(n_393),
.B2(n_400),
.Y(n_633)
);

OAI211xp5_ASAP7_75t_L g634 ( 
.A1(n_602),
.A2(n_442),
.B(n_456),
.C(n_514),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_597),
.B(n_513),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_596),
.A2(n_393),
.B1(n_386),
.B2(n_388),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_600),
.B(n_603),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_565),
.B(n_513),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_596),
.A2(n_386),
.B1(n_388),
.B2(n_412),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_568),
.A2(n_384),
.B1(n_394),
.B2(n_370),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_513),
.B1(n_361),
.B2(n_370),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_599),
.A2(n_384),
.B1(n_394),
.B2(n_388),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_612),
.A2(n_361),
.B1(n_370),
.B2(n_386),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_599),
.B(n_67),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_584),
.A2(n_390),
.B1(n_382),
.B2(n_403),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_390),
.B1(n_382),
.B2(n_399),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_565),
.B(n_379),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_593),
.A2(n_390),
.B1(n_382),
.B2(n_361),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_612),
.A2(n_379),
.B1(n_377),
.B2(n_371),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_588),
.B(n_69),
.Y(n_651)
);

OAI222xp33_ASAP7_75t_L g652 ( 
.A1(n_605),
.A2(n_377),
.B1(n_371),
.B2(n_447),
.C1(n_370),
.C2(n_79),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_637),
.B(n_586),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_586),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_648),
.B(n_589),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_615),
.B(n_589),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_644),
.B(n_569),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_625),
.B(n_572),
.Y(n_658)
);

OAI221xp5_ASAP7_75t_L g659 ( 
.A1(n_616),
.A2(n_583),
.B1(n_578),
.B2(n_609),
.C(n_607),
.Y(n_659)
);

OA211x2_ASAP7_75t_L g660 ( 
.A1(n_628),
.A2(n_613),
.B(n_583),
.C(n_604),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_609),
.C(n_604),
.Y(n_661)
);

AOI221xp5_ASAP7_75t_L g662 ( 
.A1(n_622),
.A2(n_580),
.B1(n_590),
.B2(n_579),
.C(n_611),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_626),
.B(n_611),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_619),
.B(n_579),
.C(n_601),
.Y(n_664)
);

AOI221xp5_ASAP7_75t_L g665 ( 
.A1(n_635),
.A2(n_652),
.B1(n_631),
.B2(n_617),
.C(n_623),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_651),
.B(n_601),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_638),
.B(n_604),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_618),
.B(n_610),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_636),
.B(n_70),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_643),
.A2(n_368),
.B1(n_447),
.B2(n_377),
.C(n_371),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_636),
.B(n_72),
.Y(n_671)
);

OAI221xp5_ASAP7_75t_L g672 ( 
.A1(n_640),
.A2(n_377),
.B1(n_371),
.B2(n_411),
.C(n_83),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_639),
.B(n_77),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_621),
.A2(n_411),
.B1(n_82),
.B2(n_84),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_620),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_650),
.B(n_78),
.C(n_85),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_639),
.B(n_86),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_646),
.B(n_87),
.Y(n_678)
);

OAI221xp5_ASAP7_75t_SL g679 ( 
.A1(n_649),
.A2(n_627),
.B1(n_645),
.B2(n_650),
.C(n_629),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_630),
.B(n_614),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_641),
.C(n_647),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_654),
.B(n_632),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_655),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_655),
.B(n_642),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_654),
.B(n_632),
.Y(n_685)
);

INVxp33_ASAP7_75t_SL g686 ( 
.A(n_675),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_653),
.B(n_88),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_658),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_672),
.B(n_624),
.C(n_633),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_658),
.B(n_633),
.Y(n_690)
);

AO21x1_ASAP7_75t_L g691 ( 
.A1(n_661),
.A2(n_89),
.B(n_90),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_656),
.B(n_93),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_667),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_657),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_663),
.B(n_94),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_657),
.B(n_95),
.Y(n_697)
);

AND4x1_ASAP7_75t_L g698 ( 
.A(n_662),
.B(n_96),
.C(n_98),
.D(n_99),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_688),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_688),
.B(n_663),
.Y(n_700)
);

XNOR2x2_ASAP7_75t_L g701 ( 
.A(n_697),
.B(n_686),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_695),
.Y(n_702)
);

XNOR2x2_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_680),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_695),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_683),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_694),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_693),
.B(n_666),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_686),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_684),
.Y(n_709)
);

XOR2x2_ASAP7_75t_L g710 ( 
.A(n_703),
.B(n_698),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

XNOR2x1_ASAP7_75t_L g712 ( 
.A(n_701),
.B(n_696),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_709),
.B(n_684),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_706),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_712),
.A2(n_708),
.B1(n_710),
.B2(n_713),
.Y(n_715)
);

OAI22x1_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_707),
.B1(n_708),
.B2(n_700),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_711),
.Y(n_717)
);

XOR2x2_ASAP7_75t_L g718 ( 
.A(n_711),
.B(n_696),
.Y(n_718)
);

AOI22x1_ASAP7_75t_L g719 ( 
.A1(n_710),
.A2(n_707),
.B1(n_692),
.B2(n_702),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_713),
.Y(n_720)
);

XNOR2xp5_ASAP7_75t_L g721 ( 
.A(n_715),
.B(n_666),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_720),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_718),
.A2(n_691),
.B1(n_681),
.B2(n_687),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

OAI322xp33_ASAP7_75t_L g726 ( 
.A1(n_724),
.A2(n_719),
.A3(n_717),
.B1(n_700),
.B2(n_705),
.C1(n_702),
.C2(n_704),
.Y(n_726)
);

CKINVDCx16_ASAP7_75t_R g727 ( 
.A(n_721),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_725),
.A2(n_722),
.B(n_717),
.C(n_689),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_727),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_727),
.A2(n_690),
.B1(n_674),
.B2(n_660),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_730),
.A2(n_729),
.B1(n_728),
.B2(n_731),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_SL g733 ( 
.A1(n_729),
.A2(n_691),
.B1(n_676),
.B2(n_664),
.Y(n_733)
);

OAI211xp5_ASAP7_75t_SL g734 ( 
.A1(n_729),
.A2(n_665),
.B(n_671),
.C(n_670),
.Y(n_734)
);

OA22x2_ASAP7_75t_L g735 ( 
.A1(n_730),
.A2(n_692),
.B1(n_704),
.B2(n_699),
.Y(n_735)
);

OA22x2_ASAP7_75t_L g736 ( 
.A1(n_730),
.A2(n_668),
.B1(n_678),
.B2(n_669),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_729),
.B(n_685),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_737),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_738),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_678),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_660),
.B1(n_668),
.B2(n_669),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_732),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_733),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_737),
.B(n_685),
.Y(n_746)
);

AND4x1_ASAP7_75t_L g747 ( 
.A(n_744),
.B(n_677),
.C(n_673),
.D(n_664),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_739),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_746),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

AND4x1_ASAP7_75t_L g753 ( 
.A(n_742),
.B(n_677),
.C(n_673),
.D(n_682),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_743),
.A2(n_679),
.B1(n_682),
.B2(n_102),
.Y(n_754)
);

AND4x1_ASAP7_75t_L g755 ( 
.A(n_744),
.B(n_100),
.C(n_101),
.D(n_103),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_752),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_749),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_748),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_751),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_754),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_750),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_747),
.B(n_109),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_754),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_757),
.Y(n_765)
);

NAND4xp25_ASAP7_75t_L g766 ( 
.A(n_764),
.B(n_753),
.C(n_112),
.D(n_113),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_763),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_756),
.A2(n_758),
.B1(n_759),
.B2(n_762),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_761),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_765),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_769),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_768),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_771),
.A2(n_766),
.B1(n_760),
.B2(n_767),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_773),
.A2(n_770),
.B1(n_123),
.B2(n_124),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_771),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_775),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_772),
.B1(n_776),
.B2(n_774),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_778),
.Y(n_779)
);

AOI221x1_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.C(n_131),
.Y(n_780)
);

AOI211xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_781)
);


endmodule