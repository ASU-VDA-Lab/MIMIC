module fake_jpeg_6942_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_18;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx3_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_5),
.C(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_7),
.Y(n_28)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_7),
.B(n_10),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_17),
.Y(n_33)
);

OR2x2_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_17),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_49),
.B(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_10),
.B1(n_13),
.B2(n_19),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_13),
.B1(n_19),
.B2(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_26),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_44),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_54),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_42),
.B(n_47),
.C(n_11),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_35),
.C(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_33),
.C(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_33),
.B1(n_54),
.B2(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_62),
.B1(n_50),
.B2(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_41),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.C(n_58),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_25),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_60),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_60),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_18),
.Y(n_72)
);


endmodule