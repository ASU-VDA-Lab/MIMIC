module fake_jpeg_22043_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_49),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_33),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_2),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_29),
.B1(n_24),
.B2(n_21),
.Y(n_50)
);

OA22x2_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_76),
.B1(n_59),
.B2(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_28),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_27),
.B1(n_34),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_30),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_29),
.B1(n_18),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_82),
.B1(n_55),
.B2(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_86),
.B1(n_3),
.B2(n_4),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_84),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_20),
.B1(n_35),
.B2(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_20),
.B1(n_17),
.B2(n_5),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_8),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_95),
.B1(n_101),
.B2(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_100),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_7),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_15),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_60),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_53),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_69),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_143),
.B1(n_92),
.B2(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_52),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_127),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_144),
.C(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_113),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_136),
.B(n_140),
.Y(n_156)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_104),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_89),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_89),
.A2(n_85),
.B1(n_75),
.B2(n_68),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_87),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_72),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_159),
.B(n_144),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_114),
.B(n_100),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_120),
.B(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_94),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_139),
.B1(n_138),
.B2(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_165),
.B1(n_144),
.B2(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_103),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_126),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_95),
.B1(n_102),
.B2(n_91),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_143),
.B1(n_55),
.B2(n_126),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_131),
.B1(n_126),
.B2(n_140),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_188),
.B1(n_161),
.B2(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_167),
.B1(n_172),
.B2(n_155),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_106),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_110),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_133),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_197),
.B(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_196),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_142),
.B(n_134),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_204),
.B(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_166),
.C(n_159),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_206),
.C(n_212),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_158),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_156),
.B(n_163),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_171),
.C(n_170),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_162),
.C(n_151),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_220),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_187),
.B1(n_189),
.B2(n_164),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_228),
.B1(n_209),
.B2(n_168),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_182),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_224),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_184),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_210),
.Y(n_238)
);

XOR2x1_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_197),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_206),
.C(n_198),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_237),
.C(n_227),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_222),
.B(n_185),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_212),
.C(n_213),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_243),
.B(n_245),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_238),
.C(n_225),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_222),
.B(n_205),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_182),
.B1(n_216),
.B2(n_172),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_252),
.B1(n_229),
.B2(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_155),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_250),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_231),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_225),
.B(n_195),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_243),
.B1(n_249),
.B2(n_252),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_259),
.B(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_148),
.Y(n_260)
);

AOI321xp33_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_255),
.A3(n_176),
.B1(n_66),
.B2(n_14),
.C(n_13),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_93),
.C(n_10),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_261),
.Y(n_264)
);


endmodule