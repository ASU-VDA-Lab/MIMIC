module real_jpeg_32710_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_712, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_712;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_704;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_707;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_703;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_699;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_708;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_694;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_0),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_0),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_1),
.A2(n_370),
.B1(n_371),
.B2(n_373),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_1),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_1),
.A2(n_370),
.B1(n_464),
.B2(n_466),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_1),
.A2(n_370),
.B1(n_578),
.B2(n_582),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_1),
.A2(n_370),
.B1(n_616),
.B2(n_618),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_183),
.B1(n_189),
.B2(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_2),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_2),
.A2(n_102),
.B1(n_189),
.B2(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_2),
.A2(n_189),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_2),
.A2(n_189),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_4),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_176),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_4),
.A2(n_176),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_4),
.A2(n_176),
.B1(n_354),
.B2(n_358),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_5),
.A2(n_178),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_5),
.Y(n_266)
);

OAI22x1_ASAP7_75t_SL g380 ( 
.A1(n_5),
.A2(n_266),
.B1(n_381),
.B2(n_384),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_5),
.A2(n_266),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_5),
.A2(n_266),
.B1(n_540),
.B2(n_542),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_7),
.A2(n_24),
.B1(n_123),
.B2(n_127),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_24),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_7),
.A2(n_24),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_9),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_10),
.A2(n_65),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_10),
.A2(n_195),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_10),
.A2(n_195),
.B1(n_311),
.B2(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_10),
.A2(n_195),
.B1(n_508),
.B2(n_511),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_11),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_11),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_11),
.B(n_71),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_11),
.B(n_546),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_11),
.A2(n_477),
.B1(n_569),
.B2(n_572),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_11),
.B(n_83),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_L g624 ( 
.A1(n_11),
.A2(n_301),
.B(n_604),
.Y(n_624)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_14),
.B1(n_20),
.B2(n_708),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_14),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_63),
.B1(n_101),
.B2(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_15),
.A2(n_63),
.B1(n_161),
.B2(n_166),
.Y(n_160)
);

AO22x1_ASAP7_75t_SL g239 ( 
.A1(n_15),
.A2(n_63),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_16),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_16),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_17),
.A2(n_29),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_17),
.A2(n_323),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_17),
.A2(n_323),
.B1(n_529),
.B2(n_533),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_17),
.A2(n_323),
.B1(n_597),
.B2(n_602),
.Y(n_596)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_18),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_74),
.B(n_705),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_72),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_22),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_22),
.B(n_222),
.Y(n_704)
);

CKINVDCx14_ASAP7_75t_R g707 ( 
.A(n_22),
.Y(n_707)
);

AOI22x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_62),
.B2(n_70),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_23),
.A2(n_34),
.B1(n_70),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_28),
.Y(n_180)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_28),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_28),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_28),
.Y(n_374)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_32),
.Y(n_325)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_32),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_33),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_62),
.B(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_34),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_35),
.A2(n_70),
.B1(n_182),
.B2(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_35),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_35),
.B(n_322),
.Y(n_321)
);

AO22x1_ASAP7_75t_SL g368 ( 
.A1(n_35),
.A2(n_71),
.B1(n_322),
.B2(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_35),
.B(n_472),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_50),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_44),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_44),
.Y(n_432)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_46),
.Y(n_265)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_57),
.B2(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_55),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_55),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_56),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_56),
.Y(n_429)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_59),
.Y(n_571)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_67),
.Y(n_420)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_71),
.B(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_71),
.B(n_262),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_71),
.B(n_369),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_73),
.B(n_707),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_344),
.B(n_694),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_223),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_220),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_78),
.B(n_221),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_210),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_79),
.B(n_210),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_193),
.C(n_200),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_80),
.A2(n_193),
.B1(n_202),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_80),
.Y(n_339)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_169),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_131),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_82),
.B(n_212),
.C(n_213),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_100),
.B1(n_110),
.B2(n_122),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_83),
.A2(n_110),
.B1(n_122),
.B2(n_204),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g215 ( 
.A1(n_83),
.A2(n_100),
.B(n_110),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_83),
.A2(n_110),
.B1(n_204),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_83),
.A2(n_110),
.B1(n_279),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_83),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_83),
.B(n_380),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_83),
.A2(n_110),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_111),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_96),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_87),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_88),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_95),
.Y(n_560)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_105),
.Y(n_417)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_108),
.Y(n_334)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_110),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_110),
.B(n_380),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_125),
.Y(n_383)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_126),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_126),
.Y(n_409)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_130),
.Y(n_556)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_130),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_131),
.B(n_202),
.C(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_131),
.B(n_203),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_160),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_133),
.A2(n_151),
.B1(n_245),
.B2(n_252),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_133),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_133),
.A2(n_151),
.B1(n_245),
.B2(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_133),
.A2(n_151),
.B1(n_308),
.B2(n_364),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_133),
.A2(n_151),
.B1(n_528),
.B2(n_577),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_133),
.A2(n_577),
.B(n_592),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_133),
.B(n_477),
.Y(n_613)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_134),
.A2(n_276),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_134),
.B(n_482),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_152),
.Y(n_151)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_143),
.B2(n_147),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_136),
.Y(n_300)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_137),
.Y(n_441)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_138),
.Y(n_357)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_138),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_138),
.Y(n_646)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_145),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_148),
.Y(n_543)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_SL g527 ( 
.A1(n_151),
.A2(n_528),
.B(n_534),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_154),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_158),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_159),
.Y(n_532)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_159),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_160),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_165),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_168),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_181),
.B2(n_192),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_173),
.Y(n_425)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_175),
.Y(n_476)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_193),
.B(n_273),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_193),
.B(n_286),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_193),
.A2(n_202),
.B1(n_270),
.B2(n_271),
.Y(n_341)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_201),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_202),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_202),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_209),
.Y(n_465)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_209),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_216),
.C(n_218),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_220),
.B(n_699),
.Y(n_698)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_336),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_288),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g703 ( 
.A(n_226),
.B(n_288),
.Y(n_703)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_268),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_227),
.B(n_341),
.C(n_342),
.Y(n_340)
);

OA21x2_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_258),
.B(n_259),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_244),
.Y(n_228)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_260),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_229),
.A2(n_244),
.B1(n_258),
.B2(n_391),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_236),
.B(n_239),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_230),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_230),
.A2(n_353),
.B1(n_434),
.B2(n_437),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_230),
.B(n_539),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_230),
.A2(n_636),
.B1(n_637),
.B2(n_638),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_232),
.Y(n_359)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_232),
.Y(n_443)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_233),
.Y(n_512)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_233),
.Y(n_661)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_235),
.Y(n_606)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_237),
.A2(n_301),
.B1(n_438),
.B2(n_507),
.Y(n_506)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_238),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_242),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_242),
.Y(n_617)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_244),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_249),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_249),
.Y(n_666)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_251),
.Y(n_484)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_251),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_252),
.Y(n_277)
);

BUFx6f_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_261),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_284),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_283),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_271),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

OA21x2_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_274),
.B(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_276),
.B(n_482),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_276),
.B(n_669),
.Y(n_668)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_294),
.B(n_335),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_R g335 ( 
.A(n_290),
.B(n_291),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_290),
.B(n_292),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_294),
.B(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_317),
.C(n_326),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_295),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_307),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_296),
.B(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_301),
.B(n_302),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_297),
.A2(n_301),
.B1(n_352),
.B2(n_360),
.Y(n_351)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_301),
.A2(n_596),
.B(n_604),
.Y(n_595)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_303),
.Y(n_537)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_306),
.Y(n_436)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_306),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_307),
.Y(n_446)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_313),
.Y(n_533)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_315),
.Y(n_656)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_328),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_320),
.B(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_336),
.B(n_703),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_337),
.B(n_340),
.Y(n_696)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_515),
.B(n_685),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_451),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_347),
.A2(n_686),
.B(n_690),
.Y(n_685)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_395),
.B(n_397),
.Y(n_347)
);

NOR2x1_ASAP7_75t_SL g691 ( 
.A(n_348),
.B(n_395),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_348),
.B(n_395),
.Y(n_693)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_389),
.C(n_392),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_399),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_368),
.C(n_375),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_363),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_351),
.B(n_363),
.Y(n_489)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_354),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g541 ( 
.A(n_357),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx4f_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_368),
.B(n_376),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_379),
.B2(n_388),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_377),
.A2(n_504),
.B(n_505),
.Y(n_503)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_407),
.B(n_412),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_388),
.A2(n_412),
.B(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_393),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_398),
.B(n_400),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_447),
.B(n_450),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_444),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_402),
.B(n_444),
.Y(n_450)
);

XOR2x1_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.C(n_413),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_404),
.B1(n_406),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_456),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_433),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_414),
.B(n_433),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_418),
.B1(n_424),
.B2(n_426),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_424),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_453),
.A2(n_490),
.B(n_493),
.Y(n_452)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_453),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.C(n_489),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_454),
.A2(n_455),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_489),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_470),
.C(n_479),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_461),
.B(n_480),
.Y(n_499)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_463),
.Y(n_504)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_470),
.B(n_499),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_477),
.B(n_478),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_477),
.B(n_553),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_627),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_477),
.B(n_654),
.Y(n_653)
);

OAI21xp33_ASAP7_75t_SL g669 ( 
.A1(n_477),
.A2(n_653),
.B(n_670),
.Y(n_669)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_490),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_497),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_494),
.B(n_497),
.Y(n_687)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.C(n_501),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_518),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.C(n_513),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_503),
.B(n_524),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_513),
.B1(n_514),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_506),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_507),
.A2(n_537),
.B(n_538),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_510),
.Y(n_632)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_561),
.B(n_683),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_517),
.Y(n_684)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_521),
.B(n_684),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_526),
.C(n_535),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_564),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_526),
.A2(n_527),
.B1(n_535),
.B2(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_534),
.B(n_668),
.Y(n_667)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_535),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_544),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g586 ( 
.A(n_536),
.B(n_544),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_538),
.A2(n_615),
.B(n_619),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_539),
.B(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_545),
.A2(n_549),
.B1(n_552),
.B2(n_555),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_554),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_557),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

AO21x2_ASAP7_75t_L g561 ( 
.A1(n_562),
.A2(n_587),
.B(n_682),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_563),
.B(n_566),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_563),
.B(n_566),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_575),
.C(n_585),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_576),
.Y(n_609)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx3_ASAP7_75t_SL g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_586),
.B1(n_608),
.B2(n_609),
.Y(n_607)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

OAI321xp33_ASAP7_75t_L g587 ( 
.A1(n_588),
.A2(n_610),
.A3(n_674),
.B1(n_680),
.B2(n_681),
.C(n_712),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_607),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_607),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_593),
.C(n_595),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_591),
.A2(n_593),
.B1(n_594),
.B2(n_679),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_595),
.Y(n_677)
);

INVxp33_ASAP7_75t_SL g636 ( 
.A(n_596),
.Y(n_636)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_599),
.Y(n_618)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_611),
.A2(n_634),
.B(n_673),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_612),
.A2(n_623),
.B(n_633),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_614),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_613),
.B(n_614),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_615),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_617),
.Y(n_616)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_622),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_624),
.B(n_625),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_626),
.B(n_631),
.Y(n_625)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_639),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_635),
.B(n_639),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_640),
.B(n_667),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_640),
.B(n_667),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_641),
.A2(n_652),
.B1(n_657),
.B2(n_662),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_642),
.B(n_647),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_663),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

BUFx4f_ASAP7_75t_SL g670 ( 
.A(n_671),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_675),
.B(n_676),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_675),
.B(n_676),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_677),
.B(n_678),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_687),
.B(n_688),
.C(n_689),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_691),
.A2(n_692),
.B(n_693),
.Y(n_690)
);

NOR2x1_ASAP7_75t_L g694 ( 
.A(n_695),
.B(n_700),
.Y(n_694)
);

AO21x1_ASAP7_75t_L g695 ( 
.A1(n_696),
.A2(n_697),
.B(n_698),
.Y(n_695)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_697),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_701),
.A2(n_702),
.B(n_704),
.Y(n_700)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_706),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_709),
.Y(n_708)
);

BUFx12_ASAP7_75t_L g709 ( 
.A(n_710),
.Y(n_709)
);


endmodule