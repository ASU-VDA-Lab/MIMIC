module fake_jpeg_21967_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx8_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_19),
.B1(n_16),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_22),
.C(n_27),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_24),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_48),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_37),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_13),
.B1(n_19),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_39),
.B1(n_47),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_30),
.B1(n_17),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_58),
.B1(n_62),
.B2(n_65),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_67),
.B(n_10),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_10),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_10),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_6),
.B(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_76),
.B1(n_65),
.B2(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_63),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_54),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.C(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_58),
.B1(n_56),
.B2(n_62),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_58),
.C(n_57),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_65),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_74),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_53),
.B1(n_67),
.B2(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_67),
.B1(n_68),
.B2(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_83),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_107),
.C(n_94),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_82),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_108),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_82),
.C(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_106),
.A2(n_87),
.B1(n_97),
.B2(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_104),
.B1(n_105),
.B2(n_100),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_113),
.C(n_116),
.Y(n_120)
);

XOR2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_97),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_107),
.B(n_105),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_93),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_102),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.C(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_108),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_103),
.A3(n_104),
.B1(n_122),
.B2(n_118),
.C1(n_111),
.C2(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_92),
.A3(n_101),
.B1(n_116),
.B2(n_117),
.C1(n_122),
.C2(n_128),
.Y(n_130)
);


endmodule