module fake_jpeg_10792_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_566;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_22),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_22),
.B(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_67),
.B(n_107),
.Y(n_150)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_31),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_34),
.B1(n_38),
.B2(n_19),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_33),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_45),
.Y(n_151)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_19),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_100),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_30),
.B(n_2),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_47),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_4),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_52),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_111),
.B(n_120),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_123),
.A2(n_149),
.B1(n_52),
.B2(n_8),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_160),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_54),
.B1(n_29),
.B2(n_45),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_76),
.B1(n_90),
.B2(n_63),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_56),
.B(n_38),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_137),
.B(n_172),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_40),
.B1(n_23),
.B2(n_54),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_151),
.Y(n_199)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_69),
.B(n_53),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_57),
.A2(n_62),
.B1(n_60),
.B2(n_66),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_163),
.A2(n_168),
.B1(n_102),
.B2(n_99),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_68),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_176),
.Y(n_206)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_72),
.A2(n_40),
.B1(n_45),
.B2(n_51),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_75),
.B(n_41),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_96),
.B(n_41),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_91),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_100),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_177),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_214),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_51),
.B1(n_53),
.B2(n_48),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_179),
.A2(n_187),
.B1(n_220),
.B2(n_234),
.Y(n_247)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_180),
.Y(n_289)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_182),
.Y(n_280)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_184),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_205),
.Y(n_250)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_186),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_34),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_189),
.B(n_196),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_61),
.B(n_44),
.C(n_43),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_190),
.A2(n_207),
.B(n_218),
.Y(n_258)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

OR2x4_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_85),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_193),
.B(n_225),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_4),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_198),
.Y(n_294)
);

OR2x2_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_90),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_200),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_126),
.B(n_47),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_201),
.B(n_232),
.C(n_158),
.Y(n_267)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_203),
.Y(n_291)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

BUFx16f_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_104),
.B1(n_103),
.B2(n_47),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_113),
.B(n_33),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_209),
.B(n_221),
.Y(n_273)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_210),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_224),
.B1(n_230),
.B2(n_207),
.Y(n_246)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_215),
.Y(n_251)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_217),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_163),
.A2(n_170),
.B1(n_112),
.B2(n_135),
.Y(n_218)
);

CKINVDCx12_ASAP7_75t_R g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_115),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_5),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_140),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_223),
.Y(n_265)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_112),
.A2(n_47),
.B1(n_33),
.B2(n_84),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_47),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_5),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_231),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_131),
.A2(n_92),
.B1(n_86),
.B2(n_79),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_144),
.B(n_5),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_235),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_114),
.A2(n_132),
.B1(n_173),
.B2(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_114),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_132),
.B(n_6),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_239),
.Y(n_259)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_114),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_235),
.B1(n_216),
.B2(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_142),
.B(n_7),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_142),
.B1(n_124),
.B2(n_162),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_241),
.A2(n_249),
.B1(n_256),
.B2(n_264),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_147),
.C(n_139),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g338 ( 
.A(n_243),
.B(n_267),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_246),
.A2(n_284),
.B1(n_271),
.B2(n_288),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_124),
.B1(n_159),
.B2(n_117),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_193),
.B(n_147),
.CI(n_8),
.CON(n_255),
.SN(n_255)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_255),
.B(n_290),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_199),
.B1(n_218),
.B2(n_202),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_115),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_270),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_178),
.A2(n_117),
.B1(n_158),
.B2(n_154),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_263),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_232),
.A2(n_159),
.B1(n_154),
.B2(n_148),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_268),
.A2(n_243),
.B(n_247),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_148),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_130),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_275),
.B(n_285),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_178),
.B(n_129),
.C(n_130),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_288),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_205),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_190),
.A2(n_129),
.B1(n_52),
.B2(n_11),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_282),
.B1(n_292),
.B2(n_233),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_230),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_213),
.A2(n_180),
.B1(n_192),
.B2(n_214),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_224),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_201),
.B(n_12),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_12),
.C(n_13),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_SL g290 ( 
.A(n_238),
.B(n_13),
.C(n_14),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_181),
.A2(n_13),
.B1(n_14),
.B2(n_191),
.Y(n_292)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_301),
.A2(n_318),
.B1(n_322),
.B2(n_336),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_229),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_303),
.B(n_319),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_231),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_305),
.Y(n_350)
);

INVx2_ASAP7_75t_R g305 ( 
.A(n_257),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_195),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_323),
.B(n_341),
.Y(n_362)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_317),
.Y(n_347)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_310),
.Y(n_374)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_311),
.Y(n_382)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_251),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_258),
.A2(n_208),
.B1(n_182),
.B2(n_204),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_252),
.B(n_223),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_328),
.Y(n_356)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_258),
.A2(n_220),
.B1(n_197),
.B2(n_188),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_183),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_324),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_261),
.B(n_222),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_325),
.B(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_186),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_14),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_340),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_205),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_14),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_330),
.B(n_331),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_250),
.B(n_270),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_333),
.B(n_342),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_334),
.A2(n_281),
.B(n_244),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_335),
.A2(n_277),
.B1(n_264),
.B2(n_290),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_249),
.A2(n_241),
.B1(n_268),
.B2(n_271),
.Y(n_336)
);

INVx13_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_245),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_345),
.Y(n_358)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_244),
.A2(n_255),
.B(n_285),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_262),
.B(n_244),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_343),
.Y(n_359)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_344),
.B(n_286),
.Y(n_363)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_245),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g411 ( 
.A1(n_346),
.A2(n_383),
.B(n_388),
.C(n_328),
.D(n_296),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_353),
.A2(n_296),
.B1(n_301),
.B2(n_313),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_298),
.A2(n_279),
.B(n_274),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_354),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_294),
.C(n_265),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_367),
.C(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_369),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_294),
.C(n_265),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_304),
.B(n_274),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_300),
.A2(n_284),
.B1(n_286),
.B2(n_282),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_371),
.A2(n_323),
.B1(n_298),
.B2(n_341),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_335),
.A2(n_280),
.B1(n_253),
.B2(n_276),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_336),
.B1(n_313),
.B2(n_322),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_297),
.Y(n_373)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_307),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_299),
.B(n_265),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_376),
.B(n_316),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_295),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_334),
.A2(n_276),
.B(n_278),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_381),
.B(n_314),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_306),
.A2(n_295),
.B(n_278),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_299),
.B(n_289),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_387),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_305),
.B(n_316),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_306),
.A2(n_323),
.B(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_391),
.A2(n_403),
.B1(n_412),
.B2(n_418),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_315),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_396),
.C(n_398),
.Y(n_433)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_394),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_395),
.A2(n_420),
.B1(n_362),
.B2(n_388),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_315),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_369),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_414),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_332),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_400),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_364),
.A2(n_342),
.B1(n_309),
.B2(n_327),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_401),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_347),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_402),
.B(n_407),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_305),
.Y(n_404)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_421),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_411),
.B(n_423),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_344),
.B1(n_333),
.B2(n_340),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_363),
.Y(n_414)
);

CKINVDCx12_ASAP7_75t_R g415 ( 
.A(n_367),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_415),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_373),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_425),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_312),
.C(n_324),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_383),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_329),
.B1(n_345),
.B2(n_339),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_379),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_419),
.B(n_422),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_371),
.A2(n_376),
.B1(n_356),
.B2(n_354),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_379),
.B(n_321),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_329),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_352),
.B(n_310),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_350),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_375),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_431),
.A2(n_454),
.B1(n_450),
.B2(n_428),
.Y(n_462)
);

OA22x2_ASAP7_75t_L g432 ( 
.A1(n_397),
.A2(n_381),
.B1(n_346),
.B2(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_432),
.B(n_409),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_440),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_366),
.Y(n_439)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_387),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_410),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_441),
.B(n_451),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_352),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_458),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_359),
.Y(n_444)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_444),
.Y(n_480)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_404),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_350),
.Y(n_456)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_362),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_SL g459 ( 
.A(n_452),
.B(n_411),
.C(n_389),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_460),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_357),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_406),
.C(n_417),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_471),
.C(n_476),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_462),
.B(n_472),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_464),
.B(n_466),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_414),
.Y(n_465)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_457),
.A2(n_420),
.B1(n_409),
.B2(n_403),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_425),
.Y(n_467)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_470),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_406),
.C(n_412),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_427),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_437),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_434),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_355),
.C(n_380),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_431),
.A2(n_391),
.B1(n_418),
.B2(n_416),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_477),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_360),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_482),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_380),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_465),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_405),
.B1(n_370),
.B2(n_351),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_487),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_SL g486 ( 
.A(n_426),
.B(n_370),
.C(n_410),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_426),
.B(n_444),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_442),
.A2(n_385),
.B1(n_394),
.B2(n_355),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_488),
.A2(n_511),
.B(n_467),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_491),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_443),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_435),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_505),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_440),
.C(n_430),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_495),
.B(n_496),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_455),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_509),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_432),
.C(n_442),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_500),
.B(n_501),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_432),
.C(n_449),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_432),
.C(n_448),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_478),
.C(n_487),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_SL g505 ( 
.A(n_466),
.B(n_365),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_365),
.Y(n_508)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_508),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_481),
.B(n_453),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_464),
.A2(n_446),
.B1(n_436),
.B2(n_429),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_500),
.B(n_470),
.CI(n_501),
.CON(n_513),
.SN(n_513)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_523),
.Y(n_532)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_515),
.Y(n_542)
);

AOI321xp33_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_459),
.A3(n_480),
.B1(n_485),
.B2(n_478),
.C(n_486),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_516),
.Y(n_543)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_519),
.Y(n_545)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_521),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_482),
.C(n_483),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_527),
.C(n_507),
.Y(n_533)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_511),
.Y(n_523)
);

INVx13_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_528),
.B1(n_529),
.B2(n_468),
.Y(n_539)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_510),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_525),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_488),
.A2(n_485),
.B(n_479),
.C(n_469),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_503),
.B(n_519),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_527),
.B(n_513),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_539),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_498),
.C(n_494),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_535),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_495),
.C(n_492),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_525),
.A2(n_490),
.B1(n_504),
.B2(n_505),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_537),
.A2(n_540),
.B1(n_527),
.B2(n_513),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_516),
.A2(n_504),
.B1(n_507),
.B2(n_468),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_512),
.A2(n_530),
.B1(n_515),
.B2(n_526),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_541),
.B(n_544),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_524),
.A2(n_469),
.B1(n_463),
.B2(n_504),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_509),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_436),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_514),
.C(n_518),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_548),
.A2(n_549),
.B(n_555),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_514),
.C(n_527),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_557),
.Y(n_559)
);

OAI21x1_ASAP7_75t_SL g564 ( 
.A1(n_553),
.A2(n_537),
.B(n_546),
.Y(n_564)
);

BUFx12f_ASAP7_75t_SL g554 ( 
.A(n_543),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_554),
.B(n_545),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_532),
.A2(n_365),
.B(n_463),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_446),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_558),
.C(n_531),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_385),
.C(n_429),
.Y(n_558)
);

FAx1_ASAP7_75t_SL g560 ( 
.A(n_549),
.B(n_548),
.CI(n_550),
.CON(n_560),
.SN(n_560)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_562),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_542),
.C(n_540),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_552),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_564),
.A2(n_558),
.B1(n_557),
.B2(n_536),
.Y(n_568)
);

AOI322xp5_ASAP7_75t_L g566 ( 
.A1(n_565),
.A2(n_554),
.A3(n_536),
.B1(n_427),
.B2(n_311),
.C1(n_556),
.C2(n_552),
.Y(n_566)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_566),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_567),
.A2(n_563),
.B(n_560),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_568),
.B(n_561),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_570),
.B(n_569),
.C(n_567),
.Y(n_573)
);

AOI322xp5_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_559),
.A3(n_337),
.B1(n_368),
.B2(n_349),
.C1(n_382),
.C2(n_374),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_573),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_571),
.C(n_574),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_374),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_368),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g579 ( 
.A(n_578),
.B(n_382),
.CI(n_337),
.CON(n_579),
.SN(n_579)
);


endmodule