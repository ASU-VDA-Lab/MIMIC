module fake_ariane_300_n_967 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_967);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_967;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx11_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_48),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_57),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_21),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_125),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_35),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_65),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_52),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_83),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_104),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_87),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_20),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_97),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_46),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_68),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_121),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_17),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_106),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_24),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_81),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_78),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_164),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_187),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_82),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_16),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_5),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_189),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_92),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_193),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_130),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_29),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_51),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_10),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_41),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_128),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_115),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_182),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_40),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_77),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_199),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_199),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_204),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_219),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_219),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_202),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_209),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_205),
.B(n_0),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_236),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_238),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_198),
.B(n_0),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_257),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_206),
.B(n_2),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_266),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_198),
.B(n_2),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_196),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_197),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_211),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_221),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_201),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_214),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_257),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_203),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_227),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_216),
.B(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_223),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_287),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_283),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_R g335 ( 
.A(n_280),
.B(n_212),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_250),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_278),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_319),
.B(n_230),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_R g345 ( 
.A(n_297),
.B(n_213),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_319),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_224),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_258),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_298),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_322),
.B(n_230),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_282),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_290),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_258),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_239),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_305),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_246),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_307),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_310),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_272),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_292),
.A2(n_253),
.B(n_251),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_300),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_311),
.B(n_230),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_304),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_311),
.B1(n_326),
.B2(n_290),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_380),
.B(n_263),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_320),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_281),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

OR2x6_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_285),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_331),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_320),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_286),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_365),
.A2(n_259),
.B1(n_325),
.B2(n_288),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_343),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_336),
.B(n_272),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_330),
.Y(n_403)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_370),
.B(n_259),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_336),
.B(n_242),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_336),
.A2(n_303),
.B1(n_256),
.B2(n_270),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_375),
.B(n_370),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_348),
.B(n_269),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_376),
.B(n_342),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_247),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_352),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_237),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

BUFx8_ASAP7_75t_SL g420 ( 
.A(n_363),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_260),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_303),
.B1(n_274),
.B2(n_275),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_241),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_329),
.B(n_276),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_376),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_241),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_330),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_215),
.Y(n_431)
);

NAND3x1_ASAP7_75t_L g432 ( 
.A(n_363),
.B(n_241),
.C(n_3),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_353),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_220),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_332),
.B(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_328),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_340),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_339),
.B(n_267),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_276),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_340),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_346),
.B(n_355),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_337),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_333),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_337),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_346),
.B(n_276),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_362),
.B(n_222),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_357),
.B(n_225),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_338),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_396),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_389),
.B(n_342),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_344),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_354),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_358),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_411),
.B(n_358),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_361),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_386),
.B(n_361),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_398),
.A2(n_378),
.B(n_374),
.C(n_373),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_443),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_408),
.B(n_378),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_368),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_368),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_424),
.A2(n_367),
.B1(n_372),
.B2(n_349),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_390),
.B(n_356),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_373),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_424),
.A2(n_349),
.B1(n_372),
.B2(n_367),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_394),
.B(n_383),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_384),
.A2(n_374),
.B1(n_338),
.B2(n_254),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_408),
.B(n_267),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_406),
.A2(n_267),
.B1(n_276),
.B2(n_228),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_455),
.B(n_229),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_399),
.B(n_233),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_397),
.B(n_4),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_418),
.B(n_4),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_406),
.A2(n_267),
.B1(n_234),
.B2(n_273),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_429),
.B(n_6),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_450),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_406),
.A2(n_402),
.B1(n_440),
.B2(n_453),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_394),
.B(n_235),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_429),
.B(n_6),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_449),
.B(n_335),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_387),
.B(n_7),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_447),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_388),
.B(n_243),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_441),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_387),
.B(n_244),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_388),
.B(n_245),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_404),
.A2(n_265),
.B(n_264),
.C(n_261),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_402),
.A2(n_248),
.B1(n_345),
.B2(n_9),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_402),
.A2(n_454),
.B1(n_445),
.B2(n_431),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_404),
.A2(n_7),
.B(n_8),
.C(n_10),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_8),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_385),
.B(n_11),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_385),
.B(n_11),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_388),
.B(n_12),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_12),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_392),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_400),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_416),
.B(n_13),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_388),
.B(n_13),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_402),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_402),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_528)
);

BUFx4f_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_L g530 ( 
.A1(n_423),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_422),
.A2(n_102),
.B(n_194),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_428),
.B(n_18),
.C(n_19),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

INVx8_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_393),
.B(n_21),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_454),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_22),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

AO22x1_ASAP7_75t_L g540 ( 
.A1(n_430),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_393),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_435),
.B(n_26),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_535),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_472),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_501),
.B(n_405),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_SL g546 ( 
.A(n_493),
.B(n_409),
.C(n_414),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_483),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_472),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_534),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_529),
.B(n_493),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_518),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_529),
.B(n_439),
.Y(n_553)
);

BUFx4f_ASAP7_75t_SL g554 ( 
.A(n_464),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_494),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_459),
.B(n_405),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_535),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_466),
.B(n_393),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_467),
.B(n_495),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_486),
.A2(n_445),
.B1(n_391),
.B2(n_427),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_427),
.B(n_401),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_524),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_499),
.B(n_436),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_498),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_468),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_531),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_498),
.B(n_433),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_539),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

NOR2x1p5_ASAP7_75t_SL g571 ( 
.A(n_462),
.B(n_490),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_475),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_476),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_463),
.B(n_420),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_508),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_465),
.B(n_445),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_520),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_489),
.B(n_445),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_495),
.B(n_417),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_521),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_489),
.B(n_491),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_509),
.A2(n_432),
.B1(n_401),
.B2(n_415),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_500),
.A2(n_421),
.B1(n_434),
.B2(n_412),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_473),
.B(n_410),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_536),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_470),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_479),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_458),
.B(n_410),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_497),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_512),
.B(n_412),
.Y(n_597)
);

AO22x1_ASAP7_75t_L g598 ( 
.A1(n_500),
.A2(n_452),
.B1(n_434),
.B2(n_426),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_SL g600 ( 
.A(n_537),
.B(n_420),
.C(n_415),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_504),
.B(n_433),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_491),
.B(n_413),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_562),
.A2(n_474),
.B(n_532),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_588),
.A2(n_487),
.B1(n_509),
.B2(n_510),
.Y(n_607)
);

AO31x2_ASAP7_75t_L g608 ( 
.A1(n_589),
.A2(n_471),
.A3(n_511),
.B(n_522),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_568),
.A2(n_474),
.B(n_514),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_593),
.A2(n_485),
.B(n_502),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_561),
.B(n_485),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_602),
.A2(n_515),
.B(n_517),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_486),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_552),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_545),
.B(n_492),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_548),
.A2(n_517),
.B(n_526),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_559),
.B(n_492),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_548),
.A2(n_526),
.B(n_542),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_565),
.B(n_471),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_548),
.A2(n_506),
.B(n_502),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_559),
.A2(n_488),
.B1(n_528),
.B2(n_527),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_555),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_578),
.A2(n_506),
.B(n_496),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_565),
.B(n_433),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_546),
.A2(n_511),
.B(n_530),
.C(n_484),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_496),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_590),
.A2(n_413),
.B(n_421),
.Y(n_630)
);

NOR2x1_ASAP7_75t_SL g631 ( 
.A(n_561),
.B(n_426),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_556),
.B(n_533),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_554),
.Y(n_634)
);

NOR2x1_ASAP7_75t_SL g635 ( 
.A(n_561),
.B(n_538),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_556),
.B(n_477),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_573),
.A2(n_505),
.B(n_507),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_584),
.A2(n_507),
.B(n_433),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_545),
.B(n_558),
.Y(n_639)
);

AOI221x1_ASAP7_75t_L g640 ( 
.A1(n_589),
.A2(n_540),
.B1(n_482),
.B2(n_477),
.C(n_452),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_27),
.C(n_28),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_565),
.B(n_482),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_551),
.A2(n_452),
.B(n_109),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_590),
.A2(n_452),
.B(n_108),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_452),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_544),
.A2(n_582),
.B(n_580),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_598),
.A2(n_107),
.B(n_192),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_564),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_27),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_547),
.B(n_28),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_SL g653 ( 
.A1(n_561),
.A2(n_110),
.B(n_191),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_574),
.B(n_30),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_549),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_574),
.A2(n_105),
.B(n_185),
.Y(n_656)
);

AOI21x1_ASAP7_75t_L g657 ( 
.A1(n_598),
.A2(n_103),
.B(n_184),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_595),
.B(n_30),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_580),
.A2(n_111),
.B(n_178),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_636),
.B(n_596),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_606),
.A2(n_582),
.B(n_580),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_606),
.A2(n_582),
.B(n_563),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_628),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_SL g664 ( 
.A(n_624),
.B(n_561),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_650),
.B(n_553),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_650),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_609),
.A2(n_569),
.B(n_563),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_652),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_634),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_566),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_641),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_629),
.B(n_563),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_609),
.A2(n_622),
.B(n_614),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_622),
.A2(n_569),
.B(n_577),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_607),
.A2(n_575),
.B1(n_603),
.B2(n_567),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_655),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_640),
.A2(n_569),
.A3(n_587),
.B(n_594),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_647),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_655),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_SL g681 ( 
.A(n_627),
.B(n_601),
.C(n_567),
.Y(n_681)
);

AO21x2_ASAP7_75t_L g682 ( 
.A1(n_621),
.A2(n_549),
.B(n_581),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_643),
.A2(n_604),
.B(n_605),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_643),
.A2(n_604),
.B(n_605),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_647),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_614),
.A2(n_577),
.B(n_583),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_617),
.A2(n_603),
.B1(n_592),
.B2(n_594),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_632),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_639),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_630),
.A2(n_577),
.B(n_583),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_612),
.B(n_543),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_630),
.A2(n_577),
.B(n_583),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_627),
.A2(n_587),
.B(n_594),
.C(n_581),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_621),
.A2(n_587),
.B(n_565),
.C(n_597),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_649),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_611),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_623),
.A2(n_560),
.B(n_595),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_620),
.A2(n_618),
.B(n_645),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_637),
.A2(n_597),
.B(n_585),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_649),
.B(n_543),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_651),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_648),
.Y(n_702)
);

AOI221xp5_ASAP7_75t_L g703 ( 
.A1(n_652),
.A2(n_592),
.B1(n_566),
.B2(n_599),
.C(n_585),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_633),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_619),
.B(n_591),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_619),
.A2(n_591),
.B1(n_570),
.B2(n_579),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_610),
.A2(n_591),
.B(n_570),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_638),
.A2(n_571),
.A3(n_576),
.B(n_570),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_642),
.B(n_591),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_620),
.A2(n_618),
.B(n_657),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_659),
.A2(n_557),
.B(n_543),
.Y(n_711)
);

OA21x2_ASAP7_75t_L g712 ( 
.A1(n_659),
.A2(n_625),
.B(n_615),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_677),
.Y(n_713)
);

AO21x2_ASAP7_75t_L g714 ( 
.A1(n_687),
.A2(n_626),
.B(n_654),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_666),
.B(n_658),
.Y(n_715)
);

NAND3x1_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_611),
.C(n_646),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_703),
.A2(n_579),
.B1(n_586),
.B2(n_611),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_673),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_697),
.A2(n_579),
.B1(n_586),
.B2(n_576),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_689),
.B(n_608),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_681),
.B(n_626),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_680),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_676),
.A2(n_579),
.B1(n_586),
.B2(n_613),
.Y(n_723)
);

AO31x2_ASAP7_75t_L g724 ( 
.A1(n_679),
.A2(n_635),
.A3(n_631),
.B(n_656),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_663),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_705),
.A2(n_701),
.B1(n_687),
.B2(n_699),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_SL g727 ( 
.A(n_681),
.B(n_709),
.C(n_684),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_705),
.A2(n_579),
.B1(n_586),
.B2(n_576),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_669),
.B(n_31),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_704),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_664),
.B(n_576),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_669),
.B(n_31),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_704),
.A2(n_706),
.B1(n_673),
.B2(n_683),
.Y(n_733)
);

OAI222xp33_ASAP7_75t_L g734 ( 
.A1(n_706),
.A2(n_608),
.B1(n_613),
.B2(n_644),
.C1(n_571),
.C2(n_557),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_704),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_673),
.A2(n_586),
.B1(n_579),
.B2(n_576),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_666),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_695),
.A2(n_586),
.B1(n_576),
.B2(n_557),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_710),
.A2(n_653),
.B(n_608),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_672),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_691),
.B(n_700),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_688),
.A2(n_557),
.B1(n_543),
.B2(n_608),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_707),
.B(n_195),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_671),
.B(n_32),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_679),
.A2(n_101),
.A3(n_175),
.B(n_174),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_R g746 ( 
.A(n_671),
.B(n_42),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_693),
.Y(n_747)
);

NAND2x1_ASAP7_75t_L g748 ( 
.A(n_668),
.B(n_43),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_682),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_671),
.B(n_34),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_665),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_691),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_668),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_696),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_670),
.B(n_38),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_693),
.B(n_176),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_685),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_700),
.B(n_45),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_678),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_L g760 ( 
.A1(n_694),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.C(n_54),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_682),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_691),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_712),
.A2(n_700),
.B1(n_702),
.B2(n_667),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_710),
.A2(n_56),
.B(n_58),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_678),
.B(n_59),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_702),
.Y(n_766)
);

BUFx12f_ASAP7_75t_L g767 ( 
.A(n_702),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_675),
.B(n_60),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_743),
.B(n_675),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_743),
.A2(n_694),
.B(n_661),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_743),
.A2(n_661),
.B(n_711),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_749),
.A2(n_702),
.B1(n_685),
.B2(n_712),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_764),
.A2(n_674),
.B(n_698),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_749),
.B(n_751),
.C(n_754),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_744),
.A2(n_712),
.B1(n_711),
.B2(n_678),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_762),
.B(n_708),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_725),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_L g778 ( 
.A1(n_717),
.A2(n_708),
.B1(n_662),
.B2(n_674),
.C(n_686),
.Y(n_778)
);

OAI211xp5_ASAP7_75t_L g779 ( 
.A1(n_729),
.A2(n_732),
.B(n_715),
.C(n_727),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_746),
.A2(n_708),
.B1(n_692),
.B2(n_690),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_752),
.B(n_708),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_713),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_730),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_752),
.B(n_686),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_740),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_754),
.B(n_62),
.C(n_63),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_SL g787 ( 
.A1(n_765),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_727),
.A2(n_756),
.B1(n_755),
.B2(n_723),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_752),
.B(n_70),
.Y(n_789)
);

OAI221xp5_ASAP7_75t_L g790 ( 
.A1(n_717),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.C(n_76),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_721),
.A2(n_79),
.B(n_80),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_737),
.B(n_84),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_726),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.C(n_91),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_735),
.B(n_94),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_714),
.A2(n_750),
.B1(n_744),
.B2(n_747),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_730),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_726),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_L g798 ( 
.A1(n_760),
.A2(n_99),
.B1(n_100),
.B2(n_112),
.C(n_113),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_720),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_768),
.A2(n_118),
.B(n_120),
.Y(n_800)
);

AOI322xp5_ASAP7_75t_L g801 ( 
.A1(n_733),
.A2(n_123),
.A3(n_124),
.B1(n_129),
.B2(n_131),
.C1(n_133),
.C2(n_136),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_733),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_735),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_722),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_759),
.Y(n_805)
);

AO21x2_ASAP7_75t_L g806 ( 
.A1(n_761),
.A2(n_151),
.B(n_152),
.Y(n_806)
);

INVxp33_ASAP7_75t_L g807 ( 
.A(n_730),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_730),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_768),
.A2(n_156),
.B1(n_159),
.B2(n_163),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_768),
.A2(n_764),
.B(n_734),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_165),
.Y(n_811)
);

AOI222xp33_ASAP7_75t_L g812 ( 
.A1(n_750),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.C1(n_170),
.C2(n_171),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_734),
.A2(n_172),
.B1(n_173),
.B2(n_742),
.C(n_714),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_719),
.A2(n_763),
.B1(n_728),
.B2(n_738),
.C(n_731),
.Y(n_814)
);

INVx8_ASAP7_75t_L g815 ( 
.A(n_752),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_777),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_784),
.B(n_763),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_805),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_785),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_776),
.B(n_757),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_782),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_775),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_815),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_769),
.B(n_757),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_769),
.B(n_739),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_781),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_769),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_795),
.B(n_739),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_773),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_815),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_788),
.B(n_766),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_810),
.B(n_741),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_771),
.B(n_745),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_815),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_783),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_778),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_770),
.B(n_745),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_772),
.B(n_745),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_813),
.B(n_745),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_806),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_811),
.B(n_718),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_780),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_796),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_791),
.B(n_719),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_791),
.B(n_724),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_812),
.B(n_724),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_774),
.A2(n_758),
.B(n_748),
.C(n_728),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_812),
.B(n_724),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_806),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_814),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_L g851 ( 
.A(n_850),
.B(n_801),
.C(n_786),
.Y(n_851)
);

AOI31xp33_ASAP7_75t_SL g852 ( 
.A1(n_822),
.A2(n_792),
.A3(n_793),
.B(n_800),
.Y(n_852)
);

OAI221xp5_ASAP7_75t_L g853 ( 
.A1(n_822),
.A2(n_779),
.B1(n_787),
.B2(n_802),
.C(n_790),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_817),
.B(n_807),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_846),
.A2(n_798),
.B1(n_797),
.B2(n_809),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_846),
.A2(n_799),
.B1(n_736),
.B2(n_794),
.Y(n_857)
);

NAND4xp25_ASAP7_75t_L g858 ( 
.A(n_850),
.B(n_737),
.C(n_794),
.D(n_753),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_817),
.B(n_753),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_818),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_820),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_818),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_820),
.B(n_724),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_836),
.B(n_804),
.C(n_803),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_825),
.B(n_811),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_817),
.B(n_767),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_846),
.A2(n_789),
.B(n_716),
.C(n_808),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_816),
.B(n_731),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_821),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_836),
.B(n_842),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_848),
.A2(n_831),
.B1(n_844),
.B2(n_839),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_819),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_872),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_859),
.B(n_836),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_859),
.B(n_842),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_870),
.B(n_832),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_862),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_862),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_870),
.B(n_832),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_865),
.B(n_825),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_861),
.B(n_819),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_854),
.B(n_825),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_865),
.B(n_848),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_871),
.B(n_835),
.Y(n_884)
);

AOI31xp33_ASAP7_75t_SL g885 ( 
.A1(n_856),
.A2(n_831),
.A3(n_827),
.B(n_828),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_854),
.B(n_866),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_855),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_855),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_SL g889 ( 
.A(n_884),
.B(n_848),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_881),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_883),
.A2(n_851),
.B1(n_864),
.B2(n_853),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_873),
.B(n_866),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_874),
.B(n_835),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_878),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_887),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_877),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_877),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_890),
.B(n_876),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_895),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_896),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_897),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_891),
.B(n_879),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_893),
.B(n_875),
.Y(n_904)
);

NOR2x1_ASAP7_75t_L g905 ( 
.A(n_903),
.B(n_858),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_904),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_902),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_SL g908 ( 
.A1(n_898),
.A2(n_892),
.B(n_883),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_901),
.B(n_889),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_907),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_905),
.B(n_902),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_906),
.B(n_899),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_909),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_910),
.Y(n_914)
);

AND3x2_ASAP7_75t_L g915 ( 
.A(n_913),
.B(n_900),
.C(n_880),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_911),
.Y(n_916)
);

OAI322xp33_ASAP7_75t_L g917 ( 
.A1(n_912),
.A2(n_908),
.A3(n_851),
.B1(n_883),
.B2(n_900),
.C1(n_889),
.C2(n_864),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_911),
.B(n_874),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_916),
.B(n_886),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_918),
.A2(n_867),
.B(n_839),
.C(n_837),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_914),
.B(n_917),
.Y(n_921)
);

AOI222xp33_ASAP7_75t_L g922 ( 
.A1(n_915),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.C1(n_885),
.C2(n_828),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_916),
.B(n_875),
.Y(n_923)
);

AOI221xp5_ASAP7_75t_L g924 ( 
.A1(n_917),
.A2(n_837),
.B1(n_833),
.B2(n_838),
.C(n_857),
.Y(n_924)
);

OAI211xp5_ASAP7_75t_SL g925 ( 
.A1(n_921),
.A2(n_847),
.B(n_852),
.C(n_868),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_924),
.B(n_858),
.C(n_895),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_919),
.B(n_844),
.C(n_833),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_922),
.B(n_844),
.C(n_833),
.Y(n_928)
);

OAI211xp5_ASAP7_75t_SL g929 ( 
.A1(n_923),
.A2(n_868),
.B(n_829),
.C(n_863),
.Y(n_929)
);

AOI211xp5_ASAP7_75t_SL g930 ( 
.A1(n_920),
.A2(n_880),
.B(n_865),
.C(n_845),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_926),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_925),
.B(n_880),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_927),
.B(n_882),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_928),
.Y(n_934)
);

XOR2xp5_ASAP7_75t_L g935 ( 
.A(n_930),
.B(n_865),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_931),
.A2(n_929),
.B(n_882),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_934),
.A2(n_845),
.B(n_838),
.C(n_849),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_830),
.Y(n_938)
);

NAND5xp2_ASAP7_75t_L g939 ( 
.A(n_933),
.B(n_845),
.C(n_824),
.D(n_823),
.E(n_830),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_935),
.B(n_888),
.Y(n_940)
);

AND2x2_ASAP7_75t_SL g941 ( 
.A(n_931),
.B(n_830),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_941),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_887),
.C(n_849),
.Y(n_943)
);

XOR2xp5_ASAP7_75t_L g944 ( 
.A(n_936),
.B(n_863),
.Y(n_944)
);

NAND4xp25_ASAP7_75t_L g945 ( 
.A(n_939),
.B(n_823),
.C(n_843),
.D(n_829),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_849),
.C(n_840),
.Y(n_946)
);

OAI221xp5_ASAP7_75t_L g947 ( 
.A1(n_937),
.A2(n_840),
.B1(n_834),
.B2(n_823),
.C(n_829),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_SL g948 ( 
.A1(n_938),
.A2(n_834),
.B1(n_843),
.B2(n_830),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_942),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_948),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

NAND5xp2_ASAP7_75t_L g952 ( 
.A(n_943),
.B(n_824),
.C(n_826),
.D(n_830),
.E(n_834),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_949),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_951),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_950),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_952),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_953),
.Y(n_957)
);

OAI22x1_ASAP7_75t_L g958 ( 
.A1(n_955),
.A2(n_945),
.B1(n_947),
.B2(n_946),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

OAI221xp5_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_956),
.B1(n_954),
.B2(n_843),
.C(n_840),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_959),
.A2(n_860),
.B(n_841),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_960),
.B(n_860),
.Y(n_962)
);

OA21x2_ASAP7_75t_L g963 ( 
.A1(n_961),
.A2(n_841),
.B(n_827),
.Y(n_963)
);

XNOR2x1_ASAP7_75t_L g964 ( 
.A(n_962),
.B(n_827),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_964),
.A2(n_830),
.B1(n_841),
.B2(n_869),
.Y(n_965)
);

OAI221xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_963),
.B1(n_830),
.B2(n_869),
.C(n_824),
.Y(n_966)
);

AOI211xp5_ASAP7_75t_L g967 ( 
.A1(n_966),
.A2(n_841),
.B(n_826),
.C(n_821),
.Y(n_967)
);


endmodule