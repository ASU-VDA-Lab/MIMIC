module real_aes_1628_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_0), .B(n_155), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_1), .A2(n_137), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_2), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_3), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_4), .A2(n_12), .B1(n_813), .B2(n_814), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_4), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_5), .B(n_145), .Y(n_201) );
INVx1_ASAP7_75t_L g142 ( .A(n_6), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_7), .B(n_145), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_8), .B(n_132), .Y(n_474) );
INVx1_ASAP7_75t_L g502 ( .A(n_9), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_10), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_11), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_12), .Y(n_813) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_13), .B(n_149), .Y(n_182) );
INVx2_ASAP7_75t_L g134 ( .A(n_14), .Y(n_134) );
AOI221x1_ASAP7_75t_L g224 ( .A1(n_15), .A2(n_27), .B1(n_137), .B2(n_155), .C(n_225), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_16), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_17), .B(n_155), .Y(n_178) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_18), .A2(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g483 ( .A(n_19), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_20), .B(n_168), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_21), .B(n_145), .Y(n_144) );
AO21x1_ASAP7_75t_L g196 ( .A1(n_22), .A2(n_155), .B(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g481 ( .A(n_24), .Y(n_481) );
INVx1_ASAP7_75t_SL g467 ( .A(n_25), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_26), .B(n_156), .Y(n_561) );
NAND2x1_ASAP7_75t_L g210 ( .A(n_28), .B(n_145), .Y(n_210) );
AOI33xp33_ASAP7_75t_L g529 ( .A1(n_29), .A2(n_53), .A3(n_457), .B1(n_464), .B2(n_530), .B3(n_531), .Y(n_529) );
NAND2x1_ASAP7_75t_L g164 ( .A(n_30), .B(n_149), .Y(n_164) );
INVx1_ASAP7_75t_L g511 ( .A(n_31), .Y(n_511) );
OR2x2_ASAP7_75t_L g133 ( .A(n_32), .B(n_86), .Y(n_133) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_32), .A2(n_86), .B(n_134), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_33), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_34), .B(n_149), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_35), .B(n_145), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_36), .B(n_149), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_37), .A2(n_137), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g138 ( .A(n_38), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g153 ( .A(n_38), .B(n_142), .Y(n_153) );
INVx1_ASAP7_75t_L g463 ( .A(n_38), .Y(n_463) );
OR2x6_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_40), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_41), .B(n_155), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_42), .B(n_455), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_43), .A2(n_132), .B1(n_172), .B2(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_44), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_45), .B(n_156), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_46), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_47), .B(n_149), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_48), .B(n_176), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_49), .B(n_156), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_50), .A2(n_137), .B(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_51), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_52), .B(n_149), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_54), .B(n_156), .Y(n_541) );
INVx1_ASAP7_75t_L g141 ( .A(n_55), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
AND2x2_ASAP7_75t_L g542 ( .A(n_56), .B(n_168), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_57), .A2(n_75), .B1(n_455), .B2(n_461), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_58), .B(n_455), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_59), .B(n_145), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_60), .B(n_172), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_61), .Y(n_804) );
AOI21xp5_ASAP7_75t_SL g491 ( .A1(n_62), .A2(n_461), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_63), .A2(n_137), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g477 ( .A(n_64), .Y(n_477) );
AO21x1_ASAP7_75t_L g198 ( .A1(n_65), .A2(n_137), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_66), .B(n_155), .Y(n_186) );
INVx1_ASAP7_75t_L g540 ( .A(n_67), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_68), .B(n_155), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_69), .A2(n_461), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g247 ( .A(n_70), .B(n_169), .Y(n_247) );
INVx1_ASAP7_75t_L g139 ( .A(n_71), .Y(n_139) );
INVx1_ASAP7_75t_L g147 ( .A(n_71), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_72), .A2(n_97), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_72), .Y(n_119) );
AND2x2_ASAP7_75t_L g170 ( .A(n_73), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_74), .B(n_455), .Y(n_532) );
AND2x2_ASAP7_75t_L g470 ( .A(n_76), .B(n_171), .Y(n_470) );
INVx1_ASAP7_75t_L g478 ( .A(n_77), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_78), .A2(n_461), .B(n_466), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_79), .A2(n_461), .B(n_524), .C(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_81), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g184 ( .A(n_82), .B(n_171), .Y(n_184) );
AND2x2_ASAP7_75t_SL g489 ( .A(n_83), .B(n_171), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_84), .A2(n_461), .B1(n_527), .B2(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g197 ( .A(n_85), .B(n_132), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_87), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g214 ( .A(n_88), .B(n_171), .Y(n_214) );
INVx1_ASAP7_75t_L g493 ( .A(n_89), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_90), .A2(n_118), .B1(n_786), .B2(n_790), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_91), .B(n_145), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_92), .A2(n_137), .B(n_143), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_93), .B(n_149), .Y(n_226) );
AND2x2_ASAP7_75t_L g533 ( .A(n_94), .B(n_171), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_95), .B(n_145), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_96), .A2(n_509), .B(n_510), .C(n_512), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_97), .Y(n_120) );
BUFx2_ASAP7_75t_L g796 ( .A(n_98), .Y(n_796) );
BUFx2_ASAP7_75t_SL g809 ( .A(n_98), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_99), .A2(n_137), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_100), .B(n_156), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_116), .B(n_818), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx4_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g821 ( .A(n_104), .Y(n_821) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_113), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g792 ( .A(n_107), .Y(n_792) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x6_ASAP7_75t_SL g444 ( .A(n_108), .B(n_109), .Y(n_444) );
OR2x6_ASAP7_75t_SL g783 ( .A(n_108), .B(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_108), .B(n_784), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_109), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_793), .B(n_805), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B(n_785), .Y(n_117) );
INVxp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_441), .B1(n_445), .B2(n_783), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g811 ( .A1(n_123), .A2(n_124), .B1(n_812), .B2(n_815), .Y(n_811) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_124), .A2(n_446), .B1(n_787), .B2(n_788), .Y(n_786) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_339), .Y(n_124) );
NAND3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_251), .C(n_306), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_191), .B1(n_215), .B2(n_219), .C(n_229), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_174), .Y(n_127) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_128), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g250 ( .A(n_128), .Y(n_250) );
AND2x2_ASAP7_75t_L g295 ( .A(n_128), .B(n_232), .Y(n_295) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_159), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g283 ( .A(n_130), .Y(n_283) );
INVx1_ASAP7_75t_L g293 ( .A(n_130), .Y(n_293) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B(n_157), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_131), .B(n_158), .Y(n_157) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_131), .A2(n_135), .B(n_157), .Y(n_257) );
INVx1_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_132), .A2(n_178), .B(n_179), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_132), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_132), .B(n_152), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_132), .A2(n_491), .B(n_495), .Y(n_490) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_133), .B(n_134), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_154), .Y(n_135) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
BUFx3_ASAP7_75t_L g459 ( .A(n_138), .Y(n_459) );
AND2x6_ASAP7_75t_L g149 ( .A(n_139), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g465 ( .A(n_139), .Y(n_465) );
AND2x4_ASAP7_75t_L g461 ( .A(n_140), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g145 ( .A(n_141), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g457 ( .A(n_141), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_142), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_152), .Y(n_143) );
INVxp67_ASAP7_75t_L g484 ( .A(n_145), .Y(n_484) );
AND2x4_ASAP7_75t_L g156 ( .A(n_146), .B(n_150), .Y(n_156) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVxp67_ASAP7_75t_L g482 ( .A(n_149), .Y(n_482) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_152), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_152), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_152), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_152), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_152), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_152), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_152), .A2(n_244), .B(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_152), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_152), .A2(n_468), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_152), .A2(n_468), .B(n_502), .C(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g527 ( .A(n_152), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_152), .A2(n_468), .B(n_540), .C(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_152), .A2(n_561), .B(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g155 ( .A(n_153), .B(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_153), .Y(n_512) );
INVx1_ASAP7_75t_L g479 ( .A(n_156), .Y(n_479) );
OR2x2_ASAP7_75t_L g272 ( .A(n_159), .B(n_175), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_159), .B(n_218), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_159), .B(n_183), .Y(n_316) );
INVx2_ASAP7_75t_L g325 ( .A(n_159), .Y(n_325) );
AND2x2_ASAP7_75t_L g346 ( .A(n_159), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g430 ( .A(n_159), .B(n_249), .Y(n_430) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g258 ( .A(n_160), .B(n_183), .Y(n_258) );
AND2x2_ASAP7_75t_L g391 ( .A(n_160), .B(n_218), .Y(n_391) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_160), .Y(n_417) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_167), .B(n_170), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_167), .A2(n_453), .B(n_470), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_168), .A2(n_186), .B(n_187), .Y(n_185) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_168), .A2(n_224), .B(n_228), .Y(n_223) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_168), .A2(n_224), .B(n_228), .Y(n_235) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_171), .A2(n_213), .B1(n_508), .B2(n_513), .Y(n_507) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_172), .B(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_173), .Y(n_176) );
AND2x4_ASAP7_75t_L g345 ( .A(n_174), .B(n_346), .Y(n_345) );
AOI321xp33_ASAP7_75t_L g359 ( .A1(n_174), .A2(n_288), .A3(n_289), .B1(n_321), .B2(n_360), .C(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_183), .Y(n_174) );
BUFx3_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVx2_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_175), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g282 ( .A(n_175), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g315 ( .A(n_175), .Y(n_315) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_176), .A2(n_500), .B(n_504), .Y(n_499) );
INVx2_ASAP7_75t_SL g524 ( .A(n_176), .Y(n_524) );
INVx5_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
NOR2x1_ASAP7_75t_SL g267 ( .A(n_183), .B(n_257), .Y(n_267) );
BUFx2_ASAP7_75t_L g362 ( .A(n_183), .Y(n_362) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_204), .Y(n_192) );
NOR2xp33_ASAP7_75t_SL g260 ( .A(n_193), .B(n_261), .Y(n_260) );
NOR4xp25_ASAP7_75t_L g363 ( .A(n_193), .B(n_357), .C(n_361), .D(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g401 ( .A(n_193), .Y(n_401) );
AND2x2_ASAP7_75t_L g435 ( .A(n_193), .B(n_375), .Y(n_435) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g236 ( .A(n_194), .Y(n_236) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g290 ( .A(n_195), .Y(n_290) );
OAI21x1_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_198), .B(n_202), .Y(n_195) );
INVx1_ASAP7_75t_L g203 ( .A(n_197), .Y(n_203) );
AOI33xp33_ASAP7_75t_L g431 ( .A1(n_204), .A2(n_233), .A3(n_264), .B1(n_280), .B2(n_386), .B3(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g221 ( .A(n_205), .B(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g231 ( .A(n_205), .B(n_232), .Y(n_231) );
BUFx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g238 ( .A(n_206), .Y(n_238) );
INVxp67_ASAP7_75t_L g319 ( .A(n_206), .Y(n_319) );
AND2x2_ASAP7_75t_L g375 ( .A(n_206), .B(n_240), .Y(n_375) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_213), .A2(n_241), .B(n_247), .Y(n_240) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_213), .A2(n_241), .B(n_247), .Y(n_276) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_213), .A2(n_536), .B(n_542), .Y(n_535) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_213), .A2(n_536), .B(n_542), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_215), .A2(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g384 ( .A(n_216), .B(n_258), .Y(n_384) );
AND3x2_ASAP7_75t_L g386 ( .A(n_216), .B(n_270), .C(n_325), .Y(n_386) );
INVx3_ASAP7_75t_SL g338 ( .A(n_217), .Y(n_338) );
INVx4_ASAP7_75t_L g232 ( .A(n_218), .Y(n_232) );
AND2x2_ASAP7_75t_L g270 ( .A(n_218), .B(n_257), .Y(n_270) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AND2x4_ASAP7_75t_L g289 ( .A(n_222), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g352 ( .A(n_222), .B(n_240), .Y(n_352) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g322 ( .A(n_223), .Y(n_322) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_223), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_R g229 ( .A1(n_230), .A2(n_233), .B(n_237), .C(n_248), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g281 ( .A(n_232), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_232), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_232), .B(n_249), .Y(n_410) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g392 ( .A(n_234), .B(n_382), .Y(n_392) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g239 ( .A(n_235), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g261 ( .A(n_235), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g277 ( .A(n_235), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g310 ( .A(n_235), .B(n_290), .Y(n_310) );
AND2x4_ASAP7_75t_L g275 ( .A(n_236), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g299 ( .A(n_236), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g337 ( .A(n_236), .B(n_262), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_262), .Y(n_265) );
AND2x2_ASAP7_75t_L g280 ( .A(n_238), .B(n_240), .Y(n_280) );
BUFx2_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_238), .B(n_261), .Y(n_350) );
INVx2_ASAP7_75t_L g262 ( .A(n_240), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_242), .B(n_246), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g298 ( .A1(n_248), .A2(n_299), .B1(n_301), .B2(n_305), .Y(n_298) );
INVx2_ASAP7_75t_SL g329 ( .A(n_248), .Y(n_329) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x2_ASAP7_75t_L g304 ( .A(n_249), .B(n_257), .Y(n_304) );
INVx1_ASAP7_75t_L g411 ( .A(n_250), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_284), .C(n_298), .Y(n_251) );
OAI221xp5_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_259), .B1(n_263), .B2(n_266), .C(n_268), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g312 ( .A(n_256), .Y(n_312) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_256), .Y(n_440) );
INVx1_ASAP7_75t_L g403 ( .A(n_258), .Y(n_403) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_258), .B(n_282), .Y(n_413) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_262), .B(n_290), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g296 ( .A(n_264), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g374 ( .A(n_264), .Y(n_374) );
AND2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_315), .Y(n_355) );
AND2x2_ASAP7_75t_L g432 ( .A(n_267), .B(n_430), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B1(n_280), .B2(n_281), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g291 ( .A(n_272), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx2_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
AND2x4_ASAP7_75t_L g321 ( .A(n_275), .B(n_322), .Y(n_321) );
OAI21xp33_ASAP7_75t_SL g351 ( .A1(n_275), .A2(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g378 ( .A(n_275), .B(n_336), .Y(n_378) );
INVx2_ASAP7_75t_L g300 ( .A(n_276), .Y(n_300) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
INVx1_ASAP7_75t_SL g357 ( .A(n_277), .Y(n_357) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g288 ( .A(n_279), .Y(n_288) );
AND2x4_ASAP7_75t_SL g382 ( .A(n_279), .B(n_300), .Y(n_382) );
AND2x2_ASAP7_75t_L g379 ( .A(n_282), .B(n_325), .Y(n_379) );
AND2x2_ASAP7_75t_L g405 ( .A(n_282), .B(n_391), .Y(n_405) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
INVx1_ASAP7_75t_L g347 ( .A(n_283), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_291), .B1(n_294), .B2(n_296), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_289), .B(n_300), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_289), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g428 ( .A(n_289), .Y(n_428) );
INVx2_ASAP7_75t_SL g353 ( .A(n_291), .Y(n_353) );
AND2x2_ASAP7_75t_L g365 ( .A(n_293), .B(n_325), .Y(n_365) );
INVx2_ASAP7_75t_L g371 ( .A(n_293), .Y(n_371) );
INVxp33_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_299), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g421 ( .A(n_299), .Y(n_421) );
INVx1_ASAP7_75t_L g349 ( .A(n_301), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_302), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_304), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_328), .C(n_331), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_313), .B2(n_317), .C(n_320), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g426 ( .A(n_311), .Y(n_426) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g395 ( .A(n_312), .B(n_361), .Y(n_395) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_315), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g397 ( .A(n_317), .Y(n_397) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g394 ( .A(n_318), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_319), .Y(n_400) );
OR2x2_ASAP7_75t_L g423 ( .A(n_319), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_SL g332 ( .A(n_322), .Y(n_332) );
AND2x2_ASAP7_75t_L g402 ( .A(n_322), .B(n_382), .Y(n_402) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_322), .B(n_335), .Y(n_434) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g439 ( .A(n_325), .Y(n_439) );
INVx1_ASAP7_75t_L g389 ( .A(n_327), .Y(n_389) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_334), .C(n_338), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_332), .B(n_382), .Y(n_406) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_335), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g343 ( .A(n_337), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g424 ( .A(n_337), .Y(n_424) );
NAND4xp75_ASAP7_75t_L g339 ( .A(n_340), .B(n_396), .C(n_412), .D(n_433), .Y(n_339) );
NOR3x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_358), .C(n_380), .Y(n_340) );
NAND4xp75_ASAP7_75t_L g341 ( .A(n_342), .B(n_348), .C(n_351), .D(n_354), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AND2x2_ASAP7_75t_L g393 ( .A(n_344), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g418 ( .A(n_345), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_SL g407 ( .A(n_350), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_366), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_362), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_372), .B(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g398 ( .A1(n_370), .A2(n_399), .A3(n_403), .B1(n_404), .B2(n_406), .C1(n_407), .C2(n_408), .Y(n_398) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_371), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_374), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_375), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_385), .C(n_387), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B1(n_393), .B2(n_395), .Y(n_387) );
NOR2xp33_ASAP7_75t_SL g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_402), .Y(n_399) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_405), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g415 ( .A(n_410), .B(n_416), .Y(n_415) );
O2A1O1Ixp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_419), .C(n_422), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_431), .Y(n_422) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx4_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx6p67_ASAP7_75t_R g787 ( .A(n_442), .Y(n_787) );
INVx3_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR3x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_648), .C(n_719), .Y(n_446) );
NAND3x1_ASAP7_75t_SL g447 ( .A(n_448), .B(n_575), .C(n_597), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_565), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_496), .B1(n_543), .B2(n_547), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_450), .A2(n_751), .B1(n_752), .B2(n_754), .Y(n_750) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_471), .Y(n_450) );
AND2x2_ASAP7_75t_L g566 ( .A(n_451), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_451), .B(n_613), .Y(n_632) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
AND2x2_ASAP7_75t_L g600 ( .A(n_452), .B(n_473), .Y(n_600) );
INVx1_ASAP7_75t_L g639 ( .A(n_452), .Y(n_639) );
OR2x2_ASAP7_75t_L g676 ( .A(n_452), .B(n_488), .Y(n_676) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_452), .Y(n_688) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_452), .Y(n_712) );
AND2x2_ASAP7_75t_L g769 ( .A(n_452), .B(n_596), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_460), .Y(n_453) );
INVx1_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g556 ( .A(n_456), .Y(n_556) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OR2x6_ASAP7_75t_L g468 ( .A(n_457), .B(n_465), .Y(n_468) );
INVxp33_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
INVx1_ASAP7_75t_L g557 ( .A(n_459), .Y(n_557) );
INVxp67_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
NOR2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_468), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_476) );
INVxp67_ASAP7_75t_L g509 ( .A(n_468), .Y(n_509) );
INVx2_ASAP7_75t_L g563 ( .A(n_468), .Y(n_563) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_486), .Y(n_471) );
INVx1_ASAP7_75t_L g644 ( .A(n_472), .Y(n_644) );
AND2x2_ASAP7_75t_L g670 ( .A(n_472), .B(n_488), .Y(n_670) );
NAND2x1_ASAP7_75t_L g686 ( .A(n_472), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g567 ( .A(n_473), .B(n_553), .Y(n_567) );
INVx3_ASAP7_75t_L g596 ( .A(n_473), .Y(n_596) );
NOR2x1_ASAP7_75t_SL g715 ( .A(n_473), .B(n_488), .Y(n_715) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_480), .B(n_485), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_479), .B(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_480) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_486), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g594 ( .A(n_487), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g564 ( .A(n_488), .Y(n_564) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_488), .Y(n_609) );
AND2x2_ASAP7_75t_L g681 ( .A(n_488), .B(n_553), .Y(n_681) );
AND2x4_ASAP7_75t_L g698 ( .A(n_488), .B(n_642), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_488), .B(n_640), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_488), .B(n_549), .Y(n_774) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_496), .A2(n_591), .B1(n_662), .B2(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_521), .Y(n_496) );
INVx2_ASAP7_75t_L g664 ( .A(n_497), .Y(n_664) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .Y(n_497) );
BUFx3_ASAP7_75t_L g654 ( .A(n_498), .Y(n_654) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_499), .B(n_523), .Y(n_546) );
INVx2_ASAP7_75t_L g570 ( .A(n_499), .Y(n_570) );
INVx1_ASAP7_75t_L g582 ( .A(n_499), .Y(n_582) );
AND2x4_ASAP7_75t_L g589 ( .A(n_499), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g606 ( .A(n_499), .B(n_506), .Y(n_606) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_499), .Y(n_620) );
INVxp67_ASAP7_75t_L g628 ( .A(n_499), .Y(n_628) );
AND2x2_ASAP7_75t_L g657 ( .A(n_505), .B(n_573), .Y(n_657) );
AND2x2_ASAP7_75t_L g673 ( .A(n_505), .B(n_574), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g760 ( .A(n_505), .B(n_573), .Y(n_760) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g569 ( .A(n_506), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
INVx1_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_506), .B(n_535), .Y(n_630) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_514), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g753 ( .A(n_521), .Y(n_753) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_534), .Y(n_521) );
AND2x2_ASAP7_75t_L g627 ( .A(n_522), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g656 ( .A(n_522), .Y(n_656) );
AND2x2_ASAP7_75t_L g758 ( .A(n_522), .B(n_573), .Y(n_758) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_523), .B(n_535), .Y(n_618) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_533), .Y(n_523) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_524), .A2(n_525), .B(n_533), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_526), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g544 ( .A(n_534), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g733 ( .A(n_534), .B(n_654), .Y(n_733) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_535), .Y(n_647) );
AND2x2_ASAP7_75t_L g674 ( .A(n_535), .B(n_620), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g588 ( .A(n_544), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g604 ( .A(n_544), .Y(n_604) );
AND2x2_ASAP7_75t_L g692 ( .A(n_544), .B(n_569), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_544), .B(n_712), .Y(n_717) );
AND2x2_ASAP7_75t_L g727 ( .A(n_544), .B(n_606), .Y(n_727) );
OR2x2_ASAP7_75t_L g764 ( .A(n_544), .B(n_664), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_545), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g724 ( .A(n_545), .B(n_580), .Y(n_724) );
AND2x2_ASAP7_75t_L g740 ( .A(n_545), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g734 ( .A(n_546), .B(n_630), .Y(n_734) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g616 ( .A(n_548), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_548), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g714 ( .A(n_548), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_548), .B(n_595), .Y(n_739) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_550), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_551), .A2(n_584), .B1(n_602), .B2(n_605), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_551), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g718 ( .A(n_551), .Y(n_718) );
AND2x4_ASAP7_75t_SL g551 ( .A(n_552), .B(n_564), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
INVx1_ASAP7_75t_L g642 ( .A(n_553), .Y(n_642) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .C(n_558), .Y(n_555) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
AND2x4_ASAP7_75t_L g641 ( .A(n_564), .B(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_564), .B(n_671), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
AND2x2_ASAP7_75t_L g666 ( .A(n_566), .B(n_609), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_566), .A2(n_747), .B(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g624 ( .A(n_567), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_568), .A2(n_678), .B1(n_682), .B2(n_685), .Y(n_677) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_569), .Y(n_635) );
AND2x2_ASAP7_75t_L g645 ( .A(n_569), .B(n_646), .Y(n_645) );
INVx3_ASAP7_75t_L g684 ( .A(n_569), .Y(n_684) );
NAND2x1_ASAP7_75t_SL g709 ( .A(n_569), .B(n_578), .Y(n_709) );
AND2x2_ASAP7_75t_L g605 ( .A(n_571), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_573), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g578 ( .A(n_574), .Y(n_578) );
INVx2_ASAP7_75t_L g590 ( .A(n_574), .Y(n_590) );
AOI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_583), .B(n_587), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_578), .B(n_772), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_668), .B1(n_672), .B2(n_675), .Y(n_667) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
BUFx2_ASAP7_75t_L g772 ( .A(n_580), .Y(n_772) );
INVx1_ASAP7_75t_SL g779 ( .A(n_580), .Y(n_779) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_581), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .B(n_594), .Y(n_587) );
AND2x2_ASAP7_75t_L g591 ( .A(n_589), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g633 ( .A(n_589), .B(n_629), .Y(n_633) );
AND2x2_ASAP7_75t_L g748 ( .A(n_589), .B(n_646), .Y(n_748) );
AND2x2_ASAP7_75t_L g751 ( .A(n_589), .B(n_657), .Y(n_751) );
AND2x4_ASAP7_75t_L g759 ( .A(n_589), .B(n_760), .Y(n_759) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_591), .A2(n_714), .B(n_716), .Y(n_713) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g741 ( .A(n_593), .Y(n_741) );
AND2x2_ASAP7_75t_L g757 ( .A(n_593), .B(n_758), .Y(n_757) );
INVx4_ASAP7_75t_L g671 ( .A(n_595), .Y(n_671) );
INVx1_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
AND2x2_ASAP7_75t_L g662 ( .A(n_596), .B(n_615), .Y(n_662) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_621), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_607), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_600), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_SL g761 ( .A(n_600), .B(n_613), .Y(n_761) );
AND2x2_ASAP7_75t_L g782 ( .A(n_600), .B(n_698), .Y(n_782) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g708 ( .A(n_605), .Y(n_708) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .B(n_617), .Y(n_607) );
OR2x6_ASAP7_75t_L g660 ( .A(n_609), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OR2x2_ASAP7_75t_L g683 ( .A(n_618), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g780 ( .A(n_618), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_619), .B(n_753), .Y(n_752) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_634), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_631), .B2(n_633), .Y(n_622) );
OR2x2_ASAP7_75t_L g694 ( .A(n_624), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g700 ( .A(n_629), .Y(n_700) );
INVx2_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_643), .B2(n_645), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
AND2x4_ASAP7_75t_SL g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g643 ( .A(n_641), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g704 ( .A(n_644), .B(n_698), .Y(n_704) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_689), .Y(n_648) );
NOR2xp67_ASAP7_75t_L g649 ( .A(n_650), .B(n_663), .Y(n_649) );
AOI21xp33_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_658), .Y(n_650) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp33_ASAP7_75t_SL g728 ( .A1(n_660), .A2(n_729), .B1(n_731), .B2(n_734), .Y(n_728) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_661), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g711 ( .A(n_662), .B(n_712), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_667), .C(n_677), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp33_ASAP7_75t_SL g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVxp33_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g680 ( .A(n_671), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_672), .A2(n_692), .B1(n_693), .B2(n_696), .C(n_699), .Y(n_691) );
AND2x4_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g732 ( .A(n_673), .Y(n_732) );
INVx2_ASAP7_75t_SL g730 ( .A(n_676), .Y(n_730) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2x1_ASAP7_75t_L g729 ( .A(n_680), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g726 ( .A(n_686), .Y(n_726) );
INVx1_ASAP7_75t_L g755 ( .A(n_687), .Y(n_755) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_705), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_703), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g744 ( .A(n_695), .Y(n_744) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g765 ( .A(n_698), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g770 ( .A(n_698), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVxp33_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx2_ASAP7_75t_L g723 ( .A(n_702), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_710), .B(n_713), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g766 ( .A(n_712), .Y(n_766) );
AND2x2_ASAP7_75t_L g754 ( .A(n_715), .B(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_R g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_735), .C(n_762), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_722), .B(n_725), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_749), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_737), .B(n_746), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_745), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_750), .B(n_756), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g775 ( .A(n_759), .Y(n_775) );
AOI211xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B(n_767), .C(n_776), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_771), .B1(n_773), .B2(n_775), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVxp67_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_783), .Y(n_789) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_798), .A2(n_811), .B(n_816), .Y(n_810) );
NOR2xp33_ASAP7_75t_SL g798 ( .A(n_799), .B(n_804), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
BUFx3_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
BUFx2_ASAP7_75t_L g817 ( .A(n_803), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx8_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_812), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
endmodule