module fake_ibex_91_n_3464 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3464);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3464;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_2183;
wire n_1859;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_667;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_3323;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_2333;
wire n_715;
wire n_1910;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2980;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2999;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_2732;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3333;
wire n_3096;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2348;
wire n_2093;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3305;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3051;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_632;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_1532;
wire n_791;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3225;
wire n_2652;
wire n_2227;
wire n_3380;
wire n_1074;
wire n_3067;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_3124;
wire n_999;
wire n_2634;
wire n_3286;
wire n_2982;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_2186;
wire n_1843;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_683;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

INVx2_ASAP7_75t_L g630 ( 
.A(n_158),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_270),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_223),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_423),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_384),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_131),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_422),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_280),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_99),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_416),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_193),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_58),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_382),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_451),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_100),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_454),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_504),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_227),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_383),
.Y(n_650)
);

INVxp33_ASAP7_75t_SL g651 ( 
.A(n_605),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_1),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_79),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_477),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_402),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_113),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_512),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_310),
.Y(n_658)
);

CKINVDCx14_ASAP7_75t_R g659 ( 
.A(n_430),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_79),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_266),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_54),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_149),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_250),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_217),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_161),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_568),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_8),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_419),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_536),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_390),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_7),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_519),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_92),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_613),
.B(n_136),
.Y(n_675)
);

BUFx8_ASAP7_75t_SL g676 ( 
.A(n_125),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_54),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_104),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_571),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_627),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_256),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_18),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_282),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_552),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_495),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_134),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_516),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_538),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_500),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_131),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_564),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_182),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_447),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_413),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_441),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_41),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_523),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_324),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_587),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_445),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_509),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_154),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_592),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_163),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_466),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_324),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_318),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_522),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_229),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_155),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_85),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_488),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_453),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_24),
.B(n_335),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_455),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_342),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_629),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_72),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_276),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_315),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_29),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_585),
.Y(n_723)
);

BUFx5_ASAP7_75t_L g724 ( 
.A(n_498),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_462),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_276),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_107),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_582),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_548),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_549),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_321),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_414),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_434),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_426),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_576),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_136),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_42),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_604),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_101),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_338),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_496),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_184),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_530),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_228),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_513),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_207),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_597),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_506),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_23),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_268),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_350),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_529),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_228),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_562),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_457),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_511),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_118),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_94),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_339),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_317),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_279),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_85),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_223),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_14),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_40),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_116),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_599),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_201),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_45),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_461),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_21),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_542),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_217),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_591),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_401),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_351),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_399),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_269),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_247),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_534),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_1),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_567),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_63),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_566),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_395),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_66),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_203),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_147),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_113),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_590),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_596),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_238),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_520),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_235),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_403),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_301),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_73),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_569),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_71),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_9),
.B(n_226),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_484),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_602),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_199),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_535),
.B(n_481),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_326),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_550),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_537),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_318),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_518),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_372),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_545),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_429),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_281),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_21),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_64),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_159),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_114),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_63),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_505),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_628),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_45),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_565),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_547),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_62),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_399),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_624),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_486),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_316),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_43),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_32),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_558),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_256),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_617),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_157),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_135),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_468),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_174),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_336),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_365),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_198),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_185),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_293),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_449),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_14),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_382),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_246),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_351),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_431),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_330),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_176),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_224),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_178),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_581),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_446),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_463),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_316),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_232),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_282),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_331),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_271),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_373),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_321),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_393),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_91),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_92),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_84),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_203),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_398),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_433),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_479),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_573),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_208),
.Y(n_873)
);

CKINVDCx14_ASAP7_75t_R g874 ( 
.A(n_410),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_485),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_253),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_623),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_6),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_156),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_372),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_60),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_55),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_67),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_452),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_144),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_284),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_300),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_155),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_167),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_227),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_616),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_428),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_356),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_124),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_546),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_376),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_29),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_124),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_586),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_492),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_194),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_470),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_557),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_606),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_472),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_360),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_83),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_326),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_483),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_361),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_600),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_341),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_116),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_584),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_214),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_74),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_390),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_611),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_257),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_70),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_292),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_615),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_130),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_594),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_577),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_22),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_489),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_369),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_251),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_258),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_539),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_377),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_344),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_595),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_556),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_115),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_307),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_598),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_296),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_272),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_490),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_464),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_381),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_342),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_185),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_23),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_171),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_521),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_205),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_9),
.Y(n_950)
);

XOR2xp5_ASAP7_75t_L g951 ( 
.A(n_373),
.B(n_225),
.Y(n_951)
);

BUFx5_ASAP7_75t_L g952 ( 
.A(n_44),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_319),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_308),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_16),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_544),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_366),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_74),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_575),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_363),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_450),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_154),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_141),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_13),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_559),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_563),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_129),
.Y(n_967)
);

BUFx10_ASAP7_75t_L g968 ( 
.A(n_138),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_187),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_579),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_473),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_190),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_134),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_358),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_366),
.Y(n_975)
);

BUFx8_ASAP7_75t_SL g976 ( 
.A(n_601),
.Y(n_976)
);

CKINVDCx16_ASAP7_75t_R g977 ( 
.A(n_497),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_220),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_180),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_231),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_329),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_322),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_254),
.Y(n_983)
);

BUFx10_ASAP7_75t_L g984 ( 
.A(n_56),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_572),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_603),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_105),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_265),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_42),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_614),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_202),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_193),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_105),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_255),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_389),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_713),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_976),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_874),
.B(n_0),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_722),
.Y(n_999)
);

OA21x2_ASAP7_75t_L g1000 ( 
.A1(n_733),
.A2(n_421),
.B(n_420),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_903),
.Y(n_1001)
);

CKINVDCx16_ASAP7_75t_R g1002 ( 
.A(n_656),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_722),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_726),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_708),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_708),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_903),
.A2(n_425),
.B(n_424),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_733),
.A2(n_781),
.B(n_765),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_726),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_874),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_676),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_713),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_666),
.B(n_2),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_713),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_883),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_713),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_R g1017 ( 
.A(n_689),
.B(n_990),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_666),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_726),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_818),
.B(n_3),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_818),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_972),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_868),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_868),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_972),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_708),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_708),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_765),
.A2(n_432),
.B(n_427),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_630),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_652),
.B(n_5),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_630),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_718),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_868),
.Y(n_1034)
);

INVx6_ASAP7_75t_L g1035 ( 
.A(n_697),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_708),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_708),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_718),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_708),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_705),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_676),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_677),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_718),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_639),
.Y(n_1044)
);

AND2x6_ASAP7_75t_L g1045 ( 
.A(n_645),
.B(n_435),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_697),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_731),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_718),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

XNOR2xp5_ASAP7_75t_L g1050 ( 
.A(n_951),
.B(n_8),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_697),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_658),
.B(n_10),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_952),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_952),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_658),
.B(n_10),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_770),
.B(n_11),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_704),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_712),
.B(n_11),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_819),
.B(n_12),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_704),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_724),
.B(n_781),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_704),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_976),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_755),
.Y(n_1064)
);

OA21x2_ASAP7_75t_L g1065 ( 
.A1(n_875),
.A2(n_437),
.B(n_436),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_963),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_963),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_712),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_812),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_720),
.B(n_12),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_720),
.B(n_13),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_755),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_830),
.B(n_936),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_755),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_835),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_963),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_952),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_884),
.B(n_15),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_919),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_952),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_955),
.Y(n_1081)
);

BUFx8_ASAP7_75t_SL g1082 ( 
.A(n_637),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_952),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_921),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_820),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_955),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_968),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_882),
.B(n_16),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_930),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_875),
.A2(n_439),
.B(n_438),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_631),
.B(n_17),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_982),
.B(n_17),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_638),
.B(n_18),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_977),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_968),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_959),
.A2(n_442),
.B(n_440),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_997),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_997),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_1002),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1063),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1052),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1063),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1082),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1082),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_1035),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_1017),
.B(n_659),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_1011),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1061),
.A2(n_1008),
.B(n_1027),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1011),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_999),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1069),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_1041),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1052),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_1041),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1035),
.B(n_959),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1003),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1061),
.A2(n_648),
.B(n_633),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1055),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1069),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1094),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1094),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1055),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1004),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_1017),
.B(n_659),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1047),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1084),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1015),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1025),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1066),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1058),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1076),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1087),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1046),
.B(n_967),
.Y(n_1133)
);

BUFx10_ASAP7_75t_L g1134 ( 
.A(n_1035),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_1015),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1005),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1079),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1079),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1058),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1089),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1089),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1042),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1088),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_1009),
.B(n_670),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1027),
.A2(n_673),
.B(n_657),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1070),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1070),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1042),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_1009),
.B(n_670),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_1024),
.B(n_714),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1046),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1006),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_1024),
.B(n_714),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1034),
.B(n_1095),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1046),
.B(n_687),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1046),
.B(n_987),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_R g1157 ( 
.A(n_1034),
.B(n_771),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_998),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1071),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1051),
.B(n_1057),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1092),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1051),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1051),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1092),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1051),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1013),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1057),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1045),
.Y(n_1168)
);

NOR2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1095),
.B(n_1073),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1057),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1057),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_1060),
.B(n_771),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1060),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1060),
.B(n_823),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1036),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1060),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1050),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_R g1178 ( 
.A(n_1020),
.B(n_1067),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1037),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1062),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1073),
.B(n_968),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1062),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_R g1183 ( 
.A(n_1013),
.B(n_651),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_1021),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1062),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1039),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1021),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1093),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1062),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1056),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1053),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1093),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1085),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1019),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1085),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1085),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_1040),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_R g1198 ( 
.A(n_1085),
.B(n_1018),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1040),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1022),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1001),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_R g1202 ( 
.A(n_1000),
.B(n_991),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1023),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1010),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1001),
.B(n_642),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1078),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1001),
.B(n_693),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1026),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1031),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1001),
.B(n_650),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1031),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1045),
.B(n_823),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1030),
.B(n_984),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_L g1214 ( 
.A(n_1032),
.B(n_695),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1059),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1059),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1091),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1054),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1044),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1045),
.Y(n_1220)
);

INVxp33_ASAP7_75t_L g1221 ( 
.A(n_1091),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_R g1222 ( 
.A(n_1045),
.B(n_895),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1068),
.B(n_699),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1075),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1081),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1086),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1077),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1028),
.B(n_984),
.Y(n_1228)
);

CKINVDCx16_ASAP7_75t_R g1229 ( 
.A(n_1045),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_996),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1080),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1029),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1028),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1049),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1083),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_996),
.B(n_895),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_996),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1000),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1065),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1012),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1012),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_R g1242 ( 
.A(n_1012),
.B(n_900),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1014),
.B(n_980),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1065),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1090),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1096),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1014),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1014),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1090),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1016),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1007),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1016),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1016),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1033),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1033),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1033),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1038),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1038),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_R g1259 ( 
.A(n_1038),
.B(n_900),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1074),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1043),
.B(n_701),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1043),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1043),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1048),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1048),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1048),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1064),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1064),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1064),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1072),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1072),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_R g1272 ( 
.A(n_1072),
.B(n_983),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1074),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1074),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1052),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1015),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_997),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1002),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_997),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_997),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1202),
.B(n_735),
.C(n_723),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1246),
.A2(n_756),
.B(n_743),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1221),
.B(n_820),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1228),
.B(n_952),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1110),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1168),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1211),
.B(n_636),
.Y(n_1287)
);

INVxp33_ASAP7_75t_L g1288 ( 
.A(n_1276),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1215),
.B(n_643),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1216),
.B(n_646),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1201),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1181),
.B(n_647),
.Y(n_1292)
);

NAND2x1_ASAP7_75t_L g1293 ( 
.A(n_1201),
.B(n_805),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1229),
.B(n_820),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1219),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

INVx8_ASAP7_75t_L g1297 ( 
.A(n_1137),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1226),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1168),
.B(n_870),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1194),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1197),
.B(n_814),
.C(n_761),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1220),
.B(n_870),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1213),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1169),
.B(n_654),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_SL g1305 ( 
.A(n_1105),
.Y(n_1305)
);

AO221x1_ASAP7_75t_L g1306 ( 
.A1(n_1144),
.A2(n_753),
.B1(n_764),
.B2(n_707),
.C(n_637),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1126),
.Y(n_1307)
);

CKINVDCx8_ASAP7_75t_R g1308 ( 
.A(n_1103),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1206),
.B(n_870),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1108),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1200),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1203),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1127),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1208),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1224),
.B(n_667),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1225),
.B(n_669),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1166),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1187),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1138),
.B(n_984),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1115),
.B(n_679),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1101),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1233),
.B(n_680),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1205),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1220),
.B(n_1184),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1184),
.B(n_684),
.Y(n_1325)
);

INVx8_ASAP7_75t_L g1326 ( 
.A(n_1140),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1141),
.B(n_688),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1113),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1254),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1188),
.B(n_691),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1192),
.B(n_685),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1105),
.B(n_927),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1142),
.B(n_632),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1134),
.B(n_700),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1148),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1210),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1145),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1118),
.B(n_703),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1134),
.B(n_706),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1122),
.B(n_709),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1130),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1183),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1139),
.B(n_716),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1146),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1133),
.B(n_725),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1147),
.B(n_728),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1199),
.B(n_786),
.C(n_740),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1159),
.B(n_729),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1161),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_L g1351 ( 
.A(n_1202),
.B(n_803),
.C(n_794),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1260),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1212),
.B(n_730),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1251),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1125),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1164),
.B(n_734),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1123),
.B(n_1128),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1275),
.B(n_738),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_L g1359 ( 
.A(n_1204),
.B(n_1119),
.C(n_1111),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1156),
.B(n_741),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1151),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1176),
.B(n_1209),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1243),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1231),
.B(n_745),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1212),
.B(n_1198),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1198),
.B(n_747),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1214),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1207),
.A2(n_661),
.B(n_665),
.C(n_664),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1246),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1120),
.B(n_920),
.C(n_806),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1223),
.Y(n_1371)
);

OR2x2_ASAP7_75t_SL g1372 ( 
.A(n_1135),
.B(n_707),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1217),
.B(n_748),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1154),
.B(n_752),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1154),
.B(n_754),
.Y(n_1376)
);

NAND2xp33_ASAP7_75t_L g1377 ( 
.A(n_1222),
.B(n_724),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1261),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1239),
.B(n_821),
.C(n_807),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1230),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1106),
.B(n_634),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1162),
.B(n_768),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1249),
.B(n_849),
.C(n_827),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1207),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1236),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1163),
.B(n_773),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1232),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1165),
.B(n_775),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1167),
.B(n_783),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1230),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_L g1391 ( 
.A(n_1238),
.B(n_1244),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1124),
.B(n_785),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_1245),
.B(n_1172),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1241),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1160),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1155),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1155),
.Y(n_1397)
);

NOR3xp33_ASAP7_75t_L g1398 ( 
.A(n_1121),
.B(n_944),
.C(n_644),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_SL g1399 ( 
.A(n_1232),
.B(n_828),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1173),
.B(n_792),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1180),
.B(n_799),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1182),
.B(n_802),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1242),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1185),
.B(n_808),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1189),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1242),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1234),
.B(n_854),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1241),
.Y(n_1409)
);

NOR2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1129),
.B(n_640),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_L g1411 ( 
.A(n_1172),
.B(n_724),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1235),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1193),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1237),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1149),
.B(n_649),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1227),
.B(n_855),
.Y(n_1416)
);

AO221x1_ASAP7_75t_L g1417 ( 
.A1(n_1144),
.A2(n_1153),
.B1(n_1157),
.B2(n_1150),
.C(n_1174),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1195),
.B(n_810),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1196),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1240),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1136),
.B(n_813),
.Y(n_1421)
);

NAND2xp33_ASAP7_75t_L g1422 ( 
.A(n_1174),
.B(n_724),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1117),
.A2(n_871),
.B(n_856),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1152),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1175),
.B(n_824),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_L g1426 ( 
.A(n_1259),
.B(n_724),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1179),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1153),
.B(n_653),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1186),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1247),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1191),
.B(n_837),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1218),
.B(n_1178),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1190),
.B(n_844),
.Y(n_1433)
);

NOR2xp67_ASAP7_75t_L g1434 ( 
.A(n_1248),
.B(n_448),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1253),
.A2(n_877),
.B(n_872),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1158),
.B(n_892),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1273),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1259),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1143),
.B(n_899),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1157),
.B(n_902),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1250),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1252),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1255),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1256),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1257),
.B(n_909),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1131),
.B(n_914),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_L g1447 ( 
.A(n_1132),
.B(n_724),
.Y(n_1447)
);

BUFx5_ASAP7_75t_L g1448 ( 
.A(n_1262),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1263),
.Y(n_1449)
);

BUFx8_ASAP7_75t_L g1450 ( 
.A(n_1104),
.Y(n_1450)
);

NOR3xp33_ASAP7_75t_L g1451 ( 
.A(n_1097),
.B(n_660),
.C(n_655),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1280),
.B(n_832),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1099),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1265),
.B(n_918),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1266),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1267),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1098),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1268),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1278),
.B(n_924),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1100),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_L g1461 ( 
.A(n_1102),
.B(n_663),
.C(n_662),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1277),
.B(n_934),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1269),
.B(n_938),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1183),
.B(n_941),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1279),
.B(n_975),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1258),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1272),
.B(n_942),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1258),
.B(n_956),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1177),
.B(n_961),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1272),
.B(n_715),
.Y(n_1470)
);

BUFx5_ASAP7_75t_L g1471 ( 
.A(n_1264),
.Y(n_1471)
);

AND2x6_ASAP7_75t_SL g1472 ( 
.A(n_1107),
.B(n_753),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1270),
.B(n_965),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1271),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1274),
.B(n_966),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1109),
.B(n_971),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1112),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1114),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1126),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1221),
.B(n_668),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1221),
.B(n_671),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1221),
.B(n_891),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1221),
.B(n_672),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1229),
.B(n_970),
.Y(n_1484)
);

INVxp33_ASAP7_75t_L g1485 ( 
.A(n_1276),
.Y(n_1485)
);

BUFx5_ASAP7_75t_L g1486 ( 
.A(n_1168),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1221),
.B(n_674),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1105),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1204),
.A2(n_686),
.B1(n_690),
.B2(n_678),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1229),
.B(n_985),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1229),
.B(n_986),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1201),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1110),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_SL g1494 ( 
.A(n_1168),
.B(n_645),
.Y(n_1494)
);

XNOR2xp5_ASAP7_75t_L g1495 ( 
.A(n_1099),
.B(n_764),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1110),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1221),
.B(n_904),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1221),
.B(n_905),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1229),
.B(n_911),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1229),
.B(n_922),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1201),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1201),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1254),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1201),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1221),
.B(n_925),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1201),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1221),
.B(n_681),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1201),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1166),
.A2(n_694),
.B1(n_698),
.B2(n_692),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1221),
.B(n_682),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1166),
.A2(n_710),
.B1(n_727),
.B2(n_702),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1229),
.B(n_931),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1201),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1110),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1201),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1201),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1229),
.B(n_935),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1110),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1221),
.B(n_696),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1110),
.Y(n_1520)
);

NAND2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1228),
.B(n_736),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1110),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1110),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1276),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1201),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1201),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1221),
.B(n_711),
.Y(n_1527)
);

INVxp33_ASAP7_75t_L g1528 ( 
.A(n_1276),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1221),
.B(n_717),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1201),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1110),
.Y(n_1531)
);

AND2x6_ASAP7_75t_L g1532 ( 
.A(n_1168),
.B(n_948),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1105),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1221),
.B(n_719),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1221),
.B(n_721),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1201),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1105),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1110),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1281),
.A2(n_797),
.B1(n_876),
.B2(n_774),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1313),
.Y(n_1540)
);

NOR2xp67_ASAP7_75t_L g1541 ( 
.A(n_1336),
.B(n_19),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1288),
.B(n_635),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1298),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_732),
.Y(n_1544)
);

NOR2x2_ASAP7_75t_L g1545 ( 
.A(n_1355),
.B(n_1495),
.Y(n_1545)
);

INVx5_ASAP7_75t_L g1546 ( 
.A(n_1409),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1498),
.B(n_739),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1369),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1297),
.B(n_801),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_L g1550 ( 
.A(n_1410),
.B(n_1357),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1313),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1307),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1354),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1297),
.B(n_737),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1524),
.A2(n_1399),
.B1(n_1343),
.B2(n_1529),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1286),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1300),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1485),
.B(n_774),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1295),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1528),
.B(n_744),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1521),
.B(n_1317),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1297),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1334),
.B(n_797),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1307),
.Y(n_1564)
);

XOR2x2_ASAP7_75t_L g1565 ( 
.A(n_1479),
.B(n_969),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1326),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1409),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1329),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1479),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1311),
.Y(n_1570)
);

BUFx4f_ASAP7_75t_L g1571 ( 
.A(n_1326),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1409),
.B(n_750),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1318),
.B(n_751),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1312),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1281),
.A2(n_885),
.B1(n_887),
.B2(n_876),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1286),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_R g1577 ( 
.A(n_1326),
.B(n_885),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1286),
.Y(n_1578)
);

AOI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1494),
.A2(n_675),
.B(n_742),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1314),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1477),
.B(n_746),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1534),
.B(n_757),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1535),
.B(n_759),
.C(n_758),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1482),
.B(n_760),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1503),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1497),
.B(n_762),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1321),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1477),
.B(n_749),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_SL g1589 ( 
.A(n_1370),
.B(n_898),
.C(n_887),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1505),
.B(n_763),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1332),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1285),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1296),
.Y(n_1593)
);

AND2x6_ASAP7_75t_L g1594 ( 
.A(n_1387),
.B(n_755),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1351),
.A2(n_933),
.B1(n_969),
.B2(n_898),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1303),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1406),
.B(n_1413),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1301),
.A2(n_772),
.B1(n_777),
.B2(n_766),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1450),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1387),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_R g1601 ( 
.A(n_1308),
.B(n_933),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1424),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1407),
.B(n_778),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1427),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1328),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1319),
.B(n_683),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1428),
.B(n_779),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1342),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1345),
.B(n_782),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1350),
.B(n_784),
.Y(n_1610)
);

NAND2x1_ASAP7_75t_L g1611 ( 
.A(n_1532),
.B(n_791),
.Y(n_1611)
);

NAND2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1488),
.B(n_767),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1362),
.B(n_842),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1429),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1532),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1419),
.B(n_780),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1538),
.Y(n_1617)
);

INVx3_ASAP7_75t_SL g1618 ( 
.A(n_1477),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_L g1619 ( 
.A(n_1532),
.B(n_1486),
.Y(n_1619)
);

NAND2x1p5_ASAP7_75t_L g1620 ( 
.A(n_1533),
.B(n_787),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1332),
.B(n_869),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1480),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1481),
.B(n_788),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1337),
.Y(n_1624)
);

AND2x6_ASAP7_75t_L g1625 ( 
.A(n_1363),
.B(n_791),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1483),
.B(n_789),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1487),
.B(n_790),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1287),
.B(n_793),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1351),
.A2(n_798),
.B1(n_815),
.B2(n_804),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1507),
.B(n_816),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1478),
.B(n_796),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1537),
.B(n_800),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1510),
.B(n_1519),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1527),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1303),
.Y(n_1635)
);

BUFx4f_ASAP7_75t_L g1636 ( 
.A(n_1478),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1493),
.Y(n_1637)
);

BUFx8_ASAP7_75t_L g1638 ( 
.A(n_1305),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1283),
.B(n_822),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1496),
.B(n_1514),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1518),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1289),
.B(n_826),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1520),
.B(n_831),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1522),
.B(n_836),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1523),
.B(n_838),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1531),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1290),
.B(n_839),
.Y(n_1647)
);

INVx3_ASAP7_75t_SL g1648 ( 
.A(n_1478),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1442),
.B(n_840),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1532),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1292),
.B(n_841),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1323),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1361),
.B(n_809),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1450),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1442),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1442),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1361),
.B(n_811),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1331),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1412),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1372),
.A2(n_848),
.B1(n_850),
.B2(n_843),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1380),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1291),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1309),
.A2(n_858),
.B1(n_861),
.B2(n_857),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1464),
.B(n_863),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1325),
.B(n_825),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1305),
.Y(n_1666)
);

BUFx4f_ASAP7_75t_L g1667 ( 
.A(n_1457),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1472),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1452),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1452),
.Y(n_1670)
);

BUFx4f_ASAP7_75t_SL g1671 ( 
.A(n_1453),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1374),
.B(n_862),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1509),
.B(n_864),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1294),
.B(n_829),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1415),
.B(n_867),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1284),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1284),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1433),
.B(n_878),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1352),
.Y(n_1679)
);

AND3x1_ASAP7_75t_L g1680 ( 
.A(n_1359),
.B(n_845),
.C(n_833),
.Y(n_1680)
);

AND2x4_ASAP7_75t_SL g1681 ( 
.A(n_1460),
.B(n_847),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1511),
.B(n_880),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1356),
.B(n_881),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1432),
.B(n_890),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1391),
.A2(n_852),
.B1(n_853),
.B2(n_851),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1465),
.B(n_896),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1408),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1489),
.A2(n_981),
.B1(n_989),
.B2(n_978),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1408),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1492),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1437),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1322),
.B(n_901),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1367),
.B(n_860),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1315),
.B(n_908),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1436),
.B(n_910),
.Y(n_1695)
);

NOR2xp67_ASAP7_75t_L g1696 ( 
.A(n_1469),
.B(n_19),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1371),
.B(n_865),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1416),
.Y(n_1698)
);

NOR2x2_ASAP7_75t_L g1699 ( 
.A(n_1472),
.B(n_912),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1416),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1390),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1293),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1394),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1501),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1396),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1327),
.B(n_866),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1381),
.B(n_913),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1385),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1316),
.B(n_1346),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1439),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1502),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1398),
.B(n_928),
.C(n_926),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1397),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1459),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1384),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1339),
.B(n_929),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1341),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1504),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1344),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1404),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1347),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1395),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1349),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1438),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1506),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1414),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1420),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1508),
.Y(n_1728)
);

INVx5_ASAP7_75t_L g1729 ( 
.A(n_1470),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1358),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1470),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1486),
.B(n_939),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1373),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1476),
.A2(n_943),
.B1(n_945),
.B2(n_940),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1446),
.B(n_946),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1470),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1513),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1378),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1368),
.B(n_1282),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1379),
.A2(n_879),
.B1(n_886),
.B2(n_873),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1348),
.B(n_947),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1430),
.Y(n_1742)
);

NAND2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1440),
.B(n_888),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1333),
.B(n_950),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1375),
.A2(n_994),
.B1(n_995),
.B2(n_993),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1515),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_SL g1747 ( 
.A(n_1451),
.B(n_954),
.C(n_953),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1364),
.B(n_957),
.Y(n_1748)
);

BUFx8_ASAP7_75t_L g1749 ( 
.A(n_1443),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1405),
.B(n_889),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1462),
.B(n_960),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1304),
.B(n_894),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1536),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1366),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1330),
.B(n_897),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1335),
.B(n_906),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1516),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1306),
.A2(n_992),
.B1(n_915),
.B2(n_916),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1340),
.B(n_907),
.Y(n_1759)
);

BUFx8_ASAP7_75t_L g1760 ( 
.A(n_1444),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1484),
.B(n_988),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1525),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1486),
.B(n_641),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1530),
.Y(n_1764)
);

INVx5_ASAP7_75t_L g1765 ( 
.A(n_1441),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1526),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1449),
.B(n_917),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1383),
.A2(n_932),
.B1(n_937),
.B2(n_923),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1338),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1490),
.B(n_1491),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_L g1771 ( 
.A(n_1461),
.B(n_1500),
.C(n_1499),
.Y(n_1771)
);

NAND2x1p5_ASAP7_75t_L g1772 ( 
.A(n_1365),
.B(n_949),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1456),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1423),
.Y(n_1774)
);

AND2x6_ASAP7_75t_SL g1775 ( 
.A(n_1401),
.B(n_958),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1435),
.Y(n_1776)
);

AO22x1_ASAP7_75t_L g1777 ( 
.A1(n_1417),
.A2(n_964),
.B1(n_973),
.B2(n_962),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1448),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1517),
.A2(n_979),
.B1(n_974),
.B2(n_769),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_R g1780 ( 
.A(n_1392),
.B(n_641),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1400),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1486),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1512),
.B(n_641),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1376),
.B(n_641),
.Y(n_1784)
);

AND3x2_ASAP7_75t_SL g1785 ( 
.A(n_1447),
.B(n_20),
.C(n_22),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1455),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1320),
.B(n_769),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1360),
.B(n_769),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1435),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1458),
.B(n_776),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1421),
.B(n_776),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1425),
.B(n_776),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1445),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1324),
.B(n_776),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1431),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1353),
.B(n_795),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1468),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1310),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1466),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1299),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1302),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1467),
.B(n_795),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1473),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1382),
.B(n_795),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1386),
.B(n_795),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1388),
.B(n_817),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1475),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1389),
.B(n_817),
.Y(n_1808)
);

NOR2x2_ASAP7_75t_L g1809 ( 
.A(n_1426),
.B(n_24),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1402),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1403),
.B(n_817),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1418),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1454),
.B(n_1463),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1474),
.Y(n_1814)
);

OR2x4_ASAP7_75t_L g1815 ( 
.A(n_1411),
.B(n_846),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1448),
.Y(n_1816)
);

INVx3_ASAP7_75t_SL g1817 ( 
.A(n_1471),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1422),
.Y(n_1818)
);

CKINVDCx6p67_ASAP7_75t_R g1819 ( 
.A(n_1471),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1377),
.A2(n_1393),
.B1(n_846),
.B2(n_893),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1471),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1434),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1471),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1498),
.B(n_846),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1300),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1298),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1313),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1281),
.A2(n_846),
.B1(n_893),
.B2(n_859),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1369),
.Y(n_1829)
);

AO21x1_ASAP7_75t_L g1830 ( 
.A1(n_1776),
.A2(n_1789),
.B(n_1787),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1739),
.A2(n_1759),
.B(n_1756),
.C(n_1633),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1638),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1552),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1698),
.B(n_1700),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1769),
.A2(n_893),
.B(n_859),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1687),
.B(n_859),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1679),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1638),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1810),
.B(n_893),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1709),
.A2(n_444),
.B(n_443),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1655),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_R g1842 ( 
.A(n_1571),
.B(n_25),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1689),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_SL g1844 ( 
.A1(n_1554),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1733),
.B(n_30),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1546),
.B(n_1571),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1543),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1812),
.B(n_31),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1738),
.B(n_33),
.Y(n_1849)
);

NAND2xp33_ASAP7_75t_L g1850 ( 
.A(n_1817),
.B(n_456),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1553),
.A2(n_459),
.B(n_458),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1543),
.B(n_34),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1548),
.A2(n_465),
.B(n_460),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1606),
.B(n_34),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_SL g1855 ( 
.A(n_1615),
.B(n_467),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1826),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1551),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1667),
.Y(n_1858)
);

O2A1O1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1688),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1829),
.A2(n_471),
.B(n_469),
.Y(n_1860)
);

OR2x6_ASAP7_75t_L g1861 ( 
.A(n_1554),
.B(n_35),
.Y(n_1861)
);

BUFx8_ASAP7_75t_L g1862 ( 
.A(n_1599),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1601),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1612),
.B(n_36),
.Y(n_1864)
);

INVx3_ASAP7_75t_SL g1865 ( 
.A(n_1566),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1826),
.B(n_1705),
.Y(n_1866)
);

NAND2x1p5_ASAP7_75t_L g1867 ( 
.A(n_1655),
.B(n_37),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1557),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1655),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1589),
.B(n_38),
.C(n_39),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1717),
.A2(n_475),
.B(n_474),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1825),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1719),
.A2(n_1723),
.B(n_1721),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1713),
.B(n_1715),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1577),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1815),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1676),
.A2(n_1677),
.B1(n_1617),
.B2(n_1685),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1559),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1564),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1581),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1563),
.B(n_1558),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1587),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1605),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1819),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1730),
.A2(n_480),
.B(n_476),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1574),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1608),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1667),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1669),
.B(n_1622),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1597),
.B(n_46),
.Y(n_1890)
);

BUFx8_ASAP7_75t_SL g1891 ( 
.A(n_1654),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1561),
.B(n_46),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1620),
.B(n_47),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_SL g1894 ( 
.A1(n_1790),
.A2(n_1802),
.B(n_1707),
.C(n_1664),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1592),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1568),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1593),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1788),
.A2(n_487),
.B(n_482),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1634),
.B(n_47),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1781),
.B(n_48),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1675),
.B(n_48),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1591),
.B(n_49),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1617),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1795),
.B(n_49),
.Y(n_1904)
);

NOR3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1668),
.B(n_50),
.C(n_51),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1570),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1542),
.B(n_1710),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1602),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1555),
.B(n_1544),
.Y(n_1909)
);

A2O1A1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1803),
.A2(n_55),
.B(n_52),
.C(n_53),
.Y(n_1910)
);

NOR2x1_ASAP7_75t_SL g1911 ( 
.A(n_1615),
.B(n_53),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_R g1912 ( 
.A(n_1596),
.B(n_56),
.Y(n_1912)
);

O2A1O1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1547),
.A2(n_1755),
.B(n_1584),
.C(n_1590),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1771),
.B(n_57),
.Y(n_1914)
);

A2O1A1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1807),
.A2(n_60),
.B(n_57),
.C(n_59),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1613),
.B(n_1540),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1580),
.B(n_61),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1565),
.B(n_61),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1581),
.Y(n_1919)
);

CKINVDCx8_ASAP7_75t_R g1920 ( 
.A(n_1775),
.Y(n_1920)
);

OAI21xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1602),
.A2(n_62),
.B(n_64),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1761),
.B(n_65),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1767),
.B(n_65),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1597),
.B(n_66),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1588),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1767),
.B(n_67),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1604),
.Y(n_1927)
);

O2A1O1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1586),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1569),
.B(n_1621),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1637),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1636),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1650),
.B(n_73),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1641),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1588),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1646),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1604),
.B(n_75),
.Y(n_1936)
);

CKINVDCx20_ASAP7_75t_R g1937 ( 
.A(n_1671),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1618),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1821),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1539),
.B(n_1575),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1614),
.Y(n_1941)
);

OAI21xp33_ASAP7_75t_L g1942 ( 
.A1(n_1686),
.A2(n_76),
.B(n_77),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1614),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1631),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1631),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1827),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1650),
.B(n_81),
.Y(n_1947)
);

AO21x1_ASAP7_75t_L g1948 ( 
.A1(n_1619),
.A2(n_494),
.B(n_491),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1640),
.A2(n_1792),
.B(n_1791),
.Y(n_1949)
);

OR2x6_ASAP7_75t_L g1950 ( 
.A(n_1635),
.B(n_82),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1652),
.B(n_82),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1658),
.B(n_83),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1648),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1636),
.Y(n_1954)
);

AND2x6_ASAP7_75t_L g1955 ( 
.A(n_1823),
.B(n_86),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1585),
.Y(n_1956)
);

NOR3xp33_ASAP7_75t_L g1957 ( 
.A(n_1747),
.B(n_87),
.C(n_88),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1660),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1659),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1773),
.B(n_89),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1670),
.B(n_90),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_R g1962 ( 
.A(n_1562),
.B(n_90),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1556),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1595),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1964)
);

INVx6_ASAP7_75t_L g1965 ( 
.A(n_1749),
.Y(n_1965)
);

NOR3xp33_ASAP7_75t_SL g1966 ( 
.A(n_1714),
.B(n_93),
.C(n_95),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1821),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1666),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1806),
.Y(n_1969)
);

OR2x6_ASAP7_75t_L g1970 ( 
.A(n_1731),
.B(n_96),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1740),
.A2(n_1768),
.B1(n_1824),
.B2(n_1696),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1816),
.A2(n_1758),
.B1(n_1541),
.B2(n_1818),
.Y(n_1972)
);

A2O1A1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1784),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1545),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1735),
.B(n_98),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1749),
.Y(n_1976)
);

A2O1A1Ixp33_ASAP7_75t_SL g1977 ( 
.A1(n_1820),
.A2(n_1828),
.B(n_1567),
.C(n_1582),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1616),
.A2(n_1734),
.B1(n_1632),
.B2(n_1706),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1690),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1690),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1793),
.B(n_99),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1760),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1616),
.B(n_100),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1632),
.B(n_101),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1681),
.B(n_102),
.Y(n_1985)
);

NOR3xp33_ASAP7_75t_L g1986 ( 
.A(n_1712),
.B(n_102),
.C(n_103),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1798),
.A2(n_501),
.B(n_499),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1797),
.B(n_103),
.Y(n_1988)
);

O2A1O1Ixp33_ASAP7_75t_SL g1989 ( 
.A1(n_1822),
.A2(n_503),
.B(n_507),
.C(n_502),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1706),
.B(n_106),
.Y(n_1990)
);

INVx5_ASAP7_75t_L g1991 ( 
.A(n_1594),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1798),
.A2(n_510),
.B(n_508),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1624),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1764),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1691),
.A2(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1624),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1805),
.A2(n_1811),
.B(n_1808),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1754),
.B(n_108),
.Y(n_1998)
);

A2O1A1Ixp33_ASAP7_75t_L g1999 ( 
.A1(n_1764),
.A2(n_1766),
.B(n_1651),
.C(n_1573),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1732),
.A2(n_515),
.B(n_514),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1760),
.Y(n_2001)
);

INVx6_ASAP7_75t_L g2002 ( 
.A(n_1765),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1693),
.Y(n_2003)
);

A2O1A1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1609),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_2004)
);

OAI22x1_ASAP7_75t_L g2005 ( 
.A1(n_1729),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1746),
.A2(n_117),
.B(n_118),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_SL g2007 ( 
.A(n_1594),
.B(n_517),
.Y(n_2007)
);

O2A1O1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1741),
.A2(n_120),
.B(n_117),
.C(n_119),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1708),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1610),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1607),
.B(n_122),
.Y(n_2011)
);

INVx1_ASAP7_75t_SL g2012 ( 
.A(n_1653),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1560),
.B(n_122),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1653),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1672),
.B(n_123),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1779),
.A2(n_126),
.B(n_123),
.C(n_125),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1678),
.B(n_126),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1680),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1665),
.B(n_127),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1576),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1693),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1665),
.B(n_128),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1736),
.Y(n_2023)
);

O2A1O1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1623),
.A2(n_1627),
.B(n_1630),
.C(n_1626),
.Y(n_2024)
);

INVx6_ASAP7_75t_L g2025 ( 
.A(n_1765),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1745),
.B(n_1657),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1716),
.A2(n_1786),
.B(n_1644),
.C(n_1645),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_1699),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1770),
.B(n_132),
.Y(n_2029)
);

INVx4_ASAP7_75t_L g2030 ( 
.A(n_1567),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1549),
.Y(n_2031)
);

O2A1O1Ixp33_ASAP7_75t_SL g2032 ( 
.A1(n_1763),
.A2(n_1611),
.B(n_1804),
.C(n_1796),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1697),
.Y(n_2033)
);

A2O1A1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1643),
.A2(n_135),
.B(n_132),
.C(n_133),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1695),
.B(n_1751),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1750),
.B(n_137),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1657),
.B(n_138),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1750),
.B(n_139),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1694),
.A2(n_525),
.B(n_524),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1697),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1598),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_2041)
);

INVx8_ASAP7_75t_L g2042 ( 
.A(n_1729),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1549),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1748),
.A2(n_527),
.B(n_526),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1684),
.A2(n_531),
.B(n_528),
.Y(n_2045)
);

O2A1O1Ixp33_ASAP7_75t_L g2046 ( 
.A1(n_1673),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1628),
.A2(n_1647),
.B(n_1642),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1656),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1783),
.Y(n_2049)
);

CKINVDCx8_ASAP7_75t_R g2050 ( 
.A(n_1729),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1662),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1752),
.B(n_145),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1692),
.A2(n_533),
.B(n_532),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_SL g2054 ( 
.A(n_1649),
.B(n_146),
.C(n_147),
.Y(n_2054)
);

NAND3xp33_ASAP7_75t_SL g2055 ( 
.A(n_1744),
.B(n_148),
.C(n_149),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1704),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1772),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1765),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1674),
.B(n_151),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1718),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1703),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1674),
.B(n_1753),
.Y(n_2062)
);

BUFx4f_ASAP7_75t_L g2063 ( 
.A(n_1743),
.Y(n_2063)
);

OAI21xp33_ASAP7_75t_SL g2064 ( 
.A1(n_1702),
.A2(n_152),
.B(n_153),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1701),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1780),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1752),
.B(n_152),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1800),
.B(n_153),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1583),
.A2(n_156),
.B(n_157),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1725),
.Y(n_2070)
);

AND3x2_ASAP7_75t_L g2071 ( 
.A(n_1809),
.B(n_158),
.C(n_159),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1731),
.Y(n_2072)
);

NAND3xp33_ASAP7_75t_SL g2073 ( 
.A(n_1639),
.B(n_160),
.C(n_161),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1814),
.A2(n_163),
.B1(n_160),
.B2(n_162),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1682),
.B(n_162),
.Y(n_2075)
);

A2O1A1Ixp33_ASAP7_75t_L g2076 ( 
.A1(n_1683),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_2076)
);

INVx8_ASAP7_75t_L g2077 ( 
.A(n_1594),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1661),
.B(n_167),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1703),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1737),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1727),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_R g2082 ( 
.A(n_1724),
.B(n_168),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1742),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_SL g2084 ( 
.A(n_1572),
.B(n_168),
.C(n_169),
.Y(n_2084)
);

CKINVDCx16_ASAP7_75t_R g2085 ( 
.A(n_1550),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1762),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1663),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1576),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1726),
.B(n_170),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1785),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1720),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1814),
.Y(n_2092)
);

NOR3xp33_ASAP7_75t_SL g2093 ( 
.A(n_1603),
.B(n_173),
.C(n_175),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1801),
.B(n_175),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1814),
.A2(n_1757),
.B1(n_1600),
.B2(n_1578),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1794),
.Y(n_2096)
);

INVx6_ASAP7_75t_L g2097 ( 
.A(n_1724),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1757),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1711),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1578),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_R g2101 ( 
.A(n_1625),
.B(n_1579),
.Y(n_2101)
);

BUFx8_ASAP7_75t_L g2102 ( 
.A(n_1794),
.Y(n_2102)
);

BUFx12f_ASAP7_75t_L g2103 ( 
.A(n_1722),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_1629),
.A2(n_1711),
.B1(n_1728),
.B2(n_1799),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1625),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1799),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1711),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1777),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_2108)
);

BUFx8_ASAP7_75t_L g2109 ( 
.A(n_1625),
.Y(n_2109)
);

O2A1O1Ixp33_ASAP7_75t_SL g2110 ( 
.A1(n_1782),
.A2(n_541),
.B(n_543),
.C(n_540),
.Y(n_2110)
);

NOR3xp33_ASAP7_75t_L g2111 ( 
.A(n_1782),
.B(n_179),
.C(n_180),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1728),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1728),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1625),
.B(n_181),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1594),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1778),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1600),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_1698),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1813),
.A2(n_553),
.B(n_551),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1813),
.A2(n_555),
.B(n_554),
.Y(n_2120)
);

NAND3xp33_ASAP7_75t_SL g2121 ( 
.A(n_1577),
.B(n_183),
.C(n_186),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1553),
.Y(n_2122)
);

INVxp67_ASAP7_75t_SL g2123 ( 
.A(n_1551),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_1552),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1679),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1813),
.A2(n_561),
.B(n_560),
.Y(n_2126)
);

A2O1A1Ixp33_ASAP7_75t_L g2127 ( 
.A1(n_1633),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1698),
.B(n_188),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1698),
.B(n_189),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1606),
.B(n_189),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1739),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2131)
);

INVx1_ASAP7_75t_SL g2132 ( 
.A(n_1540),
.Y(n_2132)
);

BUFx2_ASAP7_75t_L g2133 ( 
.A(n_1552),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1698),
.B(n_192),
.Y(n_2134)
);

NAND2xp33_ASAP7_75t_SL g2135 ( 
.A(n_1615),
.B(n_194),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1698),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_2136)
);

O2A1O1Ixp33_ASAP7_75t_L g2137 ( 
.A1(n_1739),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1606),
.B(n_198),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1679),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1542),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_1540),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1698),
.B(n_204),
.Y(n_2142)
);

INVx3_ASAP7_75t_L g2143 ( 
.A(n_1655),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1542),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1655),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_1698),
.A2(n_209),
.B1(n_206),
.B2(n_208),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1542),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_1660),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1563),
.B(n_212),
.Y(n_2149)
);

NOR3xp33_ASAP7_75t_L g2150 ( 
.A(n_1589),
.B(n_213),
.C(n_214),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1553),
.Y(n_2151)
);

NOR2x1_ASAP7_75t_L g2152 ( 
.A(n_1654),
.B(n_215),
.Y(n_2152)
);

AOI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_1813),
.A2(n_574),
.B(n_570),
.Y(n_2153)
);

A2O1A1Ixp33_ASAP7_75t_SL g2154 ( 
.A1(n_1633),
.A2(n_580),
.B(n_583),
.C(n_578),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1606),
.B(n_215),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_R g2156 ( 
.A(n_1577),
.B(n_216),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1698),
.B(n_216),
.Y(n_2157)
);

CKINVDCx8_ASAP7_75t_R g2158 ( 
.A(n_1554),
.Y(n_2158)
);

O2A1O1Ixp33_ASAP7_75t_L g2159 ( 
.A1(n_1739),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_2159)
);

A2O1A1Ixp33_ASAP7_75t_SL g2160 ( 
.A1(n_1633),
.A2(n_589),
.B(n_593),
.C(n_588),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_1571),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1698),
.B(n_219),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1698),
.B(n_221),
.Y(n_2163)
);

AOI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_1660),
.A2(n_225),
.B1(n_221),
.B2(n_222),
.Y(n_2164)
);

BUFx12f_ASAP7_75t_L g2165 ( 
.A(n_1599),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_1552),
.Y(n_2166)
);

O2A1O1Ixp33_ASAP7_75t_L g2167 ( 
.A1(n_1739),
.A2(n_229),
.B(n_222),
.C(n_226),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1698),
.B(n_230),
.Y(n_2168)
);

NAND2x1p5_ASAP7_75t_L g2169 ( 
.A(n_1546),
.B(n_230),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1553),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1679),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1655),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_1606),
.B(n_232),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_1552),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_1660),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1552),
.Y(n_2176)
);

OAI21xp33_ASAP7_75t_SL g2177 ( 
.A1(n_1698),
.A2(n_233),
.B(n_234),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_1552),
.Y(n_2178)
);

BUFx12f_ASAP7_75t_L g2179 ( 
.A(n_1599),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1698),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_1660),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_1660),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1698),
.B(n_240),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1679),
.Y(n_2184)
);

AO31x2_ASAP7_75t_L g2185 ( 
.A1(n_1774),
.A2(n_241),
.A3(n_242),
.B(n_243),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1553),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1606),
.B(n_243),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1546),
.B(n_244),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_1810),
.B(n_244),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_R g2190 ( 
.A(n_1571),
.B(n_245),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1679),
.Y(n_2191)
);

O2A1O1Ixp33_ASAP7_75t_L g2192 ( 
.A1(n_1739),
.A2(n_245),
.B(n_247),
.C(n_248),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1679),
.Y(n_2193)
);

NOR3xp33_ASAP7_75t_SL g2194 ( 
.A(n_1668),
.B(n_248),
.C(n_249),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_1552),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1553),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1553),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_1552),
.Y(n_2198)
);

A2O1A1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_1633),
.A2(n_249),
.B(n_250),
.C(n_251),
.Y(n_2199)
);

A2O1A1Ixp33_ASAP7_75t_L g2200 ( 
.A1(n_1633),
.A2(n_252),
.B(n_253),
.C(n_254),
.Y(n_2200)
);

AOI221xp5_ASAP7_75t_L g2201 ( 
.A1(n_1688),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.C(n_259),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1679),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1679),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1698),
.B(n_259),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_1660),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1553),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1810),
.B(n_261),
.Y(n_2207)
);

AO32x1_ASAP7_75t_L g2208 ( 
.A1(n_1774),
.A2(n_262),
.A3(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1679),
.Y(n_2209)
);

A2O1A1Ixp33_ASAP7_75t_SL g2210 ( 
.A1(n_1633),
.A2(n_625),
.B(n_622),
.C(n_621),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_1606),
.B(n_263),
.Y(n_2211)
);

NAND3xp33_ASAP7_75t_SL g2212 ( 
.A(n_1577),
.B(n_264),
.C(n_266),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_1552),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1856),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1940),
.B(n_267),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1837),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2125),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_1881),
.B(n_267),
.Y(n_2218)
);

OAI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_1913),
.A2(n_268),
.B(n_269),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2132),
.B(n_270),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_1939),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1903),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2139),
.Y(n_2223)
);

AO21x2_ASAP7_75t_L g2224 ( 
.A1(n_1830),
.A2(n_608),
.B(n_607),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1907),
.B(n_271),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2132),
.Y(n_2226)
);

AO21x2_ASAP7_75t_L g2227 ( 
.A1(n_1997),
.A2(n_612),
.B(n_609),
.Y(n_2227)
);

AO21x2_ASAP7_75t_L g2228 ( 
.A1(n_1949),
.A2(n_619),
.B(n_618),
.Y(n_2228)
);

AOI22x1_ASAP7_75t_L g2229 ( 
.A1(n_2039),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1834),
.B(n_273),
.Y(n_2230)
);

AO21x2_ASAP7_75t_L g2231 ( 
.A1(n_2101),
.A2(n_620),
.B(n_274),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_1927),
.B(n_275),
.Y(n_2232)
);

AO21x2_ASAP7_75t_L g2233 ( 
.A1(n_1999),
.A2(n_275),
.B(n_277),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_1938),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2171),
.Y(n_2235)
);

AOI22x1_ASAP7_75t_L g2236 ( 
.A1(n_2044),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2184),
.Y(n_2237)
);

INVx5_ASAP7_75t_L g2238 ( 
.A(n_2077),
.Y(n_2238)
);

OAI21x1_ASAP7_75t_L g2239 ( 
.A1(n_2095),
.A2(n_281),
.B(n_283),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1953),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2141),
.B(n_284),
.Y(n_2241)
);

OAI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_1831),
.A2(n_1873),
.B(n_2027),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_1896),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1941),
.Y(n_2244)
);

OA21x2_ASAP7_75t_L g2245 ( 
.A1(n_1948),
.A2(n_285),
.B(n_286),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1979),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_2095),
.A2(n_286),
.B(n_287),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1939),
.Y(n_2248)
);

INVx4_ASAP7_75t_L g2249 ( 
.A(n_2077),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1841),
.Y(n_2250)
);

AO21x2_ASAP7_75t_L g2251 ( 
.A1(n_2154),
.A2(n_287),
.B(n_288),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1980),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_2042),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1994),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1861),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1861),
.B(n_289),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1884),
.B(n_418),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2035),
.B(n_290),
.Y(n_2258)
);

BUFx2_ASAP7_75t_L g2259 ( 
.A(n_1861),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_1884),
.B(n_418),
.Y(n_2260)
);

OAI21x1_ASAP7_75t_SL g2261 ( 
.A1(n_1911),
.A2(n_290),
.B(n_291),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2191),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2141),
.Y(n_2263)
);

AO21x2_ASAP7_75t_L g2264 ( 
.A1(n_2160),
.A2(n_291),
.B(n_292),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1878),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2193),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1886),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2012),
.B(n_294),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1967),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_1879),
.Y(n_2270)
);

BUFx2_ASAP7_75t_SL g2271 ( 
.A(n_1937),
.Y(n_2271)
);

BUFx2_ASAP7_75t_SL g2272 ( 
.A(n_2158),
.Y(n_2272)
);

NOR2x1_ASAP7_75t_R g2273 ( 
.A(n_2165),
.B(n_295),
.Y(n_2273)
);

NOR2xp67_ASAP7_75t_SL g2274 ( 
.A(n_2179),
.B(n_295),
.Y(n_2274)
);

AO21x2_ASAP7_75t_L g2275 ( 
.A1(n_2210),
.A2(n_296),
.B(n_297),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2122),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2202),
.Y(n_2277)
);

AOI22x1_ASAP7_75t_L g2278 ( 
.A1(n_2105),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_2278)
);

OAI21x1_ASAP7_75t_SL g2279 ( 
.A1(n_1876),
.A2(n_299),
.B(n_301),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_1898),
.A2(n_302),
.B(n_303),
.Y(n_2280)
);

AO21x2_ASAP7_75t_L g2281 ( 
.A1(n_1977),
.A2(n_302),
.B(n_303),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1967),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2203),
.Y(n_2283)
);

CKINVDCx20_ASAP7_75t_R g2284 ( 
.A(n_1862),
.Y(n_2284)
);

OAI21x1_ASAP7_75t_L g2285 ( 
.A1(n_1835),
.A2(n_304),
.B(n_305),
.Y(n_2285)
);

AOI22x1_ASAP7_75t_L g2286 ( 
.A1(n_1840),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_2012),
.B(n_306),
.Y(n_2287)
);

OAI21x1_ASAP7_75t_SL g2288 ( 
.A1(n_1876),
.A2(n_309),
.B(n_311),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2124),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_2145),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2209),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2014),
.B(n_311),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1868),
.Y(n_2293)
);

BUFx2_ASAP7_75t_SL g2294 ( 
.A(n_1982),
.Y(n_2294)
);

NAND2x1p5_ASAP7_75t_L g2295 ( 
.A(n_1991),
.B(n_312),
.Y(n_2295)
);

OAI21x1_ASAP7_75t_SL g2296 ( 
.A1(n_1972),
.A2(n_312),
.B(n_313),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_L g2297 ( 
.A(n_2077),
.B(n_313),
.Y(n_2297)
);

BUFx4_ASAP7_75t_SL g2298 ( 
.A(n_1832),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2151),
.Y(n_2299)
);

AO21x2_ASAP7_75t_L g2300 ( 
.A1(n_1836),
.A2(n_314),
.B(n_315),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_1833),
.Y(n_2301)
);

INVx4_ASAP7_75t_L g2302 ( 
.A(n_2042),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2170),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2133),
.Y(n_2304)
);

OAI21x1_ASAP7_75t_L g2305 ( 
.A1(n_1987),
.A2(n_1992),
.B(n_2045),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2024),
.A2(n_314),
.B(n_317),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2186),
.Y(n_2307)
);

INVx6_ASAP7_75t_L g2308 ( 
.A(n_1862),
.Y(n_2308)
);

OA21x2_ASAP7_75t_L g2309 ( 
.A1(n_2069),
.A2(n_319),
.B(n_320),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1872),
.Y(n_2310)
);

BUFx3_ASAP7_75t_L g2311 ( 
.A(n_2102),
.Y(n_2311)
);

INVx1_ASAP7_75t_SL g2312 ( 
.A(n_2176),
.Y(n_2312)
);

BUFx2_ASAP7_75t_R g2313 ( 
.A(n_1838),
.Y(n_2313)
);

BUFx5_ASAP7_75t_L g2314 ( 
.A(n_1955),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1882),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2102),
.Y(n_2316)
);

AO21x2_ASAP7_75t_L g2317 ( 
.A1(n_2069),
.A2(n_320),
.B(n_322),
.Y(n_2317)
);

BUFx4_ASAP7_75t_SL g2318 ( 
.A(n_1976),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2196),
.Y(n_2319)
);

OAI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2119),
.A2(n_323),
.B(n_325),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1874),
.B(n_323),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_1909),
.A2(n_327),
.B(n_328),
.Y(n_2322)
);

AOI22x1_ASAP7_75t_L g2323 ( 
.A1(n_2120),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_2323)
);

HB1xp67_ASAP7_75t_L g2324 ( 
.A(n_2174),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2014),
.B(n_330),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2126),
.A2(n_331),
.B(n_332),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1894),
.A2(n_332),
.B(n_333),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1866),
.B(n_333),
.Y(n_2328)
);

NAND2x1p5_ASAP7_75t_L g2329 ( 
.A(n_1991),
.B(n_334),
.Y(n_2329)
);

OA21x2_ASAP7_75t_L g2330 ( 
.A1(n_1942),
.A2(n_334),
.B(n_335),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1883),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2195),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2042),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2198),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2197),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_1887),
.B(n_336),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2090),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1906),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2062),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_1991),
.Y(n_2340)
);

AO21x2_ASAP7_75t_L g2341 ( 
.A1(n_1852),
.A2(n_343),
.B(n_344),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_2103),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2002),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_2178),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2206),
.Y(n_2345)
);

INVx5_ASAP7_75t_L g2346 ( 
.A(n_1955),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2062),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1895),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_2063),
.Y(n_2349)
);

OAI21x1_ASAP7_75t_SL g2350 ( 
.A1(n_1972),
.A2(n_343),
.B(n_345),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_1963),
.Y(n_2351)
);

AO21x2_ASAP7_75t_L g2352 ( 
.A1(n_1936),
.A2(n_345),
.B(n_346),
.Y(n_2352)
);

BUFx3_ASAP7_75t_L g2353 ( 
.A(n_2002),
.Y(n_2353)
);

OAI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_1877),
.A2(n_2075),
.B(n_1971),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2025),
.Y(n_2355)
);

BUFx2_ASAP7_75t_SL g2356 ( 
.A(n_2001),
.Y(n_2356)
);

INVx1_ASAP7_75t_SL g2357 ( 
.A(n_1946),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2081),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1897),
.Y(n_2359)
);

AO21x2_ASAP7_75t_L g2360 ( 
.A1(n_2078),
.A2(n_347),
.B(n_348),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1959),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_1889),
.B(n_348),
.Y(n_2362)
);

INVx6_ASAP7_75t_L g2363 ( 
.A(n_2025),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2097),
.Y(n_2364)
);

NAND2x1p5_ASAP7_75t_L g2365 ( 
.A(n_1846),
.B(n_349),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_1929),
.B(n_349),
.Y(n_2366)
);

BUFx3_ASAP7_75t_L g2367 ( 
.A(n_2097),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1930),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1933),
.Y(n_2369)
);

AO21x2_ASAP7_75t_L g2370 ( 
.A1(n_2073),
.A2(n_352),
.B(n_353),
.Y(n_2370)
);

INVx5_ASAP7_75t_L g2371 ( 
.A(n_1955),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1935),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_1978),
.B(n_353),
.Y(n_2373)
);

NOR2x1_ASAP7_75t_SL g2374 ( 
.A(n_1970),
.B(n_354),
.Y(n_2374)
);

NAND2x1p5_ASAP7_75t_L g2375 ( 
.A(n_2063),
.B(n_354),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2080),
.B(n_355),
.Y(n_2376)
);

OR2x6_ASAP7_75t_L g2377 ( 
.A(n_1970),
.B(n_417),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1877),
.B(n_356),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1845),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_1848),
.Y(n_2380)
);

BUFx3_ASAP7_75t_L g2381 ( 
.A(n_2109),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_1916),
.A2(n_357),
.B1(n_359),
.B2(n_360),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_1880),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_2083),
.Y(n_2384)
);

OAI21x1_ASAP7_75t_L g2385 ( 
.A1(n_2153),
.A2(n_359),
.B(n_361),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1849),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2118),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2051),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_1954),
.Y(n_2389)
);

NAND2x1p5_ASAP7_75t_L g2390 ( 
.A(n_2161),
.B(n_362),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_1857),
.B(n_2026),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2118),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2086),
.B(n_362),
.Y(n_2393)
);

OAI21x1_ASAP7_75t_L g2394 ( 
.A1(n_1851),
.A2(n_1860),
.B(n_1853),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2109),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_1993),
.B(n_364),
.Y(n_2396)
);

AO21x2_ASAP7_75t_L g2397 ( 
.A1(n_2055),
.A2(n_367),
.B(n_368),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_1890),
.B(n_368),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2056),
.Y(n_2399)
);

OA21x2_ASAP7_75t_L g2400 ( 
.A1(n_1871),
.A2(n_369),
.B(n_370),
.Y(n_2400)
);

AO21x2_ASAP7_75t_L g2401 ( 
.A1(n_2068),
.A2(n_370),
.B(n_371),
.Y(n_2401)
);

BUFx2_ASAP7_75t_SL g2402 ( 
.A(n_2050),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1867),
.B(n_371),
.Y(n_2403)
);

AO21x2_ASAP7_75t_L g2404 ( 
.A1(n_2068),
.A2(n_1989),
.B(n_1917),
.Y(n_2404)
);

AO21x2_ASAP7_75t_L g2405 ( 
.A1(n_2128),
.A2(n_374),
.B(n_375),
.Y(n_2405)
);

AOI22x1_ASAP7_75t_L g2406 ( 
.A1(n_2000),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_2406)
);

AO21x2_ASAP7_75t_L g2407 ( 
.A1(n_2129),
.A2(n_378),
.B(n_379),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_1848),
.Y(n_2408)
);

AO21x2_ASAP7_75t_L g2409 ( 
.A1(n_2134),
.A2(n_378),
.B(n_379),
.Y(n_2409)
);

OAI21x1_ASAP7_75t_L g2410 ( 
.A1(n_1885),
.A2(n_380),
.B(n_381),
.Y(n_2410)
);

INVx4_ASAP7_75t_L g2411 ( 
.A(n_1955),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_1890),
.B(n_380),
.Y(n_2412)
);

OAI21x1_ASAP7_75t_L g2413 ( 
.A1(n_1867),
.A2(n_383),
.B(n_384),
.Y(n_2413)
);

AO21x2_ASAP7_75t_L g2414 ( 
.A1(n_2142),
.A2(n_385),
.B(n_386),
.Y(n_2414)
);

BUFx2_ASAP7_75t_SL g2415 ( 
.A(n_1858),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_1850),
.A2(n_385),
.B(n_386),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2136),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_2189),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_1865),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2060),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1891),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2136),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2070),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_1869),
.Y(n_2424)
);

BUFx2_ASAP7_75t_R g2425 ( 
.A(n_1863),
.Y(n_2425)
);

AO21x2_ASAP7_75t_L g2426 ( 
.A1(n_2157),
.A2(n_387),
.B(n_388),
.Y(n_2426)
);

OAI21x1_ASAP7_75t_L g2427 ( 
.A1(n_2115),
.A2(n_391),
.B(n_392),
.Y(n_2427)
);

BUFx2_ASAP7_75t_SL g2428 ( 
.A(n_1888),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_1919),
.Y(n_2429)
);

NAND2x1p5_ASAP7_75t_L g2430 ( 
.A(n_1924),
.B(n_391),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2146),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2146),
.Y(n_2432)
);

AO21x2_ASAP7_75t_L g2433 ( 
.A1(n_2162),
.A2(n_392),
.B(n_393),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2143),
.Y(n_2434)
);

NAND2x1p5_ASAP7_75t_L g2435 ( 
.A(n_1924),
.B(n_394),
.Y(n_2435)
);

CKINVDCx20_ASAP7_75t_R g2436 ( 
.A(n_1842),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_2172),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2189),
.Y(n_2438)
);

AO21x2_ASAP7_75t_L g2439 ( 
.A1(n_2163),
.A2(n_394),
.B(n_395),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_1970),
.Y(n_2440)
);

AOI22x1_ASAP7_75t_L g2441 ( 
.A1(n_2053),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.Y(n_2441)
);

INVx8_ASAP7_75t_L g2442 ( 
.A(n_1950),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2180),
.Y(n_2443)
);

BUFx2_ASAP7_75t_SL g2444 ( 
.A(n_1988),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2180),
.Y(n_2445)
);

CKINVDCx20_ASAP7_75t_R g2446 ( 
.A(n_2190),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2149),
.B(n_2015),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2123),
.B(n_400),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2099),
.A2(n_402),
.B(n_403),
.Y(n_2449)
);

OR2x6_ASAP7_75t_L g2450 ( 
.A(n_2207),
.B(n_404),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_1925),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_1965),
.Y(n_2452)
);

INVx5_ASAP7_75t_L g2453 ( 
.A(n_2020),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2003),
.B(n_404),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_2020),
.Y(n_2455)
);

CKINVDCx11_ASAP7_75t_R g2456 ( 
.A(n_1920),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1843),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_1843),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1908),
.Y(n_2459)
);

INVx4_ASAP7_75t_L g2460 ( 
.A(n_2088),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_1996),
.B(n_416),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1908),
.Y(n_2462)
);

INVx6_ASAP7_75t_L g2463 ( 
.A(n_2030),
.Y(n_2463)
);

OAI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_1971),
.A2(n_405),
.B(n_406),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_1965),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2207),
.Y(n_2466)
);

OA21x2_ASAP7_75t_L g2467 ( 
.A1(n_2034),
.A2(n_405),
.B(n_406),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_1934),
.B(n_407),
.Y(n_2468)
);

BUFx4_ASAP7_75t_SL g2469 ( 
.A(n_1950),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2058),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2048),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1943),
.Y(n_2472)
);

NAND2x1p5_ASAP7_75t_L g2473 ( 
.A(n_2030),
.B(n_408),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_1943),
.Y(n_2474)
);

INVx8_ASAP7_75t_L g2475 ( 
.A(n_1950),
.Y(n_2475)
);

INVxp67_ASAP7_75t_SL g2476 ( 
.A(n_2166),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_1944),
.Y(n_2477)
);

OAI21x1_ASAP7_75t_L g2478 ( 
.A1(n_2112),
.A2(n_408),
.B(n_409),
.Y(n_2478)
);

OAI21x1_ASAP7_75t_L g2479 ( 
.A1(n_2112),
.A2(n_409),
.B(n_411),
.Y(n_2479)
);

AO22x1_ASAP7_75t_L g2480 ( 
.A1(n_2018),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2116),
.Y(n_2481)
);

BUFx2_ASAP7_75t_R g2482 ( 
.A(n_1974),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_L g2483 ( 
.A1(n_2113),
.A2(n_412),
.B(n_414),
.Y(n_2483)
);

OA21x2_ASAP7_75t_L g2484 ( 
.A1(n_2127),
.A2(n_415),
.B(n_2199),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2092),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_1847),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2113),
.A2(n_415),
.B(n_2100),
.Y(n_2487)
);

CKINVDCx20_ASAP7_75t_R g2488 ( 
.A(n_2023),
.Y(n_2488)
);

OR2x6_ASAP7_75t_L g2489 ( 
.A(n_1875),
.B(n_2169),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1847),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_1900),
.B(n_1985),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2059),
.Y(n_2492)
);

OAI21x1_ASAP7_75t_L g2493 ( 
.A1(n_2131),
.A2(n_2159),
.B(n_2137),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2059),
.Y(n_2494)
);

INVx5_ASAP7_75t_L g2495 ( 
.A(n_2065),
.Y(n_2495)
);

INVx1_ASAP7_75t_SL g2496 ( 
.A(n_1962),
.Y(n_2496)
);

BUFx2_ASAP7_75t_L g2497 ( 
.A(n_2213),
.Y(n_2497)
);

BUFx3_ASAP7_75t_L g2498 ( 
.A(n_1931),
.Y(n_2498)
);

BUFx2_ASAP7_75t_L g2499 ( 
.A(n_1945),
.Y(n_2499)
);

NAND2x1p5_ASAP7_75t_L g2500 ( 
.A(n_1839),
.B(n_1864),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2049),
.Y(n_2501)
);

BUFx3_ASAP7_75t_L g2502 ( 
.A(n_2169),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2185),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2168),
.Y(n_2504)
);

BUFx12f_ASAP7_75t_L g2505 ( 
.A(n_1968),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2183),
.Y(n_2506)
);

AO21x2_ASAP7_75t_L g2507 ( 
.A1(n_2204),
.A2(n_1952),
.B(n_1951),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1904),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2021),
.Y(n_2509)
);

OAI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2167),
.A2(n_2192),
.B(n_1947),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2033),
.Y(n_2511)
);

CKINVDCx6p67_ASAP7_75t_R g2512 ( 
.A(n_2085),
.Y(n_2512)
);

BUFx2_ASAP7_75t_SL g2513 ( 
.A(n_1956),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2082),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2072),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2098),
.B(n_2106),
.Y(n_2516)
);

AO21x2_ASAP7_75t_L g2517 ( 
.A1(n_1932),
.A2(n_2110),
.B(n_2111),
.Y(n_2517)
);

AO21x2_ASAP7_75t_L g2518 ( 
.A1(n_1960),
.A2(n_2200),
.B(n_2076),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2040),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_2117),
.Y(n_2520)
);

OAI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2107),
.A2(n_2104),
.B(n_2114),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_1839),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2009),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2061),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2057),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2066),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2185),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2057),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_2079),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2096),
.Y(n_2530)
);

OAI21x1_ASAP7_75t_L g2531 ( 
.A1(n_2188),
.A2(n_2046),
.B(n_1928),
.Y(n_2531)
);

INVx3_ASAP7_75t_L g2532 ( 
.A(n_1969),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2032),
.A2(n_2029),
.B(n_2047),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2293),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2310),
.Y(n_2535)
);

OAI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2450),
.A2(n_2018),
.B1(n_1964),
.B2(n_1918),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2315),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_2284),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2331),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2284),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2377),
.A2(n_1870),
.B1(n_2150),
.B2(n_2211),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2226),
.Y(n_2542)
);

OAI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2354),
.A2(n_2177),
.B(n_1921),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2216),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2217),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2223),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2214),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2411),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2235),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2237),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2262),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2450),
.A2(n_2074),
.B1(n_2087),
.B2(n_2144),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2263),
.B(n_2052),
.Y(n_2553)
);

OA21x2_ASAP7_75t_L g2554 ( 
.A1(n_2503),
.A2(n_2004),
.B(n_2010),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2411),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_2333),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2214),
.Y(n_2557)
);

BUFx4_ASAP7_75t_SL g2558 ( 
.A(n_2465),
.Y(n_2558)
);

OAI22x1_ASAP7_75t_L g2559 ( 
.A1(n_2440),
.A2(n_2028),
.B1(n_2152),
.B2(n_2067),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2266),
.Y(n_2560)
);

CKINVDCx20_ASAP7_75t_R g2561 ( 
.A(n_2488),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2277),
.Y(n_2562)
);

OAI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_2450),
.A2(n_2074),
.B1(n_2140),
.B2(n_2147),
.Y(n_2563)
);

AO21x1_ASAP7_75t_L g2564 ( 
.A1(n_2411),
.A2(n_2297),
.B(n_2464),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2283),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2369),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2377),
.A2(n_2155),
.B1(n_1854),
.B2(n_2187),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2291),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2338),
.Y(n_2569)
);

AO21x2_ASAP7_75t_L g2570 ( 
.A1(n_2242),
.A2(n_1915),
.B(n_1910),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2369),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2348),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2459),
.B(n_1892),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2359),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_SL g2575 ( 
.A1(n_2442),
.A2(n_1844),
.B1(n_2173),
.B2(n_2138),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2308),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2462),
.B(n_1902),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2346),
.B(n_1914),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2368),
.Y(n_2579)
);

CKINVDCx6p67_ASAP7_75t_R g2580 ( 
.A(n_2311),
.Y(n_2580)
);

BUFx3_ASAP7_75t_L g2581 ( 
.A(n_2308),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2372),
.Y(n_2582)
);

OAI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2450),
.A2(n_2108),
.B1(n_2041),
.B2(n_1995),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2377),
.A2(n_2130),
.B1(n_2212),
.B2(n_2121),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2333),
.Y(n_2585)
);

OAI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2377),
.A2(n_2148),
.B1(n_1958),
.B2(n_2164),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2222),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2222),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2533),
.A2(n_2007),
.B(n_1855),
.Y(n_2589)
);

INVx3_ASAP7_75t_SL g2590 ( 
.A(n_2308),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2244),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2265),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2215),
.A2(n_2156),
.B1(n_2201),
.B2(n_2017),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2298),
.Y(n_2594)
);

HB1xp67_ASAP7_75t_L g2595 ( 
.A(n_2263),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2267),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_SL g2597 ( 
.A(n_2311),
.Y(n_2597)
);

INVx6_ASAP7_75t_L g2598 ( 
.A(n_2302),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2244),
.Y(n_2599)
);

NAND2x1p5_ASAP7_75t_L g2600 ( 
.A(n_2302),
.B(n_1893),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2218),
.B(n_1966),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2318),
.Y(n_2602)
);

NAND2x1p5_ASAP7_75t_L g2603 ( 
.A(n_2302),
.B(n_2037),
.Y(n_2603)
);

BUFx2_ASAP7_75t_L g2604 ( 
.A(n_2253),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_SL g2605 ( 
.A1(n_2442),
.A2(n_2006),
.B1(n_2064),
.B2(n_1961),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2267),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2270),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2246),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2215),
.A2(n_1957),
.B1(n_1986),
.B2(n_1922),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2246),
.Y(n_2610)
);

AOI21x1_ASAP7_75t_L g2611 ( 
.A1(n_2527),
.A2(n_1975),
.B(n_2005),
.Y(n_2611)
);

INVx1_ASAP7_75t_SL g2612 ( 
.A(n_2513),
.Y(n_2612)
);

CKINVDCx20_ASAP7_75t_R g2613 ( 
.A(n_2488),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2252),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2252),
.Y(n_2615)
);

AO21x2_ASAP7_75t_L g2616 ( 
.A1(n_2219),
.A2(n_1973),
.B(n_2016),
.Y(n_2616)
);

INVx3_ASAP7_75t_L g2617 ( 
.A(n_2238),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2254),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2440),
.A2(n_2182),
.B1(n_2181),
.B2(n_2175),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2440),
.A2(n_2205),
.B1(n_2093),
.B2(n_2054),
.Y(n_2620)
);

OR2x2_ASAP7_75t_L g2621 ( 
.A(n_2289),
.B(n_1981),
.Y(n_2621)
);

INVx3_ASAP7_75t_L g2622 ( 
.A(n_2238),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2276),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2430),
.A2(n_2084),
.B1(n_2036),
.B2(n_1990),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2254),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2509),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2511),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2519),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2232),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2218),
.B(n_2194),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2419),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2232),
.Y(n_2632)
);

NAND2x1_ASAP7_75t_L g2633 ( 
.A(n_2460),
.B(n_2007),
.Y(n_2633)
);

AO21x1_ASAP7_75t_L g2634 ( 
.A1(n_2297),
.A2(n_2135),
.B(n_2008),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2525),
.A2(n_2013),
.B1(n_2038),
.B2(n_1901),
.Y(n_2635)
);

INVx1_ASAP7_75t_SL g2636 ( 
.A(n_2444),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2270),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2299),
.Y(n_2638)
);

OAI21xp5_ASAP7_75t_SL g2639 ( 
.A1(n_2430),
.A2(n_2071),
.B(n_1859),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2299),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2398),
.B(n_1905),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2232),
.Y(n_2642)
);

OAI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2306),
.A2(n_2378),
.B(n_2387),
.Y(n_2643)
);

NAND2x1p5_ASAP7_75t_L g2644 ( 
.A(n_2238),
.B(n_1912),
.Y(n_2644)
);

BUFx6f_ASAP7_75t_L g2645 ( 
.A(n_2453),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2376),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2412),
.B(n_2091),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2376),
.Y(n_2648)
);

AOI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2528),
.A2(n_2022),
.B1(n_2019),
.B2(n_2011),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2393),
.Y(n_2650)
);

BUFx4f_ASAP7_75t_L g2651 ( 
.A(n_2512),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2419),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_SL g2653 ( 
.A1(n_2442),
.A2(n_2031),
.B1(n_2043),
.B2(n_1984),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2303),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2393),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2442),
.A2(n_2089),
.B1(n_2094),
.B2(n_1926),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2491),
.B(n_1998),
.Y(n_2657)
);

BUFx2_ASAP7_75t_SL g2658 ( 
.A(n_2465),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2316),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2393),
.Y(n_2660)
);

INVx4_ASAP7_75t_SL g2661 ( 
.A(n_2316),
.Y(n_2661)
);

OAI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_2475),
.A2(n_1983),
.B1(n_1923),
.B2(n_1899),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2481),
.Y(n_2663)
);

INVx1_ASAP7_75t_SL g2664 ( 
.A(n_2301),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2253),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2303),
.Y(n_2666)
);

INVxp67_ASAP7_75t_L g2667 ( 
.A(n_2523),
.Y(n_2667)
);

CKINVDCx11_ASAP7_75t_R g2668 ( 
.A(n_2456),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2256),
.B(n_2185),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2307),
.Y(n_2670)
);

OAI21x1_ASAP7_75t_L g2671 ( 
.A1(n_2394),
.A2(n_2208),
.B(n_2305),
.Y(n_2671)
);

INVx1_ASAP7_75t_SL g2672 ( 
.A(n_2301),
.Y(n_2672)
);

INVx4_ASAP7_75t_L g2673 ( 
.A(n_2238),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_2421),
.Y(n_2674)
);

OAI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2435),
.A2(n_2408),
.B1(n_2418),
.B2(n_2380),
.Y(n_2675)
);

AOI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2472),
.A2(n_2486),
.B1(n_2490),
.B2(n_2474),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2220),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2373),
.B(n_2225),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2241),
.Y(n_2679)
);

BUFx4f_ASAP7_75t_SL g2680 ( 
.A(n_2436),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2336),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2307),
.Y(n_2682)
);

CKINVDCx20_ASAP7_75t_R g2683 ( 
.A(n_2421),
.Y(n_2683)
);

INVx3_ASAP7_75t_L g2684 ( 
.A(n_2249),
.Y(n_2684)
);

INVx2_ASAP7_75t_SL g2685 ( 
.A(n_2349),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2319),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2319),
.Y(n_2687)
);

BUFx12f_ASAP7_75t_L g2688 ( 
.A(n_2456),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2392),
.B(n_2417),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2335),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2335),
.Y(n_2691)
);

INVx1_ASAP7_75t_SL g2692 ( 
.A(n_2324),
.Y(n_2692)
);

BUFx2_ASAP7_75t_L g2693 ( 
.A(n_2475),
.Y(n_2693)
);

CKINVDCx20_ASAP7_75t_R g2694 ( 
.A(n_2512),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2249),
.Y(n_2695)
);

INVxp33_ASAP7_75t_L g2696 ( 
.A(n_2358),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2349),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2345),
.Y(n_2698)
);

CKINVDCx11_ASAP7_75t_R g2699 ( 
.A(n_2505),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2475),
.A2(n_2431),
.B1(n_2432),
.B2(n_2422),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2475),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2345),
.Y(n_2702)
);

OAI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_2435),
.A2(n_2259),
.B1(n_2255),
.B2(n_2380),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2361),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2361),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2324),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2515),
.Y(n_2707)
);

INVx4_ASAP7_75t_L g2708 ( 
.A(n_2452),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2388),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2225),
.B(n_2332),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2332),
.B(n_2334),
.Y(n_2711)
);

BUFx4f_ASAP7_75t_SL g2712 ( 
.A(n_2436),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2388),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2399),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2514),
.B(n_2357),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2399),
.Y(n_2716)
);

AND2x4_ASAP7_75t_L g2717 ( 
.A(n_2346),
.B(n_2371),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2443),
.A2(n_2457),
.B1(n_2458),
.B2(n_2445),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2420),
.Y(n_2719)
);

NOR2x1_ASAP7_75t_L g2720 ( 
.A(n_2231),
.B(n_2502),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2334),
.B(n_2366),
.Y(n_2721)
);

INVx4_ASAP7_75t_L g2722 ( 
.A(n_2452),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2420),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2423),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2391),
.A2(n_2408),
.B1(n_2438),
.B2(n_2418),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2493),
.A2(n_2510),
.B(n_2531),
.Y(n_2726)
);

CKINVDCx11_ASAP7_75t_R g2727 ( 
.A(n_2505),
.Y(n_2727)
);

INVx5_ASAP7_75t_L g2728 ( 
.A(n_2453),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2390),
.Y(n_2729)
);

AO21x1_ASAP7_75t_L g2730 ( 
.A1(n_2403),
.A2(n_2473),
.B(n_2329),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2390),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2396),
.Y(n_2732)
);

INVx6_ASAP7_75t_L g2733 ( 
.A(n_2495),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2391),
.A2(n_2438),
.B1(n_2466),
.B2(n_2366),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2501),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2396),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2466),
.A2(n_2447),
.B1(n_2489),
.B2(n_2504),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2396),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2469),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2461),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2339),
.Y(n_2741)
);

INVx4_ASAP7_75t_L g2742 ( 
.A(n_2346),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2249),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2446),
.A2(n_2454),
.B1(n_2494),
.B2(n_2492),
.Y(n_2744)
);

INVx4_ASAP7_75t_SL g2745 ( 
.A(n_2342),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2347),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2489),
.A2(n_2506),
.B1(n_2508),
.B2(n_2386),
.Y(n_2747)
);

OAI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2346),
.A2(n_2371),
.B1(n_2489),
.B2(n_2473),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2461),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_SL g2750 ( 
.A1(n_2374),
.A2(n_2446),
.B1(n_2502),
.B2(n_2288),
.Y(n_2750)
);

HB1xp67_ASAP7_75t_L g2751 ( 
.A(n_2344),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2487),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2453),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2448),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2485),
.Y(n_2755)
);

NAND2x1p5_ASAP7_75t_L g2756 ( 
.A(n_2342),
.B(n_2381),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2485),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2448),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2375),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_SL g2760 ( 
.A1(n_2279),
.A2(n_2371),
.B1(n_2314),
.B2(n_2350),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2375),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2379),
.A2(n_2268),
.B1(n_2287),
.B2(n_2296),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2239),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2497),
.B(n_2476),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2239),
.Y(n_2765)
);

INVx8_ASAP7_75t_L g2766 ( 
.A(n_2495),
.Y(n_2766)
);

OAI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2371),
.A2(n_2329),
.B1(n_2295),
.B2(n_2322),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2313),
.Y(n_2768)
);

CKINVDCx20_ASAP7_75t_R g2769 ( 
.A(n_2234),
.Y(n_2769)
);

INVx2_ASAP7_75t_SL g2770 ( 
.A(n_2381),
.Y(n_2770)
);

INVxp67_ASAP7_75t_L g2771 ( 
.A(n_2272),
.Y(n_2771)
);

OAI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2295),
.A2(n_2337),
.B1(n_2365),
.B2(n_2230),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2337),
.A2(n_2365),
.B1(n_2328),
.B2(n_2268),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2515),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2247),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2454),
.A2(n_2287),
.B1(n_2382),
.B2(n_2480),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2304),
.B(n_2312),
.Y(n_2777)
);

BUFx10_ASAP7_75t_L g2778 ( 
.A(n_2257),
.Y(n_2778)
);

BUFx8_ASAP7_75t_L g2779 ( 
.A(n_2234),
.Y(n_2779)
);

BUFx2_ASAP7_75t_R g2780 ( 
.A(n_2271),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2260),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2260),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_L g2783 ( 
.A1(n_2362),
.A2(n_2258),
.B1(n_2484),
.B2(n_2292),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2260),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2321),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2341),
.Y(n_2786)
);

AOI22xp33_ASAP7_75t_SL g2787 ( 
.A1(n_2314),
.A2(n_2278),
.B1(n_2496),
.B2(n_2395),
.Y(n_2787)
);

AOI222xp33_ASAP7_75t_L g2788 ( 
.A1(n_2536),
.A2(n_2273),
.B1(n_2274),
.B2(n_2395),
.C1(n_2526),
.C2(n_2451),
.Y(n_2788)
);

AOI21xp33_ASAP7_75t_L g2789 ( 
.A1(n_2662),
.A2(n_2518),
.B(n_2484),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2534),
.Y(n_2790)
);

CKINVDCx5p33_ASAP7_75t_R g2791 ( 
.A(n_2594),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2735),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2535),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2537),
.Y(n_2794)
);

CKINVDCx14_ASAP7_75t_R g2795 ( 
.A(n_2561),
.Y(n_2795)
);

OR2x6_ASAP7_75t_L g2796 ( 
.A(n_2602),
.B(n_2294),
.Y(n_2796)
);

NAND2xp33_ASAP7_75t_R g2797 ( 
.A(n_2768),
.B(n_2384),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2547),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2539),
.Y(n_2799)
);

HB1xp67_ASAP7_75t_L g2800 ( 
.A(n_2664),
.Y(n_2800)
);

AND2x2_ASAP7_75t_SL g2801 ( 
.A(n_2651),
.B(n_2340),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_2766),
.Y(n_2802)
);

OAI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2593),
.A2(n_2327),
.B(n_2416),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2544),
.Y(n_2804)
);

NAND2x1_ASAP7_75t_L g2805 ( 
.A(n_2548),
.B(n_2340),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2754),
.B(n_2383),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2711),
.B(n_2470),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2545),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2557),
.Y(n_2809)
);

O2A1O1Ixp5_ASAP7_75t_L g2810 ( 
.A1(n_2564),
.A2(n_2460),
.B(n_2340),
.C(n_2282),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_R g2811 ( 
.A(n_2651),
.B(n_2240),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2536),
.A2(n_2500),
.B1(n_2468),
.B2(n_2463),
.Y(n_2812)
);

AOI22xp33_ASAP7_75t_L g2813 ( 
.A1(n_2586),
.A2(n_2484),
.B1(n_2370),
.B2(n_2397),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2758),
.B(n_2429),
.Y(n_2814)
);

INVx6_ASAP7_75t_L g2815 ( 
.A(n_2745),
.Y(n_2815)
);

HB1xp67_ASAP7_75t_L g2816 ( 
.A(n_2664),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2741),
.B(n_2477),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2548),
.B(n_2453),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2696),
.B(n_2613),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_R g2820 ( 
.A(n_2694),
.B(n_2240),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2746),
.B(n_2477),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2647),
.B(n_2470),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2555),
.B(n_2530),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2546),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_SL g2825 ( 
.A1(n_2739),
.A2(n_2356),
.B1(n_2402),
.B2(n_2482),
.Y(n_2825)
);

NAND2xp33_ASAP7_75t_R g2826 ( 
.A(n_2556),
.B(n_2309),
.Y(n_2826)
);

OAI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2593),
.A2(n_2500),
.B1(n_2495),
.B2(n_2309),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2538),
.B(n_2243),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2657),
.B(n_2325),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2549),
.Y(n_2830)
);

O2A1O1Ixp33_ASAP7_75t_SL g2831 ( 
.A1(n_2748),
.A2(n_2389),
.B(n_2221),
.C(n_2282),
.Y(n_2831)
);

INVxp67_ASAP7_75t_L g2832 ( 
.A(n_2764),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2550),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2766),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2766),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2551),
.Y(n_2836)
);

OR2x2_ASAP7_75t_L g2837 ( 
.A(n_2672),
.B(n_2692),
.Y(n_2837)
);

NAND3xp33_ASAP7_75t_L g2838 ( 
.A(n_2584),
.B(n_2406),
.C(n_2441),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_R g2839 ( 
.A(n_2699),
.B(n_2243),
.Y(n_2839)
);

AOI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2601),
.A2(n_2397),
.B1(n_2370),
.B2(n_2499),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2710),
.B(n_2553),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_SL g2842 ( 
.A1(n_2639),
.A2(n_2389),
.B(n_2248),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2663),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2555),
.B(n_2530),
.Y(n_2844)
);

NAND3xp33_ASAP7_75t_SL g2845 ( 
.A(n_2639),
.B(n_2425),
.C(n_2460),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_L g2846 ( 
.A1(n_2586),
.A2(n_2314),
.B1(n_2518),
.B2(n_2522),
.Y(n_2846)
);

NAND3xp33_ASAP7_75t_L g2847 ( 
.A(n_2575),
.B(n_2236),
.C(n_2229),
.Y(n_2847)
);

NAND2xp33_ASAP7_75t_R g2848 ( 
.A(n_2585),
.B(n_2309),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2668),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2730),
.B(n_2314),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2776),
.A2(n_2463),
.B1(n_2495),
.B2(n_2522),
.Y(n_2851)
);

NAND2xp33_ASAP7_75t_R g2852 ( 
.A(n_2707),
.B(n_2330),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2721),
.B(n_2692),
.Y(n_2853)
);

NAND2xp33_ASAP7_75t_R g2854 ( 
.A(n_2774),
.B(n_2330),
.Y(n_2854)
);

AO21x2_ASAP7_75t_L g2855 ( 
.A1(n_2726),
.A2(n_2231),
.B(n_2281),
.Y(n_2855)
);

AND2x4_ASAP7_75t_L g2856 ( 
.A(n_2617),
.B(n_2530),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2718),
.B(n_2532),
.Y(n_2857)
);

CKINVDCx16_ASAP7_75t_R g2858 ( 
.A(n_2597),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2676),
.B(n_2678),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2560),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2706),
.B(n_2604),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_R g2862 ( 
.A(n_2727),
.B(n_2314),
.Y(n_2862)
);

OR2x6_ASAP7_75t_L g2863 ( 
.A(n_2644),
.B(n_2415),
.Y(n_2863)
);

OR2x6_ASAP7_75t_L g2864 ( 
.A(n_2598),
.B(n_2428),
.Y(n_2864)
);

HB1xp67_ASAP7_75t_L g2865 ( 
.A(n_2607),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2637),
.B(n_2471),
.Y(n_2866)
);

BUFx3_ASAP7_75t_L g2867 ( 
.A(n_2756),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2676),
.B(n_2532),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2562),
.Y(n_2869)
);

OR2x2_ASAP7_75t_L g2870 ( 
.A(n_2595),
.B(n_2520),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2565),
.Y(n_2871)
);

AOI222xp33_ASAP7_75t_L g2872 ( 
.A1(n_2630),
.A2(n_2261),
.B1(n_2498),
.B2(n_2532),
.C1(n_2524),
.C2(n_2529),
.Y(n_2872)
);

OA21x2_ASAP7_75t_L g2873 ( 
.A1(n_2671),
.A2(n_2521),
.B(n_2531),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2568),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_2558),
.Y(n_2875)
);

AO31x2_ASAP7_75t_L g2876 ( 
.A1(n_2763),
.A2(n_2224),
.A3(n_2404),
.B(n_2245),
.Y(n_2876)
);

AO31x2_ASAP7_75t_L g2877 ( 
.A1(n_2765),
.A2(n_2224),
.A3(n_2404),
.B(n_2245),
.Y(n_2877)
);

INVx6_ASAP7_75t_L g2878 ( 
.A(n_2745),
.Y(n_2878)
);

A2O1A1Ixp33_ASAP7_75t_L g2879 ( 
.A1(n_2767),
.A2(n_2413),
.B(n_2449),
.C(n_2478),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2612),
.Y(n_2880)
);

NAND2xp33_ASAP7_75t_SL g2881 ( 
.A(n_2748),
.B(n_2317),
.Y(n_2881)
);

CKINVDCx5p33_ASAP7_75t_R g2882 ( 
.A(n_2688),
.Y(n_2882)
);

OR2x2_ASAP7_75t_L g2883 ( 
.A(n_2542),
.B(n_2520),
.Y(n_2883)
);

OR2x6_ASAP7_75t_L g2884 ( 
.A(n_2598),
.B(n_2364),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2665),
.B(n_2343),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2569),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_2563),
.A2(n_2314),
.B1(n_2522),
.B2(n_2286),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_2580),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2777),
.B(n_2405),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2612),
.B(n_2343),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2641),
.B(n_2353),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2751),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2617),
.B(n_2221),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2566),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2572),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2542),
.B(n_2353),
.Y(n_2896)
);

BUFx3_ASAP7_75t_L g2897 ( 
.A(n_2631),
.Y(n_2897)
);

A2O1A1Ixp33_ASAP7_75t_L g2898 ( 
.A1(n_2767),
.A2(n_2413),
.B(n_2483),
.C(n_2449),
.Y(n_2898)
);

OR2x6_ASAP7_75t_L g2899 ( 
.A(n_2658),
.B(n_2364),
.Y(n_2899)
);

CKINVDCx5p33_ASAP7_75t_R g2900 ( 
.A(n_2597),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2677),
.B(n_2355),
.Y(n_2901)
);

INVx5_ASAP7_75t_L g2902 ( 
.A(n_2728),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_2563),
.A2(n_2314),
.B1(n_2522),
.B2(n_2323),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2574),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2552),
.A2(n_2317),
.B1(n_2467),
.B2(n_2507),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2626),
.B(n_2405),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2579),
.Y(n_2907)
);

OR2x6_ASAP7_75t_L g2908 ( 
.A(n_2540),
.B(n_2367),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2582),
.Y(n_2909)
);

NAND2xp33_ASAP7_75t_R g2910 ( 
.A(n_2693),
.B(n_2467),
.Y(n_2910)
);

BUFx12f_ASAP7_75t_L g2911 ( 
.A(n_2779),
.Y(n_2911)
);

AND2x4_ASAP7_75t_L g2912 ( 
.A(n_2622),
.B(n_2221),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2571),
.Y(n_2913)
);

NAND2xp33_ASAP7_75t_R g2914 ( 
.A(n_2701),
.B(n_2467),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2674),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2673),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2679),
.B(n_2355),
.Y(n_2917)
);

NAND2xp33_ASAP7_75t_R g2918 ( 
.A(n_2622),
.B(n_2400),
.Y(n_2918)
);

CKINVDCx5p33_ASAP7_75t_R g2919 ( 
.A(n_2683),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2627),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2717),
.B(n_2248),
.Y(n_2921)
);

NAND2xp33_ASAP7_75t_R g2922 ( 
.A(n_2684),
.B(n_2400),
.Y(n_2922)
);

CKINVDCx16_ASAP7_75t_R g2923 ( 
.A(n_2708),
.Y(n_2923)
);

NAND2xp33_ASAP7_75t_R g2924 ( 
.A(n_2684),
.B(n_2400),
.Y(n_2924)
);

CKINVDCx16_ASAP7_75t_R g2925 ( 
.A(n_2708),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2776),
.A2(n_2463),
.B1(n_2282),
.B2(n_2269),
.Y(n_2926)
);

INVx4_ASAP7_75t_SL g2927 ( 
.A(n_2590),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2587),
.Y(n_2928)
);

CKINVDCx16_ASAP7_75t_R g2929 ( 
.A(n_2722),
.Y(n_2929)
);

OR2x6_ASAP7_75t_L g2930 ( 
.A(n_2722),
.B(n_2367),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_R g2931 ( 
.A(n_2680),
.B(n_2363),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2552),
.A2(n_2507),
.B1(n_2439),
.B2(n_2409),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2592),
.Y(n_2933)
);

NAND2xp33_ASAP7_75t_R g2934 ( 
.A(n_2695),
.B(n_2248),
.Y(n_2934)
);

HB1xp67_ASAP7_75t_L g2935 ( 
.A(n_2588),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2669),
.B(n_2498),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2628),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2652),
.B(n_2516),
.Y(n_2938)
);

AOI22xp33_ASAP7_75t_L g2939 ( 
.A1(n_2583),
.A2(n_2407),
.B1(n_2433),
.B2(n_2414),
.Y(n_2939)
);

NAND2xp33_ASAP7_75t_R g2940 ( 
.A(n_2695),
.B(n_2269),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2591),
.Y(n_2941)
);

NOR3xp33_ASAP7_75t_SL g2942 ( 
.A(n_2620),
.B(n_2363),
.C(n_2233),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2673),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_R g2944 ( 
.A(n_2712),
.B(n_2363),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2567),
.A2(n_2269),
.B1(n_2524),
.B2(n_2529),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2596),
.Y(n_2946)
);

NAND3xp33_ASAP7_75t_SL g2947 ( 
.A(n_2636),
.B(n_2233),
.C(n_2352),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2599),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_2779),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2744),
.B(n_2407),
.Y(n_2950)
);

A2O1A1Ixp33_ASAP7_75t_L g2951 ( 
.A1(n_2620),
.A2(n_2479),
.B(n_2483),
.C(n_2478),
.Y(n_2951)
);

NOR2x1p5_ASAP7_75t_L g2952 ( 
.A(n_2576),
.B(n_2424),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2608),
.Y(n_2953)
);

CKINVDCx5p33_ASAP7_75t_R g2954 ( 
.A(n_2780),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2610),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_2780),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_2769),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2744),
.B(n_2409),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2583),
.A2(n_2439),
.B1(n_2414),
.B2(n_2433),
.Y(n_2959)
);

OR2x6_ASAP7_75t_L g2960 ( 
.A(n_2733),
.B(n_2479),
.Y(n_2960)
);

NAND2xp33_ASAP7_75t_R g2961 ( 
.A(n_2743),
.B(n_2290),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2685),
.B(n_2516),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2728),
.Y(n_2963)
);

NOR3xp33_ASAP7_75t_SL g2964 ( 
.A(n_2703),
.B(n_2426),
.C(n_2352),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2606),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2614),
.Y(n_2966)
);

INVxp67_ASAP7_75t_L g2967 ( 
.A(n_2715),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2697),
.B(n_2516),
.Y(n_2968)
);

OR2x2_ASAP7_75t_L g2969 ( 
.A(n_2615),
.B(n_2401),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2618),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2625),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_R g2972 ( 
.A(n_2581),
.B(n_2290),
.Y(n_2972)
);

HB1xp67_ASAP7_75t_L g2973 ( 
.A(n_2667),
.Y(n_2973)
);

HB1xp67_ASAP7_75t_L g2974 ( 
.A(n_2682),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2619),
.A2(n_2426),
.B1(n_2341),
.B2(n_2401),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2659),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_2661),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_R g2978 ( 
.A(n_2743),
.B(n_2290),
.Y(n_2978)
);

OAI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2609),
.A2(n_2410),
.B(n_2385),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2623),
.Y(n_2980)
);

HB1xp67_ASAP7_75t_L g2981 ( 
.A(n_2686),
.Y(n_2981)
);

NOR3xp33_ASAP7_75t_SL g2982 ( 
.A(n_2624),
.B(n_2360),
.C(n_2427),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2687),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2621),
.B(n_2770),
.Y(n_2984)
);

BUFx2_ASAP7_75t_L g2985 ( 
.A(n_2733),
.Y(n_2985)
);

CKINVDCx16_ASAP7_75t_R g2986 ( 
.A(n_2778),
.Y(n_2986)
);

NOR3xp33_ASAP7_75t_SL g2987 ( 
.A(n_2624),
.B(n_2360),
.C(n_2427),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2619),
.A2(n_2605),
.B1(n_2541),
.B2(n_2773),
.Y(n_2988)
);

HB1xp67_ASAP7_75t_L g2989 ( 
.A(n_2690),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2661),
.Y(n_2990)
);

BUFx2_ASAP7_75t_SL g2991 ( 
.A(n_2728),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2691),
.Y(n_2992)
);

NAND2xp33_ASAP7_75t_SL g2993 ( 
.A(n_2675),
.B(n_2300),
.Y(n_2993)
);

INVxp67_ASAP7_75t_SL g2994 ( 
.A(n_2675),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2734),
.B(n_2300),
.Y(n_2995)
);

BUFx3_ASAP7_75t_L g2996 ( 
.A(n_2645),
.Y(n_2996)
);

CKINVDCx14_ASAP7_75t_R g2997 ( 
.A(n_2778),
.Y(n_2997)
);

AND2x2_ASAP7_75t_L g2998 ( 
.A(n_2759),
.B(n_2434),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_SL g2999 ( 
.A1(n_2772),
.A2(n_2228),
.B1(n_2227),
.B2(n_2517),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2761),
.B(n_2437),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2928),
.Y(n_3001)
);

NOR2x1_ASAP7_75t_L g3002 ( 
.A(n_2845),
.B(n_2729),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2841),
.B(n_2689),
.Y(n_3003)
);

AOI33xp33_ASAP7_75t_L g3004 ( 
.A1(n_2988),
.A2(n_2750),
.A3(n_2747),
.B1(n_2737),
.B2(n_2653),
.B3(n_2700),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2790),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2793),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2794),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2799),
.Y(n_3008)
);

AND2x4_ASAP7_75t_SL g3009 ( 
.A(n_2802),
.B(n_2834),
.Y(n_3009)
);

HB1xp67_ASAP7_75t_L g3010 ( 
.A(n_2935),
.Y(n_3010)
);

INVx5_ASAP7_75t_L g3011 ( 
.A(n_2902),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2853),
.B(n_2689),
.Y(n_3012)
);

AO21x2_ASAP7_75t_L g3013 ( 
.A1(n_2947),
.A2(n_2726),
.B(n_2786),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2804),
.Y(n_3014)
);

OAI211xp5_ASAP7_75t_L g3015 ( 
.A1(n_2788),
.A2(n_2609),
.B(n_2543),
.C(n_2762),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2808),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2807),
.B(n_2725),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2832),
.B(n_2698),
.Y(n_3018)
);

CKINVDCx14_ASAP7_75t_R g3019 ( 
.A(n_2839),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2837),
.B(n_2704),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2859),
.B(n_2577),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2936),
.B(n_2713),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2829),
.B(n_2714),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2824),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2798),
.Y(n_3025)
);

AND2x2_ASAP7_75t_L g3026 ( 
.A(n_2822),
.B(n_2716),
.Y(n_3026)
);

HB1xp67_ASAP7_75t_L g3027 ( 
.A(n_2974),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2809),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2984),
.B(n_2719),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2895),
.B(n_2577),
.Y(n_3030)
);

INVxp67_ASAP7_75t_SL g3031 ( 
.A(n_2981),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2861),
.B(n_2724),
.Y(n_3032)
);

OR2x2_ASAP7_75t_L g3033 ( 
.A(n_2865),
.B(n_2638),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2830),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2833),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2978),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2904),
.B(n_2573),
.Y(n_3037)
);

NAND2x1p5_ASAP7_75t_SL g3038 ( 
.A(n_2850),
.B(n_2720),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2836),
.Y(n_3039)
);

AND2x2_ASAP7_75t_SL g3040 ( 
.A(n_2835),
.B(n_2717),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2972),
.Y(n_3041)
);

INVx2_ASAP7_75t_R g3042 ( 
.A(n_2902),
.Y(n_3042)
);

HB1xp67_ASAP7_75t_L g3043 ( 
.A(n_2989),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2907),
.B(n_2573),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2894),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2860),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2995),
.B(n_2775),
.Y(n_3047)
);

AND2x4_ASAP7_75t_L g3048 ( 
.A(n_2994),
.B(n_2720),
.Y(n_3048)
);

HB1xp67_ASAP7_75t_L g3049 ( 
.A(n_2800),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2869),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2871),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2874),
.Y(n_3052)
);

NOR2xp67_ASAP7_75t_L g3053 ( 
.A(n_2902),
.B(n_2559),
.Y(n_3053)
);

NOR2x1_ASAP7_75t_SL g3054 ( 
.A(n_2864),
.B(n_2742),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2901),
.B(n_2781),
.Y(n_3055)
);

BUFx2_ASAP7_75t_L g3056 ( 
.A(n_2864),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2917),
.B(n_2782),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2896),
.B(n_2784),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2938),
.B(n_2629),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2891),
.B(n_2632),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2802),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2886),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2920),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2913),
.Y(n_3064)
);

INVxp67_ASAP7_75t_L g3065 ( 
.A(n_2816),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2937),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2880),
.B(n_2642),
.Y(n_3067)
);

BUFx2_ASAP7_75t_L g3068 ( 
.A(n_2862),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2909),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2892),
.Y(n_3070)
);

AOI22xp33_ASAP7_75t_SL g3071 ( 
.A1(n_2812),
.A2(n_2772),
.B1(n_2731),
.B2(n_2648),
.Y(n_3071)
);

INVx3_ASAP7_75t_L g3072 ( 
.A(n_2960),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2933),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2941),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2890),
.B(n_2646),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2948),
.Y(n_3076)
);

HB1xp67_ASAP7_75t_L g3077 ( 
.A(n_2843),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_2916),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_2847),
.A2(n_2634),
.B1(n_2846),
.B2(n_2785),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_2946),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2965),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2897),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2883),
.B(n_2973),
.Y(n_3083)
);

BUFx2_ASAP7_75t_L g3084 ( 
.A(n_2916),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2962),
.B(n_2650),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2968),
.B(n_2655),
.Y(n_3086)
);

OA332x1_ASAP7_75t_L g3087 ( 
.A1(n_2851),
.A2(n_2681),
.A3(n_2649),
.B1(n_2635),
.B2(n_2771),
.B3(n_2783),
.C1(n_2611),
.C2(n_2643),
.Y(n_3087)
);

CKINVDCx6p67_ASAP7_75t_R g3088 ( 
.A(n_2796),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_2866),
.B(n_2640),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2953),
.Y(n_3090)
);

HB1xp67_ASAP7_75t_L g3091 ( 
.A(n_2980),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2955),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2966),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2970),
.B(n_2752),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2813),
.A2(n_2635),
.B1(n_2649),
.B2(n_2643),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2870),
.B(n_2660),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_2817),
.B(n_2654),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2971),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2821),
.B(n_2666),
.Y(n_3099)
);

OAI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_2997),
.A2(n_2787),
.B1(n_2656),
.B2(n_2603),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2960),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2983),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2885),
.B(n_2670),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2838),
.A2(n_2616),
.B1(n_2570),
.B2(n_2578),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2806),
.B(n_2702),
.Y(n_3105)
);

OR2x2_ASAP7_75t_L g3106 ( 
.A(n_2889),
.B(n_2705),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2943),
.Y(n_3107)
);

OAI21xp33_ASAP7_75t_L g3108 ( 
.A1(n_2942),
.A2(n_2760),
.B(n_2749),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_2943),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2814),
.B(n_2709),
.Y(n_3110)
);

HB1xp67_ASAP7_75t_L g3111 ( 
.A(n_2792),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2992),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2976),
.B(n_2723),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2998),
.B(n_2732),
.Y(n_3114)
);

INVx4_ASAP7_75t_SL g3115 ( 
.A(n_2815),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_3000),
.B(n_2736),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2969),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2906),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2840),
.B(n_2738),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_2868),
.B(n_2740),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2967),
.B(n_2755),
.Y(n_3121)
);

INVx3_ASAP7_75t_L g3122 ( 
.A(n_2823),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2857),
.B(n_2757),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2905),
.B(n_2554),
.Y(n_3124)
);

OR2x2_ASAP7_75t_L g3125 ( 
.A(n_2923),
.B(n_2645),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2932),
.B(n_2578),
.Y(n_3126)
);

HB1xp67_ASAP7_75t_L g3127 ( 
.A(n_2934),
.Y(n_3127)
);

INVx2_ASAP7_75t_SL g3128 ( 
.A(n_2815),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_2925),
.B(n_2645),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_3025),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_3088),
.Y(n_3131)
);

AND2x4_ASAP7_75t_L g3132 ( 
.A(n_3072),
.B(n_2950),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_3025),
.Y(n_3133)
);

OR2x2_ASAP7_75t_L g3134 ( 
.A(n_3001),
.B(n_2929),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3001),
.B(n_2958),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3010),
.Y(n_3136)
);

AND2x4_ASAP7_75t_L g3137 ( 
.A(n_3072),
.B(n_2855),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_3028),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_3047),
.B(n_2873),
.Y(n_3139)
);

NOR3xp33_ASAP7_75t_L g3140 ( 
.A(n_3015),
.B(n_2842),
.C(n_2803),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3010),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3027),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3027),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3043),
.Y(n_3144)
);

OR2x2_ASAP7_75t_L g3145 ( 
.A(n_3043),
.B(n_2979),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_3047),
.B(n_3120),
.Y(n_3146)
);

NOR2xp67_ASAP7_75t_L g3147 ( 
.A(n_3011),
.B(n_2911),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3031),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3031),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3077),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_3120),
.B(n_3124),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_3077),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_3003),
.B(n_2939),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_3124),
.B(n_2876),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_3072),
.B(n_2879),
.Y(n_3155)
);

AND2x6_ASAP7_75t_L g3156 ( 
.A(n_3107),
.B(n_2802),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_3053),
.B(n_2796),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_3021),
.B(n_2959),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3005),
.Y(n_3159)
);

OAI221xp5_ASAP7_75t_SL g3160 ( 
.A1(n_3004),
.A2(n_2975),
.B1(n_2863),
.B2(n_2887),
.C(n_2903),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3006),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3007),
.Y(n_3162)
);

NAND2xp33_ASAP7_75t_SL g3163 ( 
.A(n_3127),
.B(n_2811),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3008),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_3118),
.B(n_2876),
.Y(n_3165)
);

AND2x4_ASAP7_75t_SL g3166 ( 
.A(n_3088),
.B(n_2834),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3012),
.B(n_2872),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_3045),
.Y(n_3168)
);

OAI221xp5_ASAP7_75t_SL g3169 ( 
.A1(n_3004),
.A2(n_2863),
.B1(n_2951),
.B2(n_2827),
.C(n_2795),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_3064),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3117),
.B(n_3094),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3014),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_3049),
.B(n_2876),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3117),
.B(n_2877),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_3070),
.B(n_2926),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3105),
.B(n_2964),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3016),
.Y(n_3177)
);

AND2x4_ASAP7_75t_SL g3178 ( 
.A(n_3127),
.B(n_2834),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3094),
.B(n_2877),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_3101),
.B(n_2898),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_3094),
.B(n_2877),
.Y(n_3181)
);

OAI221xp5_ASAP7_75t_SL g3182 ( 
.A1(n_3095),
.A2(n_2899),
.B1(n_2908),
.B2(n_2930),
.C(n_2884),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_3112),
.B(n_2789),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3024),
.Y(n_3184)
);

AOI221xp5_ASAP7_75t_L g3185 ( 
.A1(n_3095),
.A2(n_2993),
.B1(n_2881),
.B2(n_2819),
.C(n_2828),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_3073),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_3073),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3034),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_3081),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_3049),
.B(n_2858),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_3110),
.B(n_2856),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3035),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3023),
.B(n_2856),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_3157),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_3166),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3136),
.B(n_3141),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3152),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3150),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3142),
.Y(n_3199)
);

INVx1_ASAP7_75t_SL g3200 ( 
.A(n_3131),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3143),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3144),
.Y(n_3202)
);

INVx1_ASAP7_75t_SL g3203 ( 
.A(n_3134),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3159),
.Y(n_3204)
);

OR2x2_ASAP7_75t_L g3205 ( 
.A(n_3135),
.B(n_3146),
.Y(n_3205)
);

AND2x4_ASAP7_75t_SL g3206 ( 
.A(n_3171),
.B(n_3107),
.Y(n_3206)
);

BUFx2_ASAP7_75t_L g3207 ( 
.A(n_3163),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3158),
.B(n_3065),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_L g3209 ( 
.A(n_3167),
.B(n_3082),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3151),
.B(n_3101),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_3151),
.B(n_3101),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3161),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_3166),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3146),
.B(n_3048),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3162),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3163),
.A2(n_3040),
.B(n_2831),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3164),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3139),
.B(n_3048),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3172),
.Y(n_3219)
);

NOR2xp33_ASAP7_75t_L g3220 ( 
.A(n_3190),
.B(n_3065),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3139),
.B(n_3048),
.Y(n_3221)
);

OR2x2_ASAP7_75t_L g3222 ( 
.A(n_3148),
.B(n_3080),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3171),
.B(n_3083),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_3185),
.B(n_3040),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3177),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3154),
.B(n_3058),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_3132),
.B(n_3155),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3130),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3130),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3153),
.B(n_3032),
.Y(n_3230)
);

AND2x4_ASAP7_75t_L g3231 ( 
.A(n_3132),
.B(n_3122),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3184),
.Y(n_3232)
);

NAND3xp33_ASAP7_75t_L g3233 ( 
.A(n_3140),
.B(n_3104),
.C(n_3071),
.Y(n_3233)
);

INVx3_ASAP7_75t_L g3234 ( 
.A(n_3156),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3154),
.B(n_3013),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3149),
.B(n_3018),
.Y(n_3236)
);

NAND2xp33_ASAP7_75t_R g3237 ( 
.A(n_3155),
.B(n_3036),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3133),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3175),
.B(n_3029),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3133),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_3179),
.B(n_3181),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_3156),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3179),
.B(n_3013),
.Y(n_3243)
);

HB1xp67_ASAP7_75t_L g3244 ( 
.A(n_3138),
.Y(n_3244)
);

OR2x2_ASAP7_75t_L g3245 ( 
.A(n_3145),
.B(n_3080),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3181),
.B(n_3132),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3188),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3192),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3138),
.Y(n_3249)
);

NOR2xp67_ASAP7_75t_L g3250 ( 
.A(n_3216),
.B(n_3147),
.Y(n_3250)
);

OR2x2_ASAP7_75t_L g3251 ( 
.A(n_3205),
.B(n_3145),
.Y(n_3251)
);

OAI32xp33_ASAP7_75t_L g3252 ( 
.A1(n_3237),
.A2(n_3176),
.A3(n_3125),
.B1(n_3129),
.B2(n_3100),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3197),
.B(n_3183),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3245),
.Y(n_3254)
);

INVxp67_ASAP7_75t_L g3255 ( 
.A(n_3209),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_3205),
.B(n_3173),
.Y(n_3256)
);

INVx2_ASAP7_75t_SL g3257 ( 
.A(n_3195),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_3244),
.Y(n_3258)
);

OAI32xp33_ASAP7_75t_L g3259 ( 
.A1(n_3237),
.A2(n_2940),
.A3(n_3109),
.B1(n_3107),
.B2(n_2986),
.Y(n_3259)
);

OR2x2_ASAP7_75t_L g3260 ( 
.A(n_3208),
.B(n_3173),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3228),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3196),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_R g3263 ( 
.A(n_3195),
.B(n_3019),
.Y(n_3263)
);

NOR2x1_ASAP7_75t_R g3264 ( 
.A(n_3194),
.B(n_2888),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3228),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3246),
.B(n_3155),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_3234),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3226),
.B(n_3183),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_SL g3269 ( 
.A(n_3207),
.B(n_3182),
.Y(n_3269)
);

OAI22xp5_ASAP7_75t_L g3270 ( 
.A1(n_3224),
.A2(n_3169),
.B1(n_3071),
.B2(n_3019),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3204),
.Y(n_3271)
);

OAI31xp33_ASAP7_75t_L g3272 ( 
.A1(n_3224),
.A2(n_3041),
.A3(n_3160),
.B(n_3056),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3246),
.B(n_3180),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3236),
.B(n_3106),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3212),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3215),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3226),
.B(n_3165),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3217),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3229),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3219),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3241),
.B(n_3180),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_3229),
.Y(n_3282)
);

AOI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_3233),
.A2(n_3175),
.B1(n_3180),
.B2(n_3002),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3238),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3198),
.B(n_3165),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3225),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_3209),
.A2(n_3220),
.B1(n_3200),
.B2(n_3203),
.Y(n_3287)
);

OAI22xp33_ASAP7_75t_SL g3288 ( 
.A1(n_3213),
.A2(n_2878),
.B1(n_3068),
.B2(n_3078),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3235),
.B(n_3174),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3232),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3247),
.Y(n_3291)
);

NAND4xp25_ASAP7_75t_L g3292 ( 
.A(n_3220),
.B(n_2825),
.C(n_3079),
.D(n_3104),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3248),
.Y(n_3293)
);

OAI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_3213),
.A2(n_3193),
.B1(n_3084),
.B2(n_3191),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_3239),
.B(n_2949),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3222),
.Y(n_3296)
);

OAI32xp33_ASAP7_75t_L g3297 ( 
.A1(n_3234),
.A2(n_3109),
.A3(n_2961),
.B1(n_2797),
.B2(n_3061),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3199),
.Y(n_3298)
);

XOR2x2_ASAP7_75t_L g3299 ( 
.A(n_3270),
.B(n_2849),
.Y(n_3299)
);

NOR3xp33_ASAP7_75t_L g3300 ( 
.A(n_3270),
.B(n_3108),
.C(n_3243),
.Y(n_3300)
);

OAI221xp5_ASAP7_75t_L g3301 ( 
.A1(n_3272),
.A2(n_3230),
.B1(n_3079),
.B2(n_3243),
.C(n_3235),
.Y(n_3301)
);

OAI221xp5_ASAP7_75t_L g3302 ( 
.A1(n_3272),
.A2(n_2878),
.B1(n_2954),
.B2(n_2956),
.C(n_2977),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3288),
.A2(n_3054),
.B(n_3234),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3285),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3285),
.Y(n_3305)
);

OAI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_3269),
.A2(n_3250),
.B1(n_3294),
.B2(n_3283),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_3281),
.B(n_3241),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_3258),
.Y(n_3308)
);

AO22x1_ASAP7_75t_L g3309 ( 
.A1(n_3257),
.A2(n_3242),
.B1(n_3156),
.B2(n_2990),
.Y(n_3309)
);

XOR2x2_ASAP7_75t_L g3310 ( 
.A(n_3264),
.B(n_2801),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3256),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3251),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3253),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3261),
.Y(n_3314)
);

INVxp67_ASAP7_75t_SL g3315 ( 
.A(n_3288),
.Y(n_3315)
);

OAI22xp33_ASAP7_75t_L g3316 ( 
.A1(n_3269),
.A2(n_3242),
.B1(n_3109),
.B2(n_3227),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3254),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3260),
.Y(n_3318)
);

XOR2x2_ASAP7_75t_L g3319 ( 
.A(n_3287),
.B(n_2882),
.Y(n_3319)
);

NAND3xp33_ASAP7_75t_L g3320 ( 
.A(n_3292),
.B(n_3202),
.C(n_3201),
.Y(n_3320)
);

AOI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3292),
.A2(n_3227),
.B1(n_3231),
.B2(n_3221),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3294),
.A2(n_3242),
.B1(n_3206),
.B2(n_3227),
.Y(n_3322)
);

OR4x1_ASAP7_75t_L g3323 ( 
.A(n_3252),
.B(n_3128),
.C(n_3249),
.D(n_3087),
.Y(n_3323)
);

AOI22xp33_ASAP7_75t_L g3324 ( 
.A1(n_3255),
.A2(n_3231),
.B1(n_3137),
.B2(n_3221),
.Y(n_3324)
);

OAI31xp33_ASAP7_75t_SL g3325 ( 
.A1(n_3263),
.A2(n_3231),
.A3(n_3214),
.B(n_3210),
.Y(n_3325)
);

BUFx4f_ASAP7_75t_SL g3326 ( 
.A(n_3274),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3271),
.B(n_3238),
.Y(n_3327)
);

A2O1A1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_3259),
.A2(n_3206),
.B(n_3178),
.C(n_3128),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3300),
.A2(n_3267),
.B1(n_3296),
.B2(n_3262),
.Y(n_3329)
);

NOR2xp67_ASAP7_75t_SL g3330 ( 
.A(n_3302),
.B(n_3011),
.Y(n_3330)
);

OAI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3302),
.A2(n_3267),
.B1(n_3268),
.B2(n_3277),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3312),
.Y(n_3332)
);

AOI21xp33_ASAP7_75t_L g3333 ( 
.A1(n_3306),
.A2(n_2875),
.B(n_2957),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3326),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3318),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3327),
.Y(n_3336)
);

NAND2x1p5_ASAP7_75t_L g3337 ( 
.A(n_3303),
.B(n_3011),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3304),
.B(n_3275),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3327),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_3315),
.B(n_3295),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3317),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3314),
.Y(n_3342)
);

OAI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3322),
.A2(n_3321),
.B1(n_3301),
.B2(n_3320),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3325),
.B(n_3266),
.Y(n_3344)
);

O2A1O1Ixp33_ASAP7_75t_L g3345 ( 
.A1(n_3316),
.A2(n_3297),
.B(n_3278),
.C(n_3280),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3311),
.Y(n_3346)
);

OAI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3322),
.A2(n_3289),
.B1(n_3273),
.B2(n_3011),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3325),
.B(n_3214),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3305),
.Y(n_3349)
);

INVxp67_ASAP7_75t_SL g3350 ( 
.A(n_3319),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3313),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3324),
.B(n_3210),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3308),
.Y(n_3353)
);

OAI22xp33_ASAP7_75t_SL g3354 ( 
.A1(n_3323),
.A2(n_3286),
.B1(n_3290),
.B2(n_3276),
.Y(n_3354)
);

AOI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_3299),
.A2(n_3218),
.B1(n_3293),
.B2(n_3291),
.Y(n_3355)
);

INVxp67_ASAP7_75t_L g3356 ( 
.A(n_3310),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3307),
.Y(n_3357)
);

AOI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3309),
.A2(n_3328),
.B1(n_3218),
.B2(n_3211),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_3326),
.B(n_2900),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3312),
.Y(n_3360)
);

AOI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3302),
.A2(n_3211),
.B1(n_3298),
.B2(n_3017),
.Y(n_3361)
);

OAI21xp33_ASAP7_75t_L g3362 ( 
.A1(n_3356),
.A2(n_2820),
.B(n_3121),
.Y(n_3362)
);

NOR3x1_ASAP7_75t_L g3363 ( 
.A(n_3350),
.B(n_2927),
.C(n_2985),
.Y(n_3363)
);

NOR2xp67_ASAP7_75t_L g3364 ( 
.A(n_3343),
.B(n_2791),
.Y(n_3364)
);

OAI211xp5_ASAP7_75t_L g3365 ( 
.A1(n_3333),
.A2(n_2944),
.B(n_2931),
.C(n_2915),
.Y(n_3365)
);

AOI221x1_ASAP7_75t_L g3366 ( 
.A1(n_3333),
.A2(n_2963),
.B1(n_2991),
.B2(n_3038),
.C(n_3062),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_SL g3367 ( 
.A(n_3354),
.B(n_2927),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_3334),
.B(n_3115),
.Y(n_3368)
);

BUFx2_ASAP7_75t_L g3369 ( 
.A(n_3337),
.Y(n_3369)
);

OA22x2_ASAP7_75t_L g3370 ( 
.A1(n_3343),
.A2(n_2899),
.B1(n_3178),
.B2(n_2908),
.Y(n_3370)
);

AND2x2_ASAP7_75t_L g3371 ( 
.A(n_3348),
.B(n_3223),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3338),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3338),
.Y(n_3373)
);

AOI211xp5_ASAP7_75t_SL g3374 ( 
.A1(n_3331),
.A2(n_2963),
.B(n_2945),
.C(n_3087),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_3337),
.B(n_3115),
.Y(n_3375)
);

AOI211xp5_ASAP7_75t_L g3376 ( 
.A1(n_3330),
.A2(n_2919),
.B(n_2867),
.C(n_3061),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3351),
.B(n_3223),
.Y(n_3377)
);

OAI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_3340),
.A2(n_2987),
.B(n_2982),
.Y(n_3378)
);

AOI221xp5_ASAP7_75t_L g3379 ( 
.A1(n_3329),
.A2(n_3039),
.B1(n_3069),
.B2(n_3046),
.C(n_3050),
.Y(n_3379)
);

OR2x2_ASAP7_75t_L g3380 ( 
.A(n_3332),
.B(n_3265),
.Y(n_3380)
);

XNOR2xp5_ASAP7_75t_L g3381 ( 
.A(n_3355),
.B(n_3361),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_3345),
.B(n_3115),
.Y(n_3382)
);

OAI322xp33_ASAP7_75t_L g3383 ( 
.A1(n_3347),
.A2(n_3030),
.A3(n_3063),
.B1(n_3052),
.B2(n_3066),
.C1(n_3051),
.C2(n_3037),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_L g3384 ( 
.A(n_3359),
.B(n_3279),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3335),
.B(n_3284),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3346),
.B(n_3282),
.Y(n_3386)
);

OAI21xp5_ASAP7_75t_SL g3387 ( 
.A1(n_3374),
.A2(n_3344),
.B(n_3358),
.Y(n_3387)
);

OAI211xp5_ASAP7_75t_SL g3388 ( 
.A1(n_3362),
.A2(n_3367),
.B(n_3382),
.C(n_3376),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_SL g3389 ( 
.A1(n_3370),
.A2(n_3369),
.B1(n_3373),
.B2(n_3372),
.Y(n_3389)
);

AOI221x1_ASAP7_75t_SL g3390 ( 
.A1(n_3364),
.A2(n_3360),
.B1(n_3336),
.B2(n_3339),
.C(n_3349),
.Y(n_3390)
);

NOR3xp33_ASAP7_75t_L g3391 ( 
.A(n_3362),
.B(n_3341),
.C(n_3353),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3379),
.B(n_3357),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3377),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3363),
.B(n_3352),
.Y(n_3394)
);

AOI21xp33_ASAP7_75t_L g3395 ( 
.A1(n_3381),
.A2(n_3342),
.B(n_2930),
.Y(n_3395)
);

NAND3xp33_ASAP7_75t_SL g3396 ( 
.A(n_3378),
.B(n_2600),
.C(n_2742),
.Y(n_3396)
);

NOR3xp33_ASAP7_75t_L g3397 ( 
.A(n_3365),
.B(n_2810),
.C(n_2999),
.Y(n_3397)
);

NOR3xp33_ASAP7_75t_L g3398 ( 
.A(n_3375),
.B(n_2326),
.C(n_2320),
.Y(n_3398)
);

AO22x2_ASAP7_75t_L g3399 ( 
.A1(n_3366),
.A2(n_3113),
.B1(n_3092),
.B2(n_3076),
.Y(n_3399)
);

NOR3xp33_ASAP7_75t_L g3400 ( 
.A(n_3383),
.B(n_2326),
.C(n_2320),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3368),
.A2(n_3137),
.B(n_3126),
.Y(n_3401)
);

OAI211xp5_ASAP7_75t_SL g3402 ( 
.A1(n_3384),
.A2(n_3044),
.B(n_3119),
.C(n_3122),
.Y(n_3402)
);

OAI211xp5_ASAP7_75t_SL g3403 ( 
.A1(n_3385),
.A2(n_3122),
.B(n_3033),
.C(n_3090),
.Y(n_3403)
);

NAND3xp33_ASAP7_75t_L g3404 ( 
.A(n_3386),
.B(n_3137),
.C(n_2914),
.Y(n_3404)
);

OA22x2_ASAP7_75t_L g3405 ( 
.A1(n_3368),
.A2(n_2884),
.B1(n_3009),
.B2(n_3026),
.Y(n_3405)
);

NOR3x1_ASAP7_75t_L g3406 ( 
.A(n_3387),
.B(n_3380),
.C(n_2805),
.Y(n_3406)
);

OAI211xp5_ASAP7_75t_SL g3407 ( 
.A1(n_3389),
.A2(n_3102),
.B(n_3074),
.C(n_3093),
.Y(n_3407)
);

AOI221xp5_ASAP7_75t_L g3408 ( 
.A1(n_3390),
.A2(n_3371),
.B1(n_3098),
.B2(n_3038),
.C(n_3067),
.Y(n_3408)
);

NAND2xp33_ASAP7_75t_R g3409 ( 
.A(n_3394),
.B(n_2818),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3399),
.Y(n_3410)
);

O2A1O1Ixp33_ASAP7_75t_L g3411 ( 
.A1(n_3388),
.A2(n_2633),
.B(n_2952),
.C(n_2589),
.Y(n_3411)
);

AOI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3391),
.A2(n_3156),
.B1(n_2910),
.B2(n_2848),
.Y(n_3412)
);

OAI221xp5_ASAP7_75t_L g3413 ( 
.A1(n_3395),
.A2(n_2826),
.B1(n_2854),
.B2(n_2852),
.C(n_2922),
.Y(n_3413)
);

O2A1O1Ixp33_ASAP7_75t_L g3414 ( 
.A1(n_3396),
.A2(n_2616),
.B(n_2570),
.C(n_2996),
.Y(n_3414)
);

AOI221xp5_ASAP7_75t_SL g3415 ( 
.A1(n_3392),
.A2(n_3055),
.B1(n_3057),
.B2(n_3123),
.C(n_3075),
.Y(n_3415)
);

AOI222xp33_ASAP7_75t_L g3416 ( 
.A1(n_3393),
.A2(n_3156),
.B1(n_3240),
.B2(n_3103),
.C1(n_3060),
.C2(n_3099),
.Y(n_3416)
);

AOI211xp5_ASAP7_75t_L g3417 ( 
.A1(n_3400),
.A2(n_2818),
.B(n_2753),
.C(n_2893),
.Y(n_3417)
);

INVx2_ASAP7_75t_SL g3418 ( 
.A(n_3405),
.Y(n_3418)
);

AOI222xp33_ASAP7_75t_L g3419 ( 
.A1(n_3399),
.A2(n_3156),
.B1(n_3240),
.B2(n_3097),
.C1(n_3112),
.C2(n_3009),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3397),
.B(n_3022),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3403),
.Y(n_3421)
);

AOI221xp5_ASAP7_75t_L g3422 ( 
.A1(n_3404),
.A2(n_3091),
.B1(n_3111),
.B2(n_3096),
.C(n_3114),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_3410),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3418),
.A2(n_3402),
.B1(n_3398),
.B2(n_3401),
.Y(n_3424)
);

NOR2x1_ASAP7_75t_L g3425 ( 
.A(n_3407),
.B(n_2251),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3420),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3421),
.Y(n_3427)
);

AOI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3409),
.A2(n_2924),
.B1(n_2918),
.B2(n_2921),
.Y(n_3428)
);

AOI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_3415),
.A2(n_2921),
.B1(n_2844),
.B2(n_2823),
.Y(n_3429)
);

NOR2x1p5_ASAP7_75t_L g3430 ( 
.A(n_3406),
.B(n_2753),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3414),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3411),
.Y(n_3432)
);

NOR2xp33_ASAP7_75t_L g3433 ( 
.A(n_3408),
.B(n_3089),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_3412),
.B(n_3020),
.Y(n_3434)
);

NAND2x1p5_ASAP7_75t_L g3435 ( 
.A(n_3423),
.B(n_2753),
.Y(n_3435)
);

NAND4xp75_ASAP7_75t_L g3436 ( 
.A(n_3427),
.B(n_3422),
.C(n_3417),
.D(n_3419),
.Y(n_3436)
);

NOR3xp33_ASAP7_75t_SL g3437 ( 
.A(n_3432),
.B(n_3413),
.C(n_3416),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3431),
.A2(n_2893),
.B(n_2912),
.Y(n_3438)
);

AOI221xp5_ASAP7_75t_L g3439 ( 
.A1(n_3426),
.A2(n_2912),
.B1(n_2844),
.B2(n_3091),
.C(n_3111),
.Y(n_3439)
);

XNOR2x1_ASAP7_75t_L g3440 ( 
.A(n_3430),
.B(n_3424),
.Y(n_3440)
);

NOR3xp33_ASAP7_75t_L g3441 ( 
.A(n_3433),
.B(n_2285),
.C(n_2280),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3429),
.B(n_3085),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_3434),
.Y(n_3443)
);

HB1xp67_ASAP7_75t_L g3444 ( 
.A(n_3443),
.Y(n_3444)
);

CKINVDCx14_ASAP7_75t_R g3445 ( 
.A(n_3443),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3437),
.B(n_3428),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_3438),
.Y(n_3447)
);

CKINVDCx16_ASAP7_75t_R g3448 ( 
.A(n_3442),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3444),
.Y(n_3449)
);

XNOR2xp5_ASAP7_75t_L g3450 ( 
.A(n_3446),
.B(n_3440),
.Y(n_3450)
);

AO22x1_ASAP7_75t_SL g3451 ( 
.A1(n_3445),
.A2(n_3435),
.B1(n_3436),
.B2(n_3441),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3448),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3447),
.Y(n_3453)
);

AO22x2_ASAP7_75t_L g3454 ( 
.A1(n_3452),
.A2(n_3439),
.B1(n_3425),
.B2(n_3042),
.Y(n_3454)
);

OAI22xp5_ASAP7_75t_L g3455 ( 
.A1(n_3449),
.A2(n_3189),
.B1(n_3187),
.B2(n_3186),
.Y(n_3455)
);

AO22x2_ASAP7_75t_L g3456 ( 
.A1(n_3451),
.A2(n_3042),
.B1(n_3170),
.B2(n_3168),
.Y(n_3456)
);

INVx1_ASAP7_75t_SL g3457 ( 
.A(n_3453),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3457),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3456),
.A2(n_3450),
.B1(n_3453),
.B2(n_3116),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3458),
.A2(n_3454),
.B(n_3455),
.Y(n_3460)
);

AOI22x1_ASAP7_75t_L g3461 ( 
.A1(n_3460),
.A2(n_3459),
.B1(n_2455),
.B2(n_2351),
.Y(n_3461)
);

AOI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_3461),
.A2(n_2275),
.B1(n_2264),
.B2(n_2251),
.Y(n_3462)
);

OR2x6_ASAP7_75t_L g3463 ( 
.A(n_3462),
.B(n_2250),
.Y(n_3463)
);

AOI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3463),
.A2(n_2264),
.B1(n_3059),
.B2(n_3086),
.Y(n_3464)
);


endmodule