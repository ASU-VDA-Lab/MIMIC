module fake_jpeg_683_n_702 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_702);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_702;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_62),
.B(n_89),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_67),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_26),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_73),
.A2(n_51),
.B1(n_45),
.B2(n_32),
.Y(n_199)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_76),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_85),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_80),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_81),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_7),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_86),
.Y(n_206)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_33),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_93),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_104),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_38),
.B(n_10),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_107),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_60),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

CKINVDCx10_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_29),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_13),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_38),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_127),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_119),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_39),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_39),
.B(n_0),
.CON(n_129),
.SN(n_129)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_40),
.Y(n_191)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_42),
.Y(n_132)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

BUFx2_ASAP7_75t_R g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_140),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_144),
.B(n_156),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_79),
.B(n_57),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_147),
.B(n_208),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_31),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_39),
.B1(n_21),
.B2(n_55),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_162),
.A2(n_174),
.B1(n_184),
.B2(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_95),
.B(n_57),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_170),
.B(n_220),
.Y(n_294)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_70),
.A2(n_39),
.B1(n_21),
.B2(n_55),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_58),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_188),
.Y(n_241)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_90),
.A2(n_58),
.B1(n_40),
.B2(n_29),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_116),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_191),
.B(n_129),
.Y(n_250)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_65),
.Y(n_194)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_31),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_219),
.Y(n_251)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_64),
.B(n_51),
.C(n_45),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_75),
.Y(n_210)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_77),
.B(n_32),
.C(n_48),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_212),
.B(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_216),
.Y(n_308)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_78),
.B(n_14),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_84),
.B(n_14),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_121),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_226),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_88),
.B(n_14),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_93),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_213),
.Y(n_231)
);

INVx4_ASAP7_75t_SL g325 ( 
.A(n_231),
.Y(n_325)
);

CKINVDCx12_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

BUFx24_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_237),
.B(n_244),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_94),
.B1(n_103),
.B2(n_120),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_238),
.A2(n_239),
.B1(n_249),
.B2(n_280),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_121),
.B1(n_108),
.B2(n_102),
.Y(n_239)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_245),
.Y(n_343)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_246),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_157),
.A2(n_110),
.B1(n_104),
.B2(n_119),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_248),
.A2(n_177),
.B1(n_214),
.B2(n_203),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_179),
.A2(n_100),
.B1(n_96),
.B2(n_126),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_218),
.Y(n_330)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_190),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_268),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_192),
.B(n_105),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_259),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_16),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_262),
.Y(n_350)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_171),
.Y(n_263)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_263),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_147),
.B(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_267),
.Y(n_320)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_160),
.Y(n_265)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_265),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_164),
.B(n_15),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_157),
.B(n_124),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_164),
.B(n_14),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_273),
.Y(n_322)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_142),
.B(n_151),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_145),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_150),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_278),
.Y(n_332)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_154),
.B(n_19),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_159),
.B(n_12),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_283),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_223),
.A2(n_80),
.B1(n_54),
.B2(n_44),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_137),
.A2(n_48),
.B1(n_122),
.B2(n_54),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_281),
.A2(n_285),
.B1(n_288),
.B2(n_290),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_150),
.B(n_0),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_137),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_301),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_226),
.A2(n_122),
.B1(n_80),
.B2(n_42),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_184),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_163),
.Y(n_289)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_187),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_302),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_162),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_292),
.A2(n_263),
.B1(n_231),
.B2(n_274),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_169),
.A2(n_4),
.B1(n_12),
.B2(n_1),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_296),
.A2(n_298),
.B1(n_312),
.B2(n_155),
.Y(n_361)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_141),
.Y(n_297)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_187),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_207),
.Y(n_336)
);

CKINVDCx12_ASAP7_75t_R g300 ( 
.A(n_207),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_300),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_178),
.B(n_1),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_196),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_135),
.B(n_2),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_305),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_153),
.B(n_136),
.Y(n_305)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_163),
.Y(n_306)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_138),
.B(n_201),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_311),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_196),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_309),
.B(n_266),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_145),
.Y(n_310)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_139),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_213),
.A2(n_185),
.B1(n_152),
.B2(n_205),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_315),
.A2(n_348),
.B1(n_360),
.B2(n_365),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_255),
.A2(n_177),
.B1(n_206),
.B2(n_165),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_323),
.A2(n_355),
.B1(n_362),
.B2(n_373),
.Y(n_408)
);

AO22x2_ASAP7_75t_L g324 ( 
.A1(n_248),
.A2(n_174),
.B1(n_168),
.B2(n_200),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_328),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_268),
.B(n_211),
.CI(n_213),
.CON(n_327),
.SN(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_327),
.A2(n_256),
.B(n_293),
.C(n_269),
.Y(n_420)
);

AO22x1_ASAP7_75t_SL g328 ( 
.A1(n_299),
.A2(n_206),
.B1(n_165),
.B2(n_146),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g329 ( 
.A1(n_238),
.A2(n_181),
.B1(n_172),
.B2(n_211),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_336),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_330),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_347),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_299),
.A2(n_181),
.B1(n_214),
.B2(n_203),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_193),
.C(n_202),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_261),
.C(n_310),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_294),
.B1(n_254),
.B2(n_251),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_175),
.B1(n_221),
.B2(n_186),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_361),
.A2(n_242),
.B1(n_246),
.B2(n_235),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_295),
.A2(n_167),
.B1(n_221),
.B2(n_186),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_233),
.B(n_175),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_364),
.B(n_230),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_241),
.A2(n_167),
.B1(n_148),
.B2(n_134),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_237),
.A2(n_134),
.B1(n_148),
.B2(n_222),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_366),
.A2(n_234),
.B1(n_260),
.B2(n_289),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_264),
.A2(n_283),
.B(n_275),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_367),
.A2(n_285),
.B(n_286),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_266),
.B(n_209),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_368),
.Y(n_409)
);

AO22x1_ASAP7_75t_SL g370 ( 
.A1(n_230),
.A2(n_222),
.B1(n_236),
.B2(n_247),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_276),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_240),
.B(n_243),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_375),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_282),
.B(n_308),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_336),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_252),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_377),
.B(n_407),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_287),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_371),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_253),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_386),
.B(n_391),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_392),
.Y(n_439)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

BUFx4f_ASAP7_75t_SL g466 ( 
.A(n_388),
.Y(n_466)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_326),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_311),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_320),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_393),
.B(n_368),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_321),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_394),
.B(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_341),
.B(n_236),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_403),
.B(n_404),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_322),
.B(n_337),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_405),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_344),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_410),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_321),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_323),
.A2(n_306),
.B1(n_245),
.B2(n_265),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_360),
.B1(n_396),
.B2(n_390),
.Y(n_426)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_417),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_247),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_419),
.Y(n_463)
);

INVx13_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_415),
.Y(n_436)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_416),
.Y(n_440)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

OA22x2_ASAP7_75t_L g451 ( 
.A1(n_418),
.A2(n_358),
.B1(n_297),
.B2(n_318),
.Y(n_451)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_420),
.A2(n_358),
.B(n_314),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_332),
.B(n_262),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_422),
.Y(n_429)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_424),
.Y(n_462)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_425),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_426),
.A2(n_428),
.B1(n_446),
.B2(n_447),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_381),
.A2(n_319),
.B1(n_315),
.B2(n_324),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_381),
.A2(n_345),
.B1(n_335),
.B2(n_366),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_430),
.A2(n_441),
.B1(n_448),
.B2(n_458),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_433),
.A2(n_467),
.B(n_377),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_381),
.A2(n_348),
.B1(n_327),
.B2(n_365),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_398),
.A2(n_336),
.B(n_327),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_461),
.B(n_379),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_397),
.A2(n_324),
.B1(n_362),
.B2(n_328),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_400),
.A2(n_324),
.B1(n_328),
.B2(n_334),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_329),
.B1(n_340),
.B2(n_343),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_385),
.Y(n_449)
);

INVx13_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_451),
.B(n_383),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_382),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_416),
.Y(n_453)
);

INVx13_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_408),
.A2(n_329),
.B1(n_343),
.B2(n_356),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_368),
.B(n_325),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_420),
.A2(n_329),
.B1(n_356),
.B2(n_313),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_465),
.A2(n_458),
.B1(n_448),
.B2(n_461),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_459),
.B1(n_430),
.B2(n_441),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_468),
.A2(n_475),
.B1(n_489),
.B2(n_497),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_443),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_491),
.Y(n_515)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_485),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_474),
.A2(n_487),
.B(n_490),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_455),
.A2(n_396),
.B1(n_401),
.B2(n_400),
.Y(n_475)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_433),
.B(n_434),
.CI(n_392),
.CON(n_477),
.SN(n_477)
);

A2O1A1O1Ixp25_ASAP7_75t_L g511 ( 
.A1(n_477),
.A2(n_439),
.B(n_444),
.C(n_465),
.D(n_463),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_429),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_478),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g512 ( 
.A1(n_479),
.A2(n_467),
.B(n_447),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_399),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_480),
.B(n_494),
.Y(n_509)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_481),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_409),
.Y(n_529)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_484),
.Y(n_526)
);

AOI322xp5_ASAP7_75t_SL g485 ( 
.A1(n_453),
.A2(n_457),
.A3(n_429),
.B1(n_399),
.B2(n_388),
.C1(n_414),
.C2(n_415),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_428),
.A2(n_376),
.B1(n_407),
.B2(n_411),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_486),
.A2(n_488),
.B1(n_467),
.B2(n_446),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_445),
.A2(n_377),
.B(n_379),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_459),
.A2(n_407),
.B1(n_378),
.B2(n_377),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_426),
.A2(n_418),
.B1(n_387),
.B2(n_393),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_435),
.A2(n_406),
.B(n_413),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_435),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_433),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_462),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_440),
.B(n_425),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_466),
.Y(n_496)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_419),
.Y(n_498)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_413),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_434),
.C(n_452),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_466),
.Y(n_500)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_500),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_502),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_405),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_503),
.A2(n_451),
.B(n_462),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_466),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_504),
.B(n_454),
.Y(n_523)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_437),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_409),
.Y(n_517)
);

MAJx2_ASAP7_75t_L g553 ( 
.A(n_510),
.B(n_511),
.C(n_529),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_512),
.A2(n_522),
.B(n_528),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_513),
.A2(n_483),
.B1(n_476),
.B2(n_497),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_436),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_518),
.B(n_520),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_454),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_525),
.Y(n_552)
);

AO22x1_ASAP7_75t_L g525 ( 
.A1(n_468),
.A2(n_451),
.B1(n_460),
.B2(n_442),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_499),
.B(n_450),
.C(n_422),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_491),
.C(n_502),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_493),
.A2(n_460),
.B(n_442),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_531),
.Y(n_549)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_532),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_481),
.B(n_350),
.Y(n_533)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_533),
.B(n_534),
.C(n_538),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_484),
.B(n_350),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_492),
.B(n_456),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_498),
.B(n_437),
.Y(n_539)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_474),
.B(n_451),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_542),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_493),
.B(n_423),
.Y(n_542)
);

AOI21xp33_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_424),
.B(n_389),
.Y(n_543)
);

OAI21xp33_ASAP7_75t_L g559 ( 
.A1(n_543),
.A2(n_488),
.B(n_503),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_476),
.B(n_331),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_490),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_547),
.A2(n_554),
.B1(n_559),
.B2(n_560),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_510),
.B(n_489),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_548),
.B(n_558),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_515),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_561),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_521),
.A2(n_486),
.B1(n_475),
.B2(n_503),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_528),
.A2(n_524),
.B(n_479),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_556),
.A2(n_524),
.B(n_540),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_557),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_521),
.A2(n_495),
.B1(n_470),
.B2(n_471),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_509),
.B(n_507),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_562),
.B(n_563),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_483),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_506),
.C(n_477),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_564),
.B(n_519),
.C(n_544),
.Y(n_581)
);

XNOR2x1_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_477),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g585 ( 
.A(n_565),
.B(n_574),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_515),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_566),
.B(n_567),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_537),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_509),
.B(n_501),
.Y(n_569)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_569),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_570),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_530),
.A2(n_495),
.B1(n_506),
.B2(n_504),
.Y(n_571)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_571),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_535),
.A2(n_505),
.B1(n_500),
.B2(n_496),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_573),
.A2(n_541),
.B1(n_526),
.B2(n_516),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_473),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_537),
.B(n_417),
.Y(n_576)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_576),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_539),
.B(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_577),
.Y(n_604)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_578),
.B(n_532),
.Y(n_586)
);

XNOR2x1_ASAP7_75t_L g615 ( 
.A(n_580),
.B(n_595),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_573),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_547),
.A2(n_512),
.B1(n_511),
.B2(n_525),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_582),
.A2(n_583),
.B1(n_587),
.B2(n_596),
.Y(n_613)
);

OAI22x1_ASAP7_75t_L g583 ( 
.A1(n_552),
.A2(n_522),
.B1(n_525),
.B2(n_512),
.Y(n_583)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_552),
.A2(n_522),
.B1(n_532),
.B2(n_526),
.Y(n_587)
);

AOI211xp5_ASAP7_75t_SL g588 ( 
.A1(n_557),
.A2(n_473),
.B(n_523),
.C(n_536),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_588),
.A2(n_568),
.B(n_577),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_548),
.B(n_564),
.C(n_562),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_589),
.B(n_591),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_553),
.B(n_541),
.C(n_536),
.Y(n_591)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_553),
.B(n_531),
.C(n_516),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_594),
.B(n_597),
.C(n_600),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_565),
.B(n_514),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_546),
.A2(n_514),
.B1(n_508),
.B2(n_412),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_508),
.C(n_363),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_545),
.B(n_363),
.C(n_342),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_545),
.B(n_342),
.C(n_410),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_568),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_607),
.B(n_606),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_608),
.B(n_611),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_583),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_592),
.B(n_555),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_567),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_612),
.B(n_614),
.Y(n_643)
);

FAx1_ASAP7_75t_SL g614 ( 
.A(n_587),
.B(n_546),
.CI(n_557),
.CON(n_614),
.SN(n_614)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_579),
.A2(n_550),
.B1(n_575),
.B2(n_549),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_616),
.A2(n_629),
.B1(n_630),
.B2(n_550),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_598),
.B(n_605),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_617),
.B(n_618),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_556),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_558),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_619),
.B(n_621),
.Y(n_645)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_593),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_625),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_591),
.B(n_574),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_597),
.B(n_578),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_624),
.B(n_600),
.Y(n_649)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_604),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_627),
.B(n_628),
.Y(n_646)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_596),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_602),
.Y(n_630)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_632),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_SL g633 ( 
.A(n_615),
.B(n_582),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_633),
.B(n_634),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_589),
.C(n_581),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_626),
.B(n_594),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_642),
.Y(n_659)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_636),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_618),
.B(n_590),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_637),
.B(n_639),
.Y(n_664)
);

MAJx2_ASAP7_75t_L g638 ( 
.A(n_615),
.B(n_595),
.C(n_585),
.Y(n_638)
);

FAx1_ASAP7_75t_SL g655 ( 
.A(n_638),
.B(n_619),
.CI(n_614),
.CON(n_655),
.SN(n_655)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_585),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_622),
.A2(n_599),
.B1(n_572),
.B2(n_549),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_640),
.B(n_647),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_623),
.B(n_572),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_613),
.A2(n_580),
.B1(n_557),
.B2(n_588),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_648),
.B(n_649),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_346),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_650),
.B(n_359),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_635),
.B(n_607),
.C(n_624),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_653),
.B(n_657),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_655),
.A2(n_666),
.B(n_667),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_634),
.B(n_620),
.C(n_609),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_643),
.A2(n_610),
.B(n_613),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_660),
.A2(n_661),
.B(n_272),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_631),
.A2(n_609),
.B(n_614),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_645),
.B(n_612),
.C(n_627),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_663),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_359),
.C(n_331),
.Y(n_663)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_665),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_636),
.A2(n_256),
.B(n_269),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_644),
.A2(n_271),
.B(n_276),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_637),
.C(n_650),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_669),
.B(n_672),
.Y(n_683)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_662),
.Y(n_670)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_670),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_639),
.C(n_633),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_659),
.B(n_646),
.Y(n_674)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_674),
.Y(n_688)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_638),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_675),
.B(n_679),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_659),
.B(n_293),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_676),
.A2(n_667),
.B(n_656),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_678),
.A2(n_666),
.B(n_654),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_651),
.A2(n_277),
.B1(n_303),
.B2(n_291),
.Y(n_679)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_680),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_671),
.A2(n_658),
.B(n_660),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_681),
.A2(n_684),
.B(n_655),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_682),
.A2(n_675),
.B(n_668),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_677),
.A2(n_661),
.B(n_673),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_669),
.B(n_664),
.C(n_663),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_685),
.B(n_672),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_689),
.B(n_691),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_686),
.A2(n_679),
.B1(n_655),
.B2(n_664),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_692),
.Y(n_696)
);

BUFx24_ASAP7_75t_SL g694 ( 
.A(n_693),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_695),
.A2(n_688),
.B(n_683),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_SL g699 ( 
.A(n_697),
.B(n_698),
.Y(n_699)
);

OAI311xp33_ASAP7_75t_L g698 ( 
.A1(n_694),
.A2(n_682),
.A3(n_690),
.B1(n_687),
.C1(n_685),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_699),
.B(n_696),
.Y(n_700)
);

XOR2xp5_ASAP7_75t_L g701 ( 
.A(n_700),
.B(n_303),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_701),
.B(n_291),
.Y(n_702)
);


endmodule