module real_jpeg_9397_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_13),
.CON(n_12),
.SN(n_12)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_9),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_18),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OA21x2_ASAP7_75t_L g13 ( 
.A1(n_2),
.A2(n_14),
.B(n_15),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_14),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_11),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_9),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_3),
.A2(n_18),
.B(n_24),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_17),
.B(n_25),
.C(n_34),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_8)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B(n_21),
.Y(n_19)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_23),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_30),
.B(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);


endmodule