module fake_netlist_1_10579_n_619 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_619);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_619;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_60), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_50), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_16), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_35), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_33), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_29), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_26), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_0), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_18), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_69), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_19), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_22), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_46), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_68), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_39), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_21), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_18), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_6), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_56), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_30), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_44), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_2), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_0), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_72), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_11), .Y(n_104) );
BUFx2_ASAP7_75t_SL g105 ( .A(n_42), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_32), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_65), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_24), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_63), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_48), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_52), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_34), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_5), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_81), .B(n_1), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_111), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_74), .Y(n_121) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_82), .B(n_31), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_98), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_85), .Y(n_125) );
BUFx8_ASAP7_75t_L g126 ( .A(n_75), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_105), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_78), .B(n_28), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_118), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_110), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_80), .B(n_1), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_109), .Y(n_142) );
NAND2xp33_ASAP7_75t_R g143 ( .A(n_94), .B(n_37), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_89), .B(n_3), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_100), .Y(n_146) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_89), .A2(n_38), .B(n_70), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g148 ( .A(n_76), .B(n_27), .C(n_67), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_90), .B(n_3), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_117), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_76), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_92), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_97), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_87), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_87), .B(n_4), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_159), .B(n_102), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_136), .B(n_102), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_128), .B(n_86), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_128), .B(n_150), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_159), .A2(n_103), .B1(n_93), .B2(n_113), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_131), .B(n_108), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_146), .A2(n_112), .B1(n_115), .B2(n_101), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_144), .B(n_107), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_125), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
AO22x2_ASAP7_75t_L g175 ( .A1(n_159), .A2(n_103), .B1(n_113), .B2(n_105), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_154), .B(n_116), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_126), .B(n_99), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_152), .A2(n_115), .B1(n_95), .B2(n_112), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_119), .B(n_101), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_158), .B(n_95), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_158), .B(n_104), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_131), .B(n_114), .Y(n_191) );
AO22x2_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_96), .B1(n_84), .B2(n_88), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_124), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_119), .B(n_82), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_124), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_135), .B(n_106), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_138), .B(n_4), .Y(n_200) );
INVx5_ASAP7_75t_L g201 ( .A(n_133), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_138), .A2(n_7), .B(n_9), .C(n_10), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_133), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_140), .B(n_12), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_147), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_127), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_127), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_120), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_167), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_196), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_169), .B(n_126), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_190), .B(n_126), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_126), .B1(n_155), .B2(n_143), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_200), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_195), .B(n_140), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_190), .B(n_145), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_178), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_190), .B(n_149), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_195), .Y(n_223) );
INVx6_ASAP7_75t_L g224 ( .A(n_200), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_171), .B(n_157), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_200), .Y(n_226) );
CKINVDCx11_ASAP7_75t_R g227 ( .A(n_173), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_162), .B(n_123), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_173), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_171), .B(n_121), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_182), .B(n_157), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_189), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_191), .B(n_157), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_182), .B(n_153), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_189), .B(n_153), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_165), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_189), .B(n_153), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_210), .B(n_151), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_133), .B1(n_139), .B2(n_137), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_175), .A2(n_133), .B1(n_127), .B2(n_137), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_160), .B(n_151), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_160), .B(n_133), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_185), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_161), .B(n_129), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_172), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_180), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_167), .A2(n_151), .B1(n_137), .B2(n_130), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_166), .B(n_129), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_161), .B(n_129), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_211), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_201), .Y(n_262) );
NOR2xp33_ASAP7_75t_R g263 ( .A(n_164), .B(n_122), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_196), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_175), .A2(n_130), .B1(n_120), .B2(n_129), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_199), .B(n_148), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_183), .Y(n_268) );
BUFx8_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_269), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_224), .B(n_209), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_232), .B(n_257), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_224), .A2(n_196), .B1(n_167), .B2(n_192), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_219), .A2(n_201), .B(n_206), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_226), .A2(n_208), .B(n_205), .C(n_204), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_219), .A2(n_201), .B(n_206), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_232), .B(n_167), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_257), .B(n_196), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_212), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_212), .B(n_192), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_257), .B(n_196), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_227), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_243), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_220), .B(n_179), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_269), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_220), .B(n_203), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_220), .B(n_201), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_223), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_261), .Y(n_298) );
INVx5_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_224), .B(n_192), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_269), .A2(n_192), .B1(n_181), .B2(n_202), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_254), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_265), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_170), .B(n_177), .C(n_163), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
NAND2x1_ASAP7_75t_L g307 ( .A(n_224), .B(n_206), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_229), .B(n_12), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_223), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_218), .A2(n_206), .B1(n_163), .B2(n_184), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_238), .B(n_163), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
O2A1O1Ixp5_ASAP7_75t_SL g315 ( .A1(n_253), .A2(n_207), .B(n_168), .C(n_193), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_223), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_301), .A2(n_225), .B1(n_217), .B2(n_231), .C(n_222), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_290), .B(n_218), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_300), .A2(n_247), .B1(n_228), .B2(n_249), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_295), .B(n_267), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_271), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_285), .A2(n_227), .B1(n_213), .B2(n_215), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_278), .A2(n_234), .B(n_242), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_313), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_216), .B1(n_267), .B2(n_244), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_306), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_285), .A2(n_213), .B1(n_263), .B2(n_264), .Y(n_327) );
NOR2x1_ASAP7_75t_SL g328 ( .A(n_300), .B(n_230), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_313), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_300), .B(n_248), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_283), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_292), .B(n_248), .Y(n_332) );
INVx8_ASAP7_75t_L g333 ( .A(n_283), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_283), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g336 ( .A1(n_275), .A2(n_239), .B(n_236), .C(n_245), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_293), .B(n_246), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
INVx4_ASAP7_75t_SL g341 ( .A(n_270), .Y(n_341) );
AND2x6_ASAP7_75t_L g342 ( .A(n_280), .B(n_246), .Y(n_342) );
OAI21xp33_ASAP7_75t_SL g343 ( .A1(n_271), .A2(n_241), .B(n_246), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_274), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_309), .A2(n_267), .B1(n_163), .B2(n_184), .Y(n_345) );
NAND3xp33_ASAP7_75t_SL g346 ( .A(n_309), .B(n_207), .C(n_174), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_330), .A2(n_295), .B1(n_292), .B2(n_280), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_293), .B1(n_270), .B2(n_273), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_330), .B(n_274), .Y(n_350) );
OAI211xp5_ASAP7_75t_L g351 ( .A1(n_319), .A2(n_304), .B(n_284), .C(n_281), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_332), .B(n_295), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_320), .B(n_298), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_333), .A2(n_298), .B1(n_282), .B2(n_287), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_344), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_317), .A2(n_292), .B1(n_296), .B2(n_294), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_340), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_320), .B(n_287), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_333), .B(n_288), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_323), .A2(n_315), .B(n_307), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_332), .B(n_288), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_325), .A2(n_282), .B1(n_276), .B2(n_312), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_333), .B(n_272), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g366 ( .A1(n_336), .A2(n_307), .B(n_272), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_317), .A2(n_286), .B1(n_291), .B2(n_302), .C(n_314), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_322), .A2(n_314), .B(n_168), .C(n_174), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_329), .B(n_296), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_318), .B1(n_334), .B2(n_331), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_345), .A2(n_299), .B1(n_289), .B2(n_297), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_368), .B(n_335), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_347), .B(n_340), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_363), .B(n_342), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_350), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_350), .B(n_328), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_369), .A2(n_327), .B(n_343), .C(n_323), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_363), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
AOI32xp33_ASAP7_75t_L g381 ( .A1(n_349), .A2(n_318), .A3(n_326), .B1(n_296), .B2(n_16), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_364), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_367), .A2(n_356), .B1(n_364), .B2(n_352), .C(n_348), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_365), .Y(n_386) );
INVx4_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_359), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_368), .B(n_346), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_357), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
AO21x2_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_279), .B(n_277), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_351), .B(n_326), .C(n_186), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_315), .B(n_310), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_355), .Y(n_396) );
OAI31xp33_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_306), .A3(n_310), .B(n_341), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
NOR2xp33_ASAP7_75t_R g399 ( .A(n_357), .B(n_342), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g401 ( .A1(n_353), .A2(n_370), .B1(n_358), .B2(n_361), .C1(n_342), .C2(n_341), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_358), .B(n_342), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_357), .Y(n_403) );
NAND2xp33_ASAP7_75t_R g404 ( .A(n_365), .B(n_147), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_390), .B(n_353), .Y(n_406) );
OAI31xp33_ASAP7_75t_L g407 ( .A1(n_397), .A2(n_371), .A3(n_372), .B(n_362), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_390), .B(n_370), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_400), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_400), .B(n_362), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g411 ( .A1(n_381), .A2(n_372), .B(n_366), .Y(n_411) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_387), .B(n_365), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_395), .A2(n_310), .B(n_311), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_381), .A2(n_366), .B(n_341), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_398), .B(n_365), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_385), .B(n_187), .C(n_193), .D(n_186), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_365), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_383), .B(n_337), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_401), .A2(n_337), .B1(n_316), .B2(n_289), .Y(n_423) );
AO21x2_ASAP7_75t_L g424 ( .A1(n_395), .A2(n_187), .B(n_311), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_396), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_387), .B(n_53), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_376), .B(n_13), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_396), .B(n_13), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_382), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_380), .B(n_14), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_388), .B(n_15), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_384), .B(n_374), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_397), .B(n_299), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_384), .B(n_17), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_373), .B(n_17), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_391), .B(n_20), .Y(n_441) );
INVx4_ASAP7_75t_R g442 ( .A(n_391), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_377), .B(n_20), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_402), .B(n_163), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_402), .B(n_206), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_386), .B(n_299), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_184), .Y(n_447) );
OAI33xp33_ASAP7_75t_L g448 ( .A1(n_375), .A2(n_197), .A3(n_188), .B1(n_183), .B2(n_241), .B3(n_252), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_382), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_425), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_425), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_410), .B(n_413), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_406), .B(n_377), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_415), .A2(n_399), .B(n_378), .C(n_403), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_439), .B(n_382), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_434), .A2(n_197), .A3(n_188), .B1(n_404), .B2(n_394), .B3(n_393), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_443), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_412), .A2(n_382), .B1(n_393), .B2(n_299), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_406), .B(n_393), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_408), .B(n_184), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_410), .B(n_184), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_407), .B(n_305), .C(n_308), .D(n_214), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_413), .B(n_23), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_409), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_439), .B(n_25), .Y(n_466) );
NOR2xp33_ASAP7_75t_R g467 ( .A(n_412), .B(n_40), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_426), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_441), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_440), .B(n_41), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_417), .B(n_43), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_45), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_418), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_408), .B(n_316), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_47), .Y(n_479) );
NAND2xp33_ASAP7_75t_SL g480 ( .A(n_405), .B(n_316), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_51), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_443), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_415), .B(n_308), .Y(n_483) );
OAI33xp33_ASAP7_75t_L g484 ( .A1(n_433), .A2(n_54), .A3(n_55), .B1(n_57), .B2(n_58), .B3(n_62), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
AND2x2_ASAP7_75t_SL g487 ( .A(n_412), .B(n_316), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_429), .B(n_316), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_435), .B(n_64), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_429), .B(n_297), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_438), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_438), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_431), .B(n_66), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_435), .B(n_297), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_411), .B(n_289), .C(n_297), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_407), .B(n_305), .C(n_214), .D(n_268), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_422), .B(n_297), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_420), .B(n_289), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_414), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_489), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_469), .B(n_421), .Y(n_503) );
NAND2x1_ASAP7_75t_L g504 ( .A(n_468), .B(n_442), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_455), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g507 ( .A1(n_454), .A2(n_437), .B(n_427), .Y(n_507) );
NOR2xp33_ASAP7_75t_SL g508 ( .A(n_468), .B(n_405), .Y(n_508) );
INVxp33_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_480), .A2(n_411), .B(n_436), .Y(n_510) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_480), .A2(n_426), .B(n_446), .C(n_449), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_484), .B(n_419), .C(n_427), .Y(n_512) );
AOI222xp33_ASAP7_75t_L g513 ( .A1(n_491), .A2(n_423), .B1(n_416), .B2(n_426), .C1(n_448), .C2(n_447), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_471), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_450), .B(n_449), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_486), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_497), .A2(n_437), .A3(n_426), .B(n_419), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_468), .B(n_449), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_494), .Y(n_522) );
OAI21xp33_ASAP7_75t_L g523 ( .A1(n_483), .A2(n_447), .B(n_445), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_492), .A2(n_444), .B1(n_449), .B2(n_432), .C(n_424), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_452), .B(n_432), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_482), .A2(n_432), .B1(n_442), .B2(n_289), .C(n_424), .Y(n_527) );
OAI322xp33_ASAP7_75t_L g528 ( .A1(n_458), .A2(n_460), .A3(n_456), .B1(n_453), .B2(n_466), .C1(n_470), .C2(n_495), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_487), .A2(n_252), .B1(n_268), .B2(n_237), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_452), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_457), .A2(n_251), .B1(n_250), .B2(n_240), .C(n_71), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_459), .B(n_240), .C(n_250), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_489), .Y(n_535) );
O2A1O1Ixp5_ASAP7_75t_L g536 ( .A1(n_495), .A2(n_251), .B(n_230), .C(n_259), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_466), .A2(n_470), .B1(n_496), .B2(n_499), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_476), .B(n_256), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_476), .Y(n_539) );
AOI21xp33_ASAP7_75t_SL g540 ( .A1(n_464), .A2(n_230), .B(n_256), .Y(n_540) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_493), .A2(n_230), .B(n_259), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_465), .B(n_258), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g543 ( .A1(n_464), .A2(n_258), .B1(n_262), .B2(n_472), .C1(n_474), .C2(n_477), .Y(n_543) );
NOR4xp25_ASAP7_75t_L g544 ( .A(n_472), .B(n_262), .C(n_474), .D(n_500), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_479), .A2(n_262), .B(n_481), .C(n_488), .Y(n_545) );
NOR4xp25_ASAP7_75t_SL g546 ( .A(n_527), .B(n_479), .C(n_481), .D(n_490), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_473), .Y(n_547) );
NOR3xp33_ASAP7_75t_SL g548 ( .A(n_510), .B(n_463), .C(n_461), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_524), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
INVxp33_ASAP7_75t_L g551 ( .A(n_508), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_539), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_521), .B(n_462), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_515), .B(n_493), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_511), .A2(n_501), .B(n_498), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_522), .B(n_462), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_506), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_516), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_526), .B(n_501), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_533), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_534), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_503), .B(n_502), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_535), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_537), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_518), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_509), .B(n_507), .Y(n_572) );
NOR3xp33_ASAP7_75t_SL g573 ( .A(n_510), .B(n_517), .C(n_523), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_525), .B(n_544), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_538), .Y(n_575) );
AND3x2_ASAP7_75t_L g576 ( .A(n_574), .B(n_512), .C(n_531), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_549), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_569), .A2(n_512), .B1(n_525), .B2(n_511), .C(n_531), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_570), .B(n_574), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_559), .Y(n_580) );
XNOR2x2_ASAP7_75t_L g581 ( .A(n_572), .B(n_532), .Y(n_581) );
AOI211x1_ASAP7_75t_L g582 ( .A1(n_557), .A2(n_513), .B(n_542), .C(n_543), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_568), .B(n_529), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_552), .B(n_545), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_551), .B(n_536), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
XOR2xp5_ASAP7_75t_L g587 ( .A(n_551), .B(n_541), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_575), .A2(n_541), .B1(n_536), .B2(n_540), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_565), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_561), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_563), .Y(n_591) );
XNOR2xp5_ASAP7_75t_L g592 ( .A(n_573), .B(n_567), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_592), .A2(n_571), .B1(n_562), .B2(n_548), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_579), .A2(n_555), .B1(n_562), .B2(n_547), .C(n_558), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_585), .B(n_550), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_587), .A2(n_550), .B1(n_567), .B2(n_546), .Y(n_596) );
NOR2xp33_ASAP7_75t_R g597 ( .A(n_576), .B(n_550), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g598 ( .A(n_583), .Y(n_598) );
XOR2xp5_ASAP7_75t_L g599 ( .A(n_581), .B(n_553), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_578), .A2(n_555), .B1(n_564), .B2(n_556), .Y(n_600) );
XNOR2x1_ASAP7_75t_L g601 ( .A(n_576), .B(n_556), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_577), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_585), .A2(n_588), .B(n_584), .Y(n_603) );
XNOR2x1_ASAP7_75t_L g604 ( .A(n_582), .B(n_566), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_588), .B(n_554), .C(n_580), .D(n_586), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_591), .B(n_554), .Y(n_606) );
OAI322xp33_ASAP7_75t_L g607 ( .A1(n_589), .A2(n_590), .A3(n_579), .B1(n_592), .B2(n_569), .C1(n_581), .C2(n_572), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_607), .B(n_598), .C(n_603), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_593), .A2(n_600), .B1(n_595), .B2(n_604), .C(n_599), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_602), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_597), .B(n_596), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_611), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_608), .A2(n_601), .B1(n_600), .B2(n_605), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_610), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_614), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_612), .Y(n_616) );
BUFx2_ASAP7_75t_L g617 ( .A(n_616), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_617), .A2(n_609), .B1(n_613), .B2(n_615), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_618), .A2(n_594), .B(n_606), .Y(n_619) );
endmodule