module real_jpeg_26773_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_6),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_8),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_18),
.B(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_67),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_37),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_8),
.B(n_17),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_87),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_86),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_58),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_58),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_31),
.C(n_45),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_14),
.A2(n_15),
.B1(n_31),
.B2(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B(n_25),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_16),
.A2(n_21),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_18),
.A2(n_20),
.B1(n_39),
.B2(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_18),
.A2(n_27),
.B(n_39),
.C(n_92),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_23),
.B(n_27),
.C(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_22),
.A2(n_23),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_27),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_27),
.B(n_35),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_31),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_31),
.A2(n_91),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B(n_40),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_33),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_36),
.B(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_45),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_57),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_54),
.B1(n_74),
.B2(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_80),
.B2(n_81),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_76),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_85),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_96),
.C(n_98),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_114),
.B(n_118),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_100),
.B(n_113),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_110),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_112),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_111),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);


endmodule