module fake_jpeg_29284_n_151 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_151);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_28),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_22),
.C(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_26),
.B1(n_15),
.B2(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_80),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_83),
.Y(n_94)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_87),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_79),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_57),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_81),
.C(n_88),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_41),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_17),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_47),
.B1(n_50),
.B2(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_102),
.B1(n_105),
.B2(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_11),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_16),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_87),
.B1(n_86),
.B2(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_110),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_86),
.B(n_105),
.Y(n_108)
);

XNOR2x1_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_81),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_94),
.B1(n_105),
.B2(n_75),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_82),
.C(n_75),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_116),
.C(n_117),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_8),
.B(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_59),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

NOR4xp25_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_115),
.C(n_92),
.D(n_109),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_124),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_101),
.A3(n_102),
.B1(n_96),
.B2(n_71),
.C1(n_94),
.C2(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_90),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_112),
.B1(n_110),
.B2(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_131),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_114),
.B1(n_90),
.B2(n_50),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_133),
.B(n_123),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_124),
.A3(n_123),
.B1(n_73),
.B2(n_64),
.C1(n_71),
.C2(n_1),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_134),
.B1(n_128),
.B2(n_60),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_138),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_62),
.C(n_56),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_142),
.C(n_73),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_134),
.B(n_2),
.C(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_1),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_2),
.B(n_4),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_135),
.B(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_147),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_73),
.Y(n_151)
);


endmodule