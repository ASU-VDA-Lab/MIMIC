module fake_jpeg_19471_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_19),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_31),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_20),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_16),
.CON(n_48),
.SN(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_31),
.B1(n_23),
.B2(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_18),
.C(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_60),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_65),
.Y(n_94)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_51),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_18),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_71),
.C(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_24),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_79),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_24),
.B1(n_29),
.B2(n_18),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_29),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.C(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_0),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_90),
.B1(n_93),
.B2(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_51),
.B1(n_52),
.B2(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_95),
.B1(n_74),
.B2(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_68),
.B1(n_58),
.B2(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_51),
.B1(n_52),
.B2(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_87),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_73),
.B1(n_71),
.B2(n_9),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_114),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_85),
.B(n_84),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_65),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_121),
.A3(n_125),
.B1(n_94),
.B2(n_102),
.C1(n_100),
.C2(n_8),
.Y(n_133)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_76),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.C(n_74),
.D(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_6),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_6),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_109),
.Y(n_152)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_91),
.B(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_138),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_87),
.B(n_86),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_86),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_142),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_103),
.C2(n_9),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_121),
.B(n_106),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_126),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_108),
.C(n_109),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_141),
.C(n_131),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_123),
.B1(n_112),
.B2(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_144),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_132),
.A3(n_141),
.B1(n_128),
.B2(n_144),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_171),
.C(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_136),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_143),
.C(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_173),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_165),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_151),
.B(n_135),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_151),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_157),
.C(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_165),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_187),
.C(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_130),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_163),
.C(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_135),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_196),
.B(n_181),
.Y(n_197)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_195),
.B(n_164),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_196),
.B(n_125),
.C(n_150),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_11),
.B(n_14),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_160),
.Y(n_203)
);


endmodule