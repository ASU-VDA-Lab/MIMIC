module fake_jpeg_6961_n_208 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_19),
.Y(n_49)
);

CKINVDCx9p33_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_25),
.B1(n_23),
.B2(n_18),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_36),
.B1(n_23),
.B2(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_24),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_23),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_26),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_63),
.B1(n_38),
.B2(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_61),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_52),
.C(n_47),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_49),
.C(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_15),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_47),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_33),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_58),
.Y(n_92)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_81),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_65),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_33),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_22),
.B(n_24),
.Y(n_110)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_57),
.C(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_70),
.B(n_64),
.Y(n_97)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_57),
.B(n_40),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_42),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_72),
.B(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_56),
.B1(n_38),
.B2(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_38),
.B1(n_75),
.B2(n_87),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_94),
.B1(n_92),
.B2(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_126),
.B1(n_131),
.B2(n_106),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_91),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_128),
.B(n_129),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_104),
.A3(n_96),
.B1(n_78),
.B2(n_102),
.C(n_79),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_17),
.B(n_18),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_82),
.B1(n_78),
.B2(n_79),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_110),
.B(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_27),
.B1(n_17),
.B2(n_16),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_93),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_86),
.C(n_107),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_142),
.B1(n_128),
.B2(n_123),
.C(n_16),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_99),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_100),
.C(n_97),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_109),
.B(n_105),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_143),
.B(n_19),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_126),
.C(n_119),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_74),
.C(n_39),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_129),
.C(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_136),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_29),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_107),
.B1(n_108),
.B2(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_162),
.C(n_134),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_13),
.B(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_86),
.Y(n_156)
);

OAI322xp33_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_160),
.A3(n_139),
.B1(n_41),
.B2(n_13),
.C1(n_32),
.C2(n_60),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_67),
.B1(n_41),
.B2(n_37),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_161),
.B(n_143),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_12),
.B(n_2),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_46),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_32),
.C(n_29),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_32),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_141),
.B1(n_139),
.B2(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_60),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_61),
.C(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_163),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_1),
.B(n_3),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_151),
.B1(n_161),
.B2(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_181),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_180),
.B(n_182),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_158),
.B1(n_162),
.B2(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_175),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_165),
.A3(n_172),
.B1(n_150),
.B2(n_171),
.C1(n_167),
.C2(n_9),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_5),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_183),
.C(n_181),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_190),
.B(n_192),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_1),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_183),
.Y(n_195)
);

NOR4xp25_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_190),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_194),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_197),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_11),
.B(n_12),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_8),
.B(n_10),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_10),
.B(n_11),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_205),
.B(n_200),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.Y(n_208)
);


endmodule