module fake_aes_1786_n_625 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_625);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_625;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_504;
wire n_170;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_21), .Y(n_76) );
INVxp33_ASAP7_75t_L g77 ( .A(n_28), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_13), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_32), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_25), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_71), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_72), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_67), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_22), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_60), .Y(n_88) );
BUFx2_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_3), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_7), .B(n_73), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_30), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_66), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_23), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_50), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_18), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_65), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_47), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_58), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_75), .Y(n_104) );
BUFx10_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_2), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_61), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_34), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_68), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_16), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_52), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_15), .Y(n_116) );
BUFx5_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_20), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_48), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_56), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_17), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_89), .B(n_0), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_117), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_113), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_89), .B(n_1), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_80), .B(n_2), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_117), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_117), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_117), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_117), .Y(n_134) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_76), .A2(n_36), .B(n_64), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_117), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_117), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_76), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_82), .B(n_35), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_99), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_101), .B(n_3), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
OR2x2_ASAP7_75t_L g145 ( .A(n_80), .B(n_4), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_77), .B(n_4), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_122), .Y(n_147) );
INVx2_ASAP7_75t_SL g148 ( .A(n_105), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_101), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_120), .B(n_5), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
OR2x6_ASAP7_75t_L g155 ( .A(n_84), .B(n_5), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_88), .A2(n_39), .B(n_62), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
NAND2xp33_ASAP7_75t_L g161 ( .A(n_85), .B(n_37), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_94), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_96), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_124), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_155), .A2(n_102), .B1(n_84), .B2(n_93), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_131), .B(n_100), .Y(n_173) );
OR2x2_ASAP7_75t_SL g174 ( .A(n_126), .B(n_103), .Y(n_174) );
INVx4_ASAP7_75t_SL g175 ( .A(n_139), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_128), .B(n_103), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_131), .B(n_108), .Y(n_177) );
INVx6_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_128), .B(n_102), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_128), .B(n_104), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_142), .B(n_105), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_125), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_148), .B(n_111), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_125), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_146), .B(n_105), .Y(n_192) );
INVx8_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_128), .B(n_104), .Y(n_198) );
INVx4_ASAP7_75t_SL g199 ( .A(n_139), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_133), .Y(n_201) );
INVx6_ASAP7_75t_L g202 ( .A(n_132), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_154), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_148), .B(n_98), .Y(n_206) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_143), .A2(n_97), .B(n_121), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_138), .B(n_98), .Y(n_208) );
INVx3_ASAP7_75t_R g209 ( .A(n_145), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_147), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_138), .B(n_118), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_141), .B(n_116), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_154), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_141), .B(n_107), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_146), .Y(n_218) );
INVx6_ASAP7_75t_L g219 ( .A(n_132), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
INVx6_ASAP7_75t_L g221 ( .A(n_139), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_203), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_203), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_220), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_166), .A2(n_155), .B1(n_123), .B2(n_127), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_192), .B(n_144), .Y(n_228) );
OR2x6_ASAP7_75t_L g229 ( .A(n_193), .B(n_155), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
BUFx12f_ASAP7_75t_L g231 ( .A(n_174), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_220), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_177), .B(n_144), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_193), .A2(n_163), .B1(n_162), .B2(n_152), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_193), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_194), .B(n_87), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_218), .B(n_145), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_192), .B(n_152), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_206), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_218), .B(n_156), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_181), .A2(n_163), .B1(n_162), .B2(n_160), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_206), .B(n_156), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx5_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_186), .B(n_160), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_206), .B(n_157), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_213), .B(n_217), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_181), .A2(n_157), .B1(n_161), .B2(n_78), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_194), .B(n_93), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
AOI21xp33_ASAP7_75t_L g257 ( .A1(n_173), .A2(n_153), .B(n_92), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
INVx5_ASAP7_75t_L g259 ( .A(n_181), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_174), .B(n_90), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_173), .B(n_115), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_208), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_176), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_187), .B(n_79), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_181), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_208), .B(n_83), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_208), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_176), .B(n_115), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_208), .B(n_95), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_176), .B(n_116), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_214), .B(n_149), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_198), .A2(n_139), .B1(n_122), .B2(n_149), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_214), .B(n_154), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_187), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_214), .A2(n_112), .B(n_96), .C(n_97), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_182), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_214), .B(n_139), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
NOR2x1_ASAP7_75t_L g283 ( .A(n_182), .B(n_109), .Y(n_283) );
BUFx12f_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_229), .A2(n_179), .B1(n_140), .B2(n_221), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_231), .B(n_179), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_234), .B(n_198), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_230), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_280), .B(n_209), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_230), .B(n_175), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_229), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_239), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_230), .B(n_179), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_229), .A2(n_179), .B1(n_221), .B2(n_198), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_222), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g300 ( .A1(n_229), .A2(n_207), .B(n_164), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_255), .A2(n_198), .B1(n_207), .B2(n_167), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_230), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_225), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_239), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_225), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_281), .A2(n_172), .B(n_171), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_224), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_224), .B(n_207), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_255), .A2(n_198), .B1(n_172), .B2(n_164), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_255), .A2(n_198), .B1(n_167), .B2(n_169), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_236), .Y(n_316) );
INVx3_ASAP7_75t_SL g317 ( .A(n_266), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_241), .A2(n_185), .B(n_189), .C(n_212), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_242), .B(n_198), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_236), .A2(n_171), .B1(n_169), .B2(n_168), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_257), .B(n_168), .Y(n_322) );
INVx5_ASAP7_75t_L g323 ( .A(n_248), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_242), .B(n_185), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_242), .B(n_175), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_252), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
CKINVDCx11_ASAP7_75t_R g330 ( .A(n_239), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_269), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_312), .A2(n_251), .B1(n_244), .B2(n_235), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_305), .B(n_228), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_313), .A2(n_244), .B1(n_251), .B2(n_270), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_330), .A2(n_283), .B1(n_260), .B2(n_275), .Y(n_337) );
O2A1O1Ixp5_ASAP7_75t_L g338 ( .A1(n_300), .A2(n_265), .B(n_276), .C(n_270), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_290), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_253), .B(n_243), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_287), .A2(n_240), .B(n_249), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_309), .B(n_248), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_295), .B(n_244), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_290), .B(n_248), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_290), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_320), .A2(n_251), .B1(n_270), .B2(n_272), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_284), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_311), .A2(n_260), .B1(n_275), .B2(n_261), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_297), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_275), .B1(n_261), .B2(n_272), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_272), .B1(n_227), .B2(n_245), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_290), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_285), .A2(n_250), .B1(n_237), .B2(n_256), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_322), .A2(n_254), .B1(n_267), .B2(n_271), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_291), .A2(n_279), .B1(n_273), .B2(n_232), .C(n_247), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_307), .A2(n_232), .B1(n_246), .B2(n_247), .C(n_258), .Y(n_362) );
OAI22x1_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_293), .B1(n_316), .B2(n_309), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g364 ( .A1(n_337), .A2(n_301), .B1(n_114), .B2(n_121), .C(n_274), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_356), .B(n_316), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_351), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_352), .A2(n_319), .B1(n_293), .B2(n_298), .C(n_310), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_354), .A2(n_284), .B1(n_321), .B2(n_326), .C1(n_310), .C2(n_297), .Y(n_368) );
AO222x2_ASAP7_75t_L g369 ( .A1(n_351), .A2(n_6), .B1(n_7), .B2(n_8), .C1(n_10), .C2(n_11), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_355), .A2(n_296), .B1(n_299), .B2(n_304), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_318), .B(n_306), .C(n_304), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_333), .B(n_321), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_350), .A2(n_299), .B1(n_306), .B2(n_296), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_339), .A2(n_292), .B(n_314), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_332), .A2(n_297), .B1(n_317), .B2(n_328), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_353), .B(n_258), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g378 ( .A(n_356), .Y(n_378) );
AO221x1_ASAP7_75t_L g379 ( .A1(n_339), .A2(n_303), .B1(n_290), .B2(n_114), .C(n_331), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_326), .B1(n_246), .B2(n_258), .C(n_289), .Y(n_380) );
INVxp33_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_359), .A2(n_303), .B1(n_289), .B2(n_91), .Y(n_382) );
OAI22xp5_ASAP7_75t_SL g383 ( .A1(n_357), .A2(n_317), .B1(n_303), .B2(n_328), .Y(n_383) );
INVx3_ASAP7_75t_SL g384 ( .A(n_348), .Y(n_384) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_345), .A2(n_110), .A3(n_150), .B1(n_147), .B2(n_159), .C1(n_151), .C2(n_189), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_335), .A2(n_327), .B1(n_317), .B2(n_315), .C(n_314), .Y(n_386) );
INVx8_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_336), .A2(n_327), .B1(n_303), .B2(n_259), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_344), .B(n_303), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_378), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_343), .B1(n_361), .B2(n_358), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_369), .A2(n_343), .B1(n_361), .B2(n_358), .C(n_349), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_389), .B(n_347), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_387), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_374), .B(n_347), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_365), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_349), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_364), .A2(n_344), .B1(n_341), .B2(n_362), .C(n_338), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_365), .B(n_339), .Y(n_402) );
AOI33xp33_ASAP7_75t_L g403 ( .A1(n_382), .A2(n_6), .A3(n_8), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_366), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_371), .B(n_348), .Y(n_405) );
OAI211xp5_ASAP7_75t_SL g406 ( .A1(n_368), .A2(n_188), .B(n_191), .C(n_197), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_381), .B(n_135), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_381), .B(n_371), .Y(n_411) );
OR2x6_ASAP7_75t_L g412 ( .A(n_376), .B(n_346), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_367), .A2(n_342), .B1(n_139), .B2(n_325), .C1(n_17), .C2(n_20), .Y(n_413) );
OAI22xp5_ASAP7_75t_SL g414 ( .A1(n_363), .A2(n_342), .B1(n_346), .B2(n_135), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_159), .B1(n_151), .B2(n_150), .C(n_147), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_383), .A2(n_139), .B1(n_325), .B2(n_315), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_346), .B(n_158), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_387), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_314), .B1(n_315), .B2(n_331), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g421 ( .A(n_380), .B(n_14), .C(n_15), .D(n_16), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_158), .B(n_135), .C(n_159), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_384), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_416), .B(n_372), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
OAI33xp33_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_14), .A3(n_188), .B1(n_204), .B2(n_191), .B3(n_197), .Y(n_427) );
OAI31xp33_ASAP7_75t_L g428 ( .A1(n_421), .A2(n_372), .A3(n_329), .B(n_204), .Y(n_428) );
NOR3xp33_ASAP7_75t_SL g429 ( .A(n_392), .B(n_385), .C(n_212), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_392), .B(n_159), .C(n_150), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_421), .A2(n_151), .B(n_150), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g433 ( .A1(n_404), .A2(n_150), .A3(n_151), .B1(n_159), .B2(n_135), .C1(n_158), .C2(n_329), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_413), .A2(n_158), .B1(n_331), .B2(n_329), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_393), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_410), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_390), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_403), .B(n_226), .C(n_233), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_422), .A2(n_282), .B(n_278), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_413), .A2(n_150), .B1(n_159), .B2(n_151), .C(n_178), .Y(n_440) );
OAI33xp33_ASAP7_75t_L g441 ( .A1(n_414), .A2(n_151), .A3(n_233), .B1(n_226), .B2(n_216), .B3(n_165), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_396), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_423), .Y(n_443) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_418), .A2(n_238), .B(n_282), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_416), .B(n_24), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g446 ( .A1(n_390), .A2(n_278), .B1(n_238), .B2(n_262), .C(n_201), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_423), .B(n_407), .C(n_395), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_396), .B(n_27), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g449 ( .A(n_390), .B(n_31), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_411), .A2(n_331), .B1(n_178), .B2(n_219), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_411), .A2(n_331), .B1(n_178), .B2(n_219), .Y(n_451) );
AOI21xp33_ASAP7_75t_SL g452 ( .A1(n_419), .A2(n_33), .B(n_40), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_397), .A2(n_323), .B1(n_248), .B2(n_259), .Y(n_453) );
OAI21x1_ASAP7_75t_L g454 ( .A1(n_418), .A2(n_262), .B(n_196), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_393), .B(n_41), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_399), .B(n_42), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_395), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_397), .B(n_43), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_399), .B(n_44), .Y(n_461) );
OAI321xp33_ASAP7_75t_L g462 ( .A1(n_414), .A2(n_183), .A3(n_205), .B1(n_211), .B2(n_210), .C(n_216), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_399), .B(n_45), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
OAI31xp33_ASAP7_75t_SL g465 ( .A1(n_395), .A2(n_46), .A3(n_49), .B(n_51), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_397), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_398), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_442), .B(n_455), .Y(n_469) );
AO21x1_ASAP7_75t_L g470 ( .A1(n_459), .A2(n_398), .B(n_400), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_447), .B(n_409), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_437), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_426), .B(n_408), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_465), .A2(n_417), .B(n_401), .C(n_415), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_430), .A2(n_406), .B(n_422), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_426), .B(n_408), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_436), .B(n_405), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_443), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_448), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_468), .B(n_402), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_467), .B(n_401), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_424), .B(n_412), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_444), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_457), .B(n_412), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_445), .B(n_412), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_428), .B(n_412), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_449), .B(n_406), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_463), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_458), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_461), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_431), .B(n_409), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g499 ( .A1(n_440), .A2(n_409), .B(n_415), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_461), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_464), .B(n_409), .Y(n_502) );
NAND4xp25_ASAP7_75t_SL g503 ( .A(n_452), .B(n_420), .C(n_418), .D(n_55), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_429), .B(n_434), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_450), .B(n_219), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_427), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_451), .B(n_53), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_464), .B(n_54), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_438), .A2(n_219), .B1(n_202), .B2(n_178), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_453), .Y(n_510) );
INVxp33_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_466), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_446), .B(n_57), .Y(n_513) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_444), .B(n_59), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_483), .B(n_444), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_480), .B(n_433), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_469), .B(n_439), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_506), .A2(n_487), .B1(n_484), .B2(n_501), .C(n_504), .Y(n_518) );
OR2x6_ASAP7_75t_L g519 ( .A(n_494), .B(n_454), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_481), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_473), .A2(n_441), .B1(n_439), .B2(n_323), .Y(n_522) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_479), .B(n_439), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_485), .B(n_74), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_492), .B(n_165), .C(n_170), .D(n_201), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_494), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_472), .Y(n_527) );
OAI21xp33_ASAP7_75t_L g528 ( .A1(n_493), .A2(n_205), .B(n_211), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_476), .A2(n_202), .B1(n_211), .B2(n_210), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_497), .B(n_210), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_500), .A2(n_323), .B1(n_259), .B2(n_248), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_491), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_502), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_502), .Y(n_535) );
AND2x2_ASAP7_75t_SL g536 ( .A(n_514), .B(n_210), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_513), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_488), .B(n_211), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_474), .B(n_211), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_474), .B(n_183), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_503), .A2(n_183), .B1(n_221), .B2(n_259), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_496), .A2(n_183), .B1(n_323), .B2(n_259), .Y(n_542) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_491), .B(n_170), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_478), .B(n_180), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_496), .B(n_323), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_478), .B(n_190), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_486), .B(n_190), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_512), .B(n_180), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_495), .B(n_184), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_477), .A2(n_184), .B(n_175), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_520), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_526), .Y(n_552) );
OAI22xp33_ASAP7_75t_SL g553 ( .A1(n_519), .A2(n_471), .B1(n_490), .B2(n_510), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_537), .A2(n_514), .B1(n_513), .B2(n_511), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_533), .B(n_489), .Y(n_555) );
OAI322xp33_ASAP7_75t_L g556 ( .A1(n_516), .A2(n_471), .A3(n_509), .B1(n_507), .B2(n_508), .C1(n_489), .C2(n_498), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_518), .B(n_470), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_533), .B(n_470), .Y(n_558) );
XNOR2xp5_ASAP7_75t_L g559 ( .A(n_543), .B(n_511), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_521), .B(n_499), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_535), .B(n_508), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g562 ( .A(n_536), .B(n_505), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_534), .B(n_527), .Y(n_563) );
AOI221xp5_ASAP7_75t_SL g564 ( .A1(n_520), .A2(n_223), .B1(n_249), .B2(n_277), .C(n_175), .Y(n_564) );
XOR2xp5_ASAP7_75t_L g565 ( .A(n_532), .B(n_223), .Y(n_565) );
OAI21xp33_ASAP7_75t_SL g566 ( .A1(n_519), .A2(n_199), .B(n_221), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_515), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_541), .A2(n_223), .B(n_249), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_528), .B(n_249), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_519), .B(n_277), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_517), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_538), .Y(n_572) );
XOR2x2_ASAP7_75t_L g573 ( .A(n_524), .B(n_546), .Y(n_573) );
XNOR2x2_ASAP7_75t_L g574 ( .A(n_525), .B(n_545), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_530), .Y(n_575) );
AOI31xp33_ASAP7_75t_L g576 ( .A1(n_550), .A2(n_544), .A3(n_529), .B(n_549), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_548), .Y(n_577) );
OA22x2_ASAP7_75t_L g578 ( .A1(n_522), .A2(n_523), .B1(n_542), .B2(n_550), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_531), .A2(n_539), .B1(n_540), .B2(n_547), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_548), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
OAI221xp5_ASAP7_75t_SL g582 ( .A1(n_518), .A2(n_392), .B1(n_537), .B2(n_516), .C(n_506), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_518), .A2(n_392), .B1(n_537), .B2(n_506), .C(n_543), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_537), .A2(n_392), .B1(n_483), .B2(n_518), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_516), .B(n_521), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_518), .B(n_516), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_518), .A2(n_392), .B1(n_506), .B2(n_391), .C(n_516), .Y(n_587) );
XNOR2x1_ASAP7_75t_L g588 ( .A(n_543), .B(n_473), .Y(n_588) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_543), .B(n_473), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_521), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_521), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g592 ( .A1(n_582), .A2(n_586), .B(n_584), .C(n_587), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
NAND4xp75_ASAP7_75t_L g594 ( .A(n_557), .B(n_560), .C(n_558), .D(n_574), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_591), .Y(n_595) );
AO22x2_ASAP7_75t_L g596 ( .A1(n_551), .A2(n_588), .B1(n_552), .B2(n_585), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_559), .B(n_589), .Y(n_597) );
OAI211xp5_ASAP7_75t_SL g598 ( .A1(n_583), .A2(n_585), .B(n_554), .C(n_575), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_571), .B(n_558), .Y(n_599) );
AOI31xp33_ASAP7_75t_L g600 ( .A1(n_559), .A2(n_565), .A3(n_562), .B(n_577), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_571), .B(n_572), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_590), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_553), .A2(n_556), .B(n_579), .C(n_562), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_578), .A2(n_553), .B(n_565), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_595), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_604), .A2(n_556), .B(n_577), .C(n_566), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_600), .A2(n_569), .B(n_573), .Y(n_607) );
OAI211xp5_ASAP7_75t_SL g608 ( .A1(n_592), .A2(n_567), .B(n_566), .C(n_581), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_601), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_596), .A2(n_580), .B1(n_572), .B2(n_576), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g611 ( .A(n_603), .B(n_564), .C(n_555), .D(n_561), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_596), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_605), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_609), .Y(n_614) );
NAND5xp2_ASAP7_75t_L g615 ( .A(n_607), .B(n_594), .C(n_570), .D(n_597), .E(n_568), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_609), .Y(n_616) );
NAND5xp2_ASAP7_75t_L g617 ( .A(n_614), .B(n_606), .C(n_612), .D(n_611), .E(n_610), .Y(n_617) );
XOR2xp5_ASAP7_75t_L g618 ( .A(n_616), .B(n_593), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_613), .B(n_602), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_618), .B(n_613), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_619), .B(n_615), .Y(n_621) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_620), .Y(n_622) );
XNOR2x1_ASAP7_75t_L g623 ( .A(n_622), .B(n_621), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_623), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_624), .A2(n_617), .B1(n_598), .B2(n_608), .C(n_599), .Y(n_625) );
endmodule