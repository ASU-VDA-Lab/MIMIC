module fake_jpeg_19664_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_22),
.B1(n_28),
.B2(n_23),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_18),
.C(n_11),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_41),
.B1(n_31),
.B2(n_23),
.Y(n_47)
);

OAI22x1_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_25),
.B1(n_23),
.B2(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_29),
.B1(n_30),
.B2(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_14),
.B1(n_19),
.B2(n_13),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_36),
.B(n_38),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_44),
.B(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_16),
.B1(n_33),
.B2(n_31),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_26),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_44),
.B1(n_37),
.B2(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_59),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_47),
.B1(n_44),
.B2(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_66),
.B1(n_56),
.B2(n_24),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_46),
.C(n_42),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_24),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_60),
.B(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_64),
.B1(n_63),
.B2(n_58),
.C(n_60),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_76),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_56),
.B1(n_62),
.B2(n_65),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_82),
.B(n_67),
.C(n_21),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_87),
.B(n_7),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_81),
.B(n_84),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_70),
.C(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_93),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_89),
.B1(n_37),
.B2(n_3),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.C(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_10),
.C(n_2),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.C(n_0),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_103),
.B(n_4),
.Y(n_106)
);


endmodule