module real_aes_9032_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g466 ( .A(n_0), .Y(n_466) );
INVx1_ASAP7_75t_L g501 ( .A(n_1), .Y(n_501) );
INVx1_ASAP7_75t_L g207 ( .A(n_2), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_3), .A2(n_37), .B1(n_168), .B2(n_531), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g175 ( .A1(n_4), .A2(n_149), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_5), .B(n_142), .Y(n_514) );
AND2x6_ASAP7_75t_L g154 ( .A(n_6), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_7), .A2(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_8), .B(n_38), .Y(n_467) );
INVx1_ASAP7_75t_L g182 ( .A(n_9), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_10), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g147 ( .A(n_11), .Y(n_147) );
INVx1_ASAP7_75t_L g495 ( .A(n_12), .Y(n_495) );
INVx1_ASAP7_75t_L g263 ( .A(n_13), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_14), .B(n_190), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_15), .B(n_143), .Y(n_572) );
AO32x2_ASAP7_75t_L g544 ( .A1(n_16), .A2(n_142), .A3(n_187), .B1(n_523), .B2(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_17), .A2(n_63), .B1(n_131), .B2(n_132), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_17), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_18), .B(n_168), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_19), .B(n_163), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_20), .B(n_143), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_21), .A2(n_51), .B1(n_168), .B2(n_531), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_22), .B(n_149), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_23), .A2(n_80), .B1(n_168), .B2(n_190), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_24), .B(n_168), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_25), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_26), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_28), .B(n_184), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_29), .B(n_180), .Y(n_209) );
INVx1_ASAP7_75t_L g196 ( .A(n_30), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_31), .A2(n_32), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
INVxp67_ASAP7_75t_L g125 ( .A(n_32), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_32), .B(n_184), .Y(n_561) );
INVx2_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_34), .B(n_168), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_35), .B(n_184), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_36), .A2(n_154), .B(n_158), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_38), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g194 ( .A(n_39), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_40), .A2(n_475), .B1(n_478), .B2(n_479), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_40), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_41), .B(n_180), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_42), .A2(n_105), .B1(n_106), .B2(n_117), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_43), .B(n_168), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_44), .A2(n_90), .B1(n_226), .B2(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_45), .B(n_168), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_46), .B(n_168), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_47), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_48), .A2(n_70), .B1(n_476), .B2(n_477), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_48), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_49), .B(n_500), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_50), .B(n_149), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_52), .A2(n_61), .B1(n_168), .B2(n_190), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_53), .A2(n_158), .B1(n_190), .B2(n_192), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_54), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_55), .B(n_168), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_56), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_57), .B(n_168), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_58), .A2(n_167), .B(n_179), .C(n_181), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_59), .Y(n_239) );
INVx1_ASAP7_75t_L g177 ( .A(n_60), .Y(n_177) );
INVx1_ASAP7_75t_L g155 ( .A(n_62), .Y(n_155) );
INVx1_ASAP7_75t_L g131 ( .A(n_63), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_64), .B(n_168), .Y(n_502) );
INVx1_ASAP7_75t_L g146 ( .A(n_65), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_67), .A2(n_142), .A3(n_243), .B1(n_523), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g521 ( .A(n_68), .Y(n_521) );
INVx1_ASAP7_75t_L g556 ( .A(n_69), .Y(n_556) );
INVx1_ASAP7_75t_L g476 ( .A(n_70), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_SL g162 ( .A1(n_71), .A2(n_163), .B(n_164), .C(n_167), .Y(n_162) );
INVxp67_ASAP7_75t_L g165 ( .A(n_72), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_73), .B(n_190), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_74), .A2(n_473), .B1(n_474), .B2(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_74), .Y(n_473) );
INVx1_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_76), .B(n_462), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_77), .A2(n_464), .B1(n_471), .B2(n_775), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_78), .Y(n_200) );
INVx1_ASAP7_75t_L g232 ( .A(n_79), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_81), .A2(n_154), .B(n_158), .C(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_82), .B(n_531), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_83), .B(n_190), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_84), .B(n_208), .Y(n_222) );
INVx2_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_86), .B(n_163), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_87), .B(n_190), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_88), .A2(n_154), .B(n_158), .C(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
OR2x2_ASAP7_75t_L g463 ( .A(n_89), .B(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_91), .A2(n_103), .B1(n_190), .B2(n_191), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_92), .B(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_93), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_94), .A2(n_154), .B(n_158), .C(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_95), .Y(n_253) );
INVx1_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_97), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_98), .B(n_208), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_99), .B(n_190), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_100), .B(n_142), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_101), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_102), .A2(n_149), .B(n_156), .Y(n_148) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_SL g481 ( .A1(n_113), .A2(n_133), .B1(n_482), .B2(n_774), .Y(n_481) );
INVx2_ASAP7_75t_L g774 ( .A(n_113), .Y(n_774) );
NOR2x2_ASAP7_75t_L g777 ( .A(n_113), .B(n_464), .Y(n_777) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_469), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g779 ( .A(n_121), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_460), .B(n_468), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B1(n_128), .B2(n_459), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_124), .Y(n_459) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B1(n_133), .B2(n_458), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g458 ( .A(n_133), .Y(n_458) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND4x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_376), .C(n_423), .D(n_443), .Y(n_134) );
NOR3xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_306), .C(n_331), .Y(n_135) );
OAI211xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_214), .B(n_266), .C(n_296), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_185), .Y(n_138) );
INVx3_ASAP7_75t_SL g348 ( .A(n_139), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_139), .B(n_279), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_139), .B(n_201), .Y(n_429) );
AND2x2_ASAP7_75t_L g452 ( .A(n_139), .B(n_318), .Y(n_452) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_173), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g270 ( .A(n_141), .B(n_174), .Y(n_270) );
INVx3_ASAP7_75t_L g283 ( .A(n_141), .Y(n_283) );
AND2x2_ASAP7_75t_L g288 ( .A(n_141), .B(n_173), .Y(n_288) );
OR2x2_ASAP7_75t_L g339 ( .A(n_141), .B(n_280), .Y(n_339) );
BUFx2_ASAP7_75t_L g359 ( .A(n_141), .Y(n_359) );
AND2x2_ASAP7_75t_L g369 ( .A(n_141), .B(n_280), .Y(n_369) );
AND2x2_ASAP7_75t_L g375 ( .A(n_141), .B(n_186), .Y(n_375) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_170), .Y(n_141) );
INVx4_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_142), .A2(n_507), .B(n_514), .Y(n_506) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_144), .B(n_145), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx2_ASAP7_75t_L g257 ( .A(n_149), .Y(n_257) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_150), .B(n_154), .Y(n_198) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g500 ( .A(n_151), .Y(n_500) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
INVx1_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
INVx1_ASAP7_75t_L g163 ( .A(n_153), .Y(n_163) );
INVx3_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx4_ASAP7_75t_SL g169 ( .A(n_154), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_154), .A2(n_494), .B(n_498), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_154), .A2(n_508), .B(n_511), .Y(n_507) );
BUFx3_ASAP7_75t_L g523 ( .A(n_154), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_154), .A2(n_536), .B(n_540), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_154), .A2(n_555), .B(n_558), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_161), .B(n_162), .C(n_169), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_157), .A2(n_169), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_157), .A2(n_169), .B(n_259), .C(n_260), .Y(n_258) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
BUFx3_ASAP7_75t_L g226 ( .A(n_159), .Y(n_226) );
INVx1_ASAP7_75t_L g531 ( .A(n_159), .Y(n_531) );
INVx1_ASAP7_75t_L g539 ( .A(n_163), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_166), .B(n_182), .Y(n_181) );
INVx5_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g529 ( .A1(n_166), .A2(n_180), .B1(n_530), .B2(n_532), .Y(n_529) );
O2A1O1Ixp5_ASAP7_75t_SL g555 ( .A1(n_167), .A2(n_208), .B(n_556), .C(n_557), .Y(n_555) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_169), .A2(n_189), .B1(n_197), .B2(n_198), .Y(n_188) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_171), .A2(n_175), .B(n_183), .Y(n_174) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g228 ( .A(n_172), .B(n_229), .Y(n_228) );
AO21x1_ASAP7_75t_L g567 ( .A1(n_172), .A2(n_568), .B(n_571), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_172), .B(n_523), .C(n_568), .Y(n_586) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_174), .B(n_280), .Y(n_294) );
INVx2_ASAP7_75t_L g304 ( .A(n_174), .Y(n_304) );
AND2x2_ASAP7_75t_L g317 ( .A(n_174), .B(n_283), .Y(n_317) );
OR2x2_ASAP7_75t_L g328 ( .A(n_174), .B(n_280), .Y(n_328) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_174), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g386 ( .A(n_174), .Y(n_386) );
AND2x2_ASAP7_75t_L g432 ( .A(n_174), .B(n_186), .Y(n_432) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_179), .A2(n_499), .B(n_521), .C(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_179), .A2(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_180), .A2(n_503), .B1(n_546), .B2(n_547), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_180), .A2(n_503), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g213 ( .A(n_184), .Y(n_213) );
INVx2_ASAP7_75t_L g243 ( .A(n_184), .Y(n_243) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_184), .A2(n_256), .B(n_265), .Y(n_255) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_184), .A2(n_535), .B(n_543), .Y(n_534) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_184), .A2(n_554), .B(n_561), .Y(n_553) );
INVx3_ASAP7_75t_SL g305 ( .A(n_185), .Y(n_305) );
OR2x2_ASAP7_75t_L g358 ( .A(n_185), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_201), .Y(n_185) );
INVx3_ASAP7_75t_L g280 ( .A(n_186), .Y(n_280) );
AND2x2_ASAP7_75t_L g347 ( .A(n_186), .B(n_202), .Y(n_347) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_186), .Y(n_415) );
AOI33xp33_ASAP7_75t_L g419 ( .A1(n_186), .A2(n_348), .A3(n_355), .B1(n_364), .B2(n_420), .B3(n_421), .Y(n_419) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_199), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_187), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_187), .A2(n_203), .B(n_211), .Y(n_202) );
INVx2_ASAP7_75t_L g227 ( .A(n_187), .Y(n_227) );
INVx2_ASAP7_75t_L g210 ( .A(n_190), .Y(n_210) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g195 ( .A(n_193), .Y(n_195) );
INVx4_ASAP7_75t_L g261 ( .A(n_193), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_232), .B(n_233), .Y(n_231) );
INVx1_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_201), .B(n_283), .Y(n_282) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_201), .B(n_343), .C(n_345), .Y(n_342) );
AND2x2_ASAP7_75t_L g368 ( .A(n_201), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_201), .B(n_375), .Y(n_378) );
AND2x2_ASAP7_75t_L g431 ( .A(n_201), .B(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
OR2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_280), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .C(n_210), .Y(n_206) );
INVx2_ASAP7_75t_L g503 ( .A(n_208), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_208), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_208), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_210), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_213), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_213), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_240), .Y(n_214) );
AOI32xp33_ASAP7_75t_L g332 ( .A1(n_215), .A2(n_333), .A3(n_335), .B1(n_337), .B2(n_340), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_215), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g435 ( .A(n_215), .Y(n_435) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_351), .Y(n_367) );
AND2x2_ASAP7_75t_L g387 ( .A(n_216), .B(n_313), .Y(n_387) );
AND2x2_ASAP7_75t_L g455 ( .A(n_216), .B(n_373), .Y(n_455) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_230), .Y(n_216) );
INVx3_ASAP7_75t_L g276 ( .A(n_217), .Y(n_276) );
AND2x2_ASAP7_75t_L g290 ( .A(n_217), .B(n_274), .Y(n_290) );
OR2x2_ASAP7_75t_L g295 ( .A(n_217), .B(n_273), .Y(n_295) );
INVx1_ASAP7_75t_L g302 ( .A(n_217), .Y(n_302) );
AND2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_284), .Y(n_310) );
AND2x2_ASAP7_75t_L g312 ( .A(n_217), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_217), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g365 ( .A(n_217), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_217), .B(n_450), .Y(n_449) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
AOI21xp5_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_220), .B(n_227), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_224), .A2(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
INVx1_ASAP7_75t_L g237 ( .A(n_227), .Y(n_237) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_227), .A2(n_493), .B(n_504), .Y(n_492) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_227), .A2(n_516), .B(n_524), .Y(n_515) );
INVx2_ASAP7_75t_L g274 ( .A(n_230), .Y(n_274) );
AND2x2_ASAP7_75t_L g320 ( .A(n_230), .B(n_241), .Y(n_320) );
AND2x2_ASAP7_75t_L g330 ( .A(n_230), .B(n_255), .Y(n_330) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_237), .B(n_238), .Y(n_230) );
INVx2_ASAP7_75t_L g450 ( .A(n_240), .Y(n_450) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_254), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_241), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g291 ( .A(n_241), .Y(n_291) );
AND2x2_ASAP7_75t_L g335 ( .A(n_241), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g351 ( .A(n_241), .B(n_314), .Y(n_351) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g299 ( .A(n_242), .Y(n_299) );
AND2x2_ASAP7_75t_L g313 ( .A(n_242), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g364 ( .A(n_242), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_242), .B(n_274), .Y(n_396) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g275 ( .A(n_254), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g336 ( .A(n_254), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_254), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g373 ( .A(n_254), .Y(n_373) );
INVx1_ASAP7_75t_L g406 ( .A(n_254), .Y(n_406) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g284 ( .A(n_255), .B(n_274), .Y(n_284) );
INVx1_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_261), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g497 ( .A(n_261), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_261), .A2(n_559), .B(n_560), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_271), .B1(n_277), .B2(n_284), .C(n_285), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_268), .B(n_288), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_268), .B(n_351), .Y(n_428) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_270), .B(n_318), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_270), .B(n_279), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_270), .B(n_293), .Y(n_422) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g344 ( .A(n_274), .Y(n_344) );
AND2x2_ASAP7_75t_L g319 ( .A(n_275), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g397 ( .A(n_275), .Y(n_397) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_276), .B(n_299), .Y(n_345) );
AND2x2_ASAP7_75t_L g409 ( .A(n_276), .B(n_335), .Y(n_409) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g318 ( .A(n_280), .B(n_287), .Y(n_318) );
AND2x2_ASAP7_75t_L g414 ( .A(n_281), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_283), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_284), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_284), .B(n_291), .Y(n_379) );
AND2x2_ASAP7_75t_L g399 ( .A(n_284), .B(n_299), .Y(n_399) );
AND2x2_ASAP7_75t_L g420 ( .A(n_284), .B(n_364), .Y(n_420) );
OAI32xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .A3(n_291), .B1(n_292), .B2(n_295), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_SL g293 ( .A(n_287), .Y(n_293) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_287), .B(n_317), .Y(n_334) );
OR2x2_ASAP7_75t_L g338 ( .A(n_287), .B(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_287), .B(n_386), .Y(n_439) );
INVx1_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
OAI221xp5_ASAP7_75t_SL g425 ( .A1(n_289), .A2(n_380), .B1(n_426), .B2(n_429), .C(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g340 ( .A(n_290), .B(n_313), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_290), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_351), .Y(n_418) );
INVxp67_ASAP7_75t_L g354 ( .A(n_291), .Y(n_354) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g424 ( .A(n_293), .B(n_411), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_293), .B(n_374), .Y(n_447) );
INVx1_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_295), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g440 ( .A(n_295), .B(n_441), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_300), .B(n_303), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_298), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g393 ( .A(n_302), .B(n_313), .Y(n_393) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g411 ( .A(n_304), .B(n_369), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_304), .B(n_368), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_305), .B(n_317), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_311), .C(n_321), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_307), .A2(n_342), .B1(n_346), .B2(n_349), .C(n_352), .Y(n_341) );
AOI31xp33_ASAP7_75t_L g436 ( .A1(n_307), .A2(n_437), .A3(n_438), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_317), .B2(n_319), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g437 ( .A(n_317), .Y(n_437) );
INVx1_ASAP7_75t_L g400 ( .A(n_318), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_320), .A2(n_444), .B(n_446), .C(n_448), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_325), .B2(n_329), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_326), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_328), .A2(n_362), .B1(n_381), .B2(n_417), .C(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g412 ( .A(n_329), .Y(n_412) );
INVx1_ASAP7_75t_L g366 ( .A(n_330), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g331 ( .A(n_332), .B(n_341), .C(n_356), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g382 ( .A1(n_333), .A2(n_383), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_335), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g442 ( .A(n_336), .Y(n_442) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_363), .Y(n_380) );
INVx1_ASAP7_75t_L g355 ( .A(n_344), .Y(n_355) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g353 ( .A(n_347), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_347), .B(n_385), .Y(n_384) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .C(n_354), .D(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B1(n_367), .B2(n_368), .C1(n_370), .C2(n_374), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g454 ( .A(n_358), .Y(n_454) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_370), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_375), .A2(n_431), .B(n_433), .Y(n_430) );
NOR4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_388), .C(n_401), .D(n_416), .Y(n_376) );
OAI221xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_379), .B1(n_380), .B2(n_381), .C(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g457 ( .A(n_378), .Y(n_457) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_385), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B1(n_394), .B2(n_395), .C1(n_398), .C2(n_400), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_424), .B(n_425), .C(n_436), .Y(n_423) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OAI222xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_407), .B1(n_408), .B2(n_410), .C1(n_412), .C2(n_413), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_418), .A2(n_421), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI211xp5_ASAP7_75t_SL g448 ( .A1(n_449), .A2(n_451), .B(n_453), .C(n_456), .Y(n_448) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_468), .A2(n_470), .B(n_778), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_474), .Y(n_480) );
INVx1_ASAP7_75t_L g478 ( .A(n_475), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_484), .B(n_740), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_644), .C(n_728), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_587), .C(n_609), .D(n_625), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_525), .B1(n_548), .B2(n_566), .C(n_573), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_505), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_489), .B(n_566), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_489), .B(n_627), .C(n_640), .D(n_642), .Y(n_639) );
INVxp67_ASAP7_75t_L g756 ( .A(n_489), .Y(n_756) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g638 ( .A(n_490), .B(n_576), .Y(n_638) );
AND2x2_ASAP7_75t_L g662 ( .A(n_490), .B(n_505), .Y(n_662) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g629 ( .A(n_491), .B(n_565), .Y(n_629) );
AND2x2_ASAP7_75t_L g669 ( .A(n_491), .B(n_650), .Y(n_669) );
AND2x2_ASAP7_75t_L g686 ( .A(n_491), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_491), .B(n_506), .Y(n_710) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g593 ( .A(n_492), .B(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_492), .B(n_515), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_501), .B(n_502), .C(n_503), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_503), .A2(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g596 ( .A(n_505), .B(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_505), .A2(n_646), .B1(n_649), .B2(n_651), .C(n_655), .Y(n_645) );
AND2x2_ASAP7_75t_L g704 ( .A(n_505), .B(n_669), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_505), .B(n_686), .Y(n_738) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx3_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
AND2x2_ASAP7_75t_L g613 ( .A(n_506), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g667 ( .A(n_506), .B(n_582), .Y(n_667) );
AND2x2_ASAP7_75t_L g725 ( .A(n_506), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g582 ( .A(n_515), .Y(n_582) );
INVx1_ASAP7_75t_L g637 ( .A(n_515), .Y(n_637) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_515), .Y(n_643) );
AND2x2_ASAP7_75t_L g688 ( .A(n_515), .B(n_565), .Y(n_688) );
OR2x2_ASAP7_75t_L g727 ( .A(n_515), .B(n_567), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_520), .B(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_525), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_533), .Y(n_525) );
AND2x2_ASAP7_75t_L g723 ( .A(n_526), .B(n_720), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_526), .B(n_705), .Y(n_755) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g654 ( .A(n_527), .B(n_578), .Y(n_654) );
AND2x2_ASAP7_75t_L g703 ( .A(n_527), .B(n_551), .Y(n_703) );
INVx1_ASAP7_75t_L g749 ( .A(n_527), .Y(n_749) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_528), .Y(n_563) );
AND2x2_ASAP7_75t_L g604 ( .A(n_528), .B(n_578), .Y(n_604) );
INVx1_ASAP7_75t_L g621 ( .A(n_528), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_528), .B(n_544), .Y(n_627) );
AND2x2_ASAP7_75t_L g695 ( .A(n_533), .B(n_603), .Y(n_695) );
INVx2_ASAP7_75t_L g760 ( .A(n_533), .Y(n_760) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_544), .Y(n_533) );
AND2x2_ASAP7_75t_L g577 ( .A(n_534), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_552), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_534), .B(n_551), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_534), .Y(n_624) );
INVx1_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_534), .Y(n_653) );
INVx2_ASAP7_75t_L g721 ( .A(n_534), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
BUFx2_ASAP7_75t_L g675 ( .A(n_544), .Y(n_675) );
AND2x2_ASAP7_75t_L g720 ( .A(n_544), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_550), .B(n_657), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_550), .A2(n_719), .B(n_733), .Y(n_743) );
AND2x2_ASAP7_75t_L g768 ( .A(n_550), .B(n_654), .Y(n_768) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g690 ( .A(n_552), .Y(n_690) );
AND2x2_ASAP7_75t_L g719 ( .A(n_552), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
INVx2_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g576 ( .A(n_563), .Y(n_576) );
OR2x2_ASAP7_75t_L g589 ( .A(n_563), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g657 ( .A(n_563), .B(n_653), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_563), .B(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g758 ( .A(n_563), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_563), .B(n_695), .Y(n_770) );
AND2x2_ASAP7_75t_L g649 ( .A(n_564), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g672 ( .A(n_564), .B(n_566), .Y(n_672) );
INVx2_ASAP7_75t_L g584 ( .A(n_565), .Y(n_584) );
AND2x2_ASAP7_75t_L g612 ( .A(n_565), .B(n_585), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_565), .B(n_637), .Y(n_693) );
AND2x2_ASAP7_75t_L g607 ( .A(n_566), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g754 ( .A(n_566), .Y(n_754) );
AND2x2_ASAP7_75t_L g766 ( .A(n_566), .B(n_629), .Y(n_766) );
AND2x2_ASAP7_75t_L g592 ( .A(n_567), .B(n_582), .Y(n_592) );
INVx1_ASAP7_75t_L g687 ( .A(n_567), .Y(n_687) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_576), .B(n_623), .Y(n_632) );
OR2x2_ASAP7_75t_L g764 ( .A(n_576), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g681 ( .A(n_577), .B(n_622), .Y(n_681) );
AND2x2_ASAP7_75t_L g689 ( .A(n_577), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g748 ( .A(n_577), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g772 ( .A(n_577), .B(n_619), .Y(n_772) );
NOR2xp67_ASAP7_75t_L g730 ( .A(n_578), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g759 ( .A(n_578), .B(n_622), .Y(n_759) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g611 ( .A(n_581), .B(n_612), .Y(n_611) );
INVxp67_ASAP7_75t_L g773 ( .A(n_581), .Y(n_773) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g608 ( .A(n_584), .Y(n_608) );
AND2x2_ASAP7_75t_L g659 ( .A(n_584), .B(n_592), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_584), .B(n_727), .Y(n_753) );
INVx2_ASAP7_75t_L g598 ( .A(n_585), .Y(n_598) );
INVx3_ASAP7_75t_L g650 ( .A(n_585), .Y(n_650) );
OR2x2_ASAP7_75t_L g678 ( .A(n_585), .B(n_679), .Y(n_678) );
AOI311xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .A3(n_593), .B(n_594), .C(n_605), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_588), .A2(n_626), .B(n_628), .C(n_630), .Y(n_625) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g610 ( .A(n_590), .Y(n_610) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g628 ( .A(n_592), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_592), .B(n_608), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_592), .B(n_593), .Y(n_761) );
AND2x2_ASAP7_75t_L g683 ( .A(n_593), .B(n_597), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B(n_600), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g741 ( .A(n_597), .B(n_629), .Y(n_741) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_598), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g635 ( .A(n_598), .Y(n_635) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g626 ( .A(n_602), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g671 ( .A(n_604), .Y(n_671) );
AND2x4_ASAP7_75t_L g733 ( .A(n_604), .B(n_702), .Y(n_733) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_607), .A2(n_673), .B1(n_685), .B2(n_689), .C1(n_691), .C2(n_695), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_613), .C(n_616), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_610), .B(n_654), .Y(n_677) );
INVx1_ASAP7_75t_L g699 ( .A(n_612), .Y(n_699) );
INVx1_ASAP7_75t_L g633 ( .A(n_614), .Y(n_633) );
OR2x2_ASAP7_75t_L g698 ( .A(n_615), .B(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .B(n_623), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_617), .B(n_635), .C(n_636), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_617), .A2(n_654), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_621), .Y(n_674) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_622), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_622), .Y(n_747) );
INVx2_ASAP7_75t_L g705 ( .A(n_623), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_627), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g679 ( .A(n_629), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_634), .B2(n_638), .C(n_639), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_633), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g767 ( .A(n_633), .Y(n_767) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g648 ( .A(n_640), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_640), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g706 ( .A(n_640), .B(n_654), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_640), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g739 ( .A(n_640), .B(n_674), .Y(n_739) );
BUFx3_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_684), .D(n_696), .E(n_711), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI32xp33_ASAP7_75t_L g736 ( .A1(n_648), .A2(n_675), .A3(n_691), .B1(n_737), .B2(n_739), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_650), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g660 ( .A(n_654), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_670), .B1(n_672), .B2(n_673), .C(n_676), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g735 ( .A(n_667), .B(n_686), .Y(n_735) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_672), .A2(n_733), .B1(n_751), .B2(n_756), .C(n_757), .Y(n_750) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx2_ASAP7_75t_L g716 ( .A(n_675), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g694 ( .A(n_686), .Y(n_694) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_707), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_705), .A2(n_752), .B1(n_754), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .B(n_724), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g765 ( .A(n_720), .Y(n_765) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B(n_734), .C(n_736), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B(n_744), .C(n_769), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_741), .Y(n_745) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_750), .C(n_762), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_761), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
endmodule