module fake_jpeg_15121_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_46),
.B1(n_59),
.B2(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_73),
.B1(n_79),
.B2(n_82),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_72),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_53),
.B1(n_51),
.B2(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_58),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_60),
.B1(n_55),
.B2(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_50),
.B1(n_45),
.B2(n_5),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_81),
.C(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_71),
.B1(n_7),
.B2(n_8),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_81),
.B(n_9),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.C(n_99),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_3),
.C(n_11),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_12),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_13),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_15),
.A3(n_16),
.B1(n_18),
.B2(n_20),
.C1(n_23),
.C2(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_26),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_33),
.Y(n_112)
);


endmodule