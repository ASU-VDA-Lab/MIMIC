module fake_jpeg_3391_n_178 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx8_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_55),
.Y(n_73)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_21),
.B(n_1),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_2),
.C(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_5),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_19),
.Y(n_76)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_5),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_29),
.A2(n_22),
.B1(n_25),
.B2(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_71),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_30),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_82),
.B1(n_69),
.B2(n_58),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_44),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_34),
.A2(n_24),
.B1(n_19),
.B2(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_32),
.B1(n_39),
.B2(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_6),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_9),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_6),
.B1(n_8),
.B2(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_76),
.B1(n_70),
.B2(n_62),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_109),
.B1(n_99),
.B2(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_65),
.B1(n_75),
.B2(n_80),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_106),
.B1(n_89),
.B2(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_84),
.C(n_75),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_104),
.C(n_107),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_60),
.CI(n_85),
.CON(n_102),
.SN(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_85),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_107),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_63),
.B1(n_74),
.B2(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_56),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_90),
.Y(n_115)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_101),
.C(n_88),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_99),
.B1(n_95),
.B2(n_102),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_102),
.B1(n_100),
.B2(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_134),
.C(n_116),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_137),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_125),
.C(n_115),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_124),
.B1(n_122),
.B2(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_129),
.B1(n_114),
.B2(n_123),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_118),
.B(n_116),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_136),
.B1(n_111),
.B2(n_122),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_136),
.B1(n_111),
.B2(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_157),
.B1(n_143),
.B2(n_110),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_136),
.A3(n_131),
.B1(n_122),
.B2(n_130),
.C(n_139),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_154),
.B(n_153),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_130),
.B(n_145),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_142),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_150),
.B1(n_162),
.B2(n_158),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_151),
.B1(n_139),
.B2(n_121),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_160),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_164),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_167),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_121),
.Y(n_178)
);


endmodule