module fake_jpeg_2190_n_611 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_58),
.Y(n_167)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_79),
.Y(n_151)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_62),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_74),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_26),
.B(n_39),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_64),
.B(n_92),
.C(n_88),
.Y(n_181)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_1),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_76),
.B(n_99),
.Y(n_199)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_1),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_82),
.B(n_115),
.Y(n_155)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_2),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_21),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_38),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_125),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_4),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_20),
.B1(n_53),
.B2(n_40),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_146),
.B1(n_197),
.B2(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_23),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_136),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_60),
.B(n_23),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_133),
.B(n_134),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_57),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_53),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_38),
.B1(n_48),
.B2(n_44),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_141),
.A2(n_196),
.B1(n_78),
.B2(n_84),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_48),
.B1(n_44),
.B2(n_40),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_145),
.A2(n_154),
.B1(n_190),
.B2(n_16),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_32),
.B1(n_28),
.B2(n_55),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_48),
.B1(n_44),
.B2(n_32),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_64),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_161),
.B(n_202),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_87),
.A2(n_55),
.A3(n_48),
.B1(n_44),
.B2(n_28),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_164),
.A2(n_102),
.B(n_121),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_111),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_178),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_105),
.A2(n_46),
.B(n_5),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_17),
.B(n_18),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_106),
.B(n_4),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_192),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_81),
.B(n_5),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_184),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_68),
.B(n_6),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_112),
.A2(n_46),
.B1(n_8),
.B2(n_9),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_72),
.B(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_204),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_108),
.A2(n_46),
.B1(n_10),
.B2(n_12),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_46),
.B1(n_10),
.B2(n_12),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_62),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_85),
.B(n_18),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_124),
.A2(n_9),
.B1(n_13),
.B2(n_16),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_212),
.B1(n_18),
.B2(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_69),
.B(n_9),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_207),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_70),
.B(n_13),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_168),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_73),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_215),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_216),
.B(n_233),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_127),
.A2(n_89),
.B1(n_93),
.B2(n_90),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_218),
.A2(n_263),
.B1(n_269),
.B2(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_220),
.Y(n_289)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_222),
.A2(n_239),
.B1(n_240),
.B2(n_250),
.Y(n_312)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_223),
.Y(n_290)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_224),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_225),
.Y(n_331)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_226),
.Y(n_344)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_230),
.B(n_231),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_188),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_132),
.A2(n_18),
.B1(n_163),
.B2(n_155),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_235),
.A2(n_241),
.B1(n_252),
.B2(n_285),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_236),
.B(n_238),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_148),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_141),
.A2(n_196),
.B1(n_144),
.B2(n_142),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_132),
.A2(n_163),
.B1(n_187),
.B2(n_159),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_243),
.Y(n_341)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_191),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_152),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_249),
.B(n_253),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_173),
.A2(n_203),
.B1(n_151),
.B2(n_171),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_255),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_199),
.B1(n_206),
.B2(n_185),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_166),
.C(n_232),
.Y(n_304)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_266),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_156),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_259),
.B(n_270),
.Y(n_327)
);

AO22x2_ASAP7_75t_L g260 ( 
.A1(n_158),
.A2(n_138),
.B1(n_139),
.B2(n_186),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_260),
.B(n_222),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_130),
.B(n_176),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_273),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_156),
.A2(n_147),
.B1(n_169),
.B2(n_182),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g264 ( 
.A1(n_135),
.A2(n_168),
.B1(n_174),
.B2(n_186),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_260),
.Y(n_316)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_153),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_126),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_267),
.B(n_268),
.Y(n_342)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_135),
.A2(n_157),
.B1(n_129),
.B2(n_137),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_189),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_126),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_271),
.B(n_272),
.Y(n_328)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_129),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_274),
.Y(n_324)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_182),
.Y(n_276)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_149),
.B(n_213),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_277),
.B(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_150),
.B(n_198),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_150),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_198),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.Y(n_291)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_180),
.B(n_165),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_282),
.B(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_200),
.A2(n_213),
.B1(n_180),
.B2(n_165),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_286),
.Y(n_343)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_166),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_288),
.A2(n_215),
.B1(n_223),
.B2(n_242),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_231),
.A2(n_143),
.B(n_166),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_299),
.A2(n_246),
.B(n_286),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_300),
.B(n_296),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_307),
.A2(n_316),
.B1(n_337),
.B2(n_281),
.Y(n_366)
);

BUFx24_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_237),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_319),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_252),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_264),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_338),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_282),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_215),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_225),
.A2(n_256),
.B1(n_214),
.B2(n_241),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_256),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_260),
.B(n_243),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_345),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_271),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_346),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_239),
.B(n_227),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_347),
.A2(n_365),
.B(n_376),
.Y(n_399)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_359),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_331),
.A2(n_312),
.B1(n_316),
.B2(n_338),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_355),
.A2(n_356),
.B1(n_385),
.B2(n_335),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_331),
.A2(n_275),
.B1(n_274),
.B2(n_247),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_323),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_294),
.B(n_219),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_362),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_319),
.A2(n_266),
.B1(n_217),
.B2(n_276),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_374),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_345),
.A2(n_226),
.B1(n_228),
.B2(n_287),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_367),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_366),
.A2(n_371),
.B1(n_382),
.B2(n_290),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_336),
.A2(n_248),
.B1(n_284),
.B2(n_340),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_310),
.B(n_299),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_368),
.A2(n_291),
.B(n_339),
.Y(n_405)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_300),
.A2(n_320),
.B1(n_336),
.B2(n_305),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_323),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_294),
.B(n_318),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_377),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_313),
.B(n_311),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_386),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_304),
.A2(n_295),
.B(n_320),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_380),
.A2(n_290),
.B(n_335),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_309),
.C(n_330),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_324),
.A2(n_321),
.B1(n_343),
.B2(n_334),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_387),
.Y(n_397)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_324),
.B(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_344),
.A2(n_291),
.B1(n_293),
.B2(n_341),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_290),
.B1(n_344),
.B2(n_308),
.Y(n_398)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_389),
.B(n_322),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_391),
.A2(n_421),
.B1(n_364),
.B2(n_362),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_381),
.C(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_402),
.C(n_406),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_414),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_398),
.A2(n_388),
.B1(n_349),
.B2(n_350),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_297),
.C(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_405),
.A2(n_415),
.B(n_425),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_317),
.C(n_339),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_308),
.C(n_330),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_411),
.C(n_352),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_303),
.C(n_301),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g413 ( 
.A(n_360),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_301),
.C(n_302),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_366),
.A2(n_298),
.B1(n_303),
.B2(n_315),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_375),
.B(n_315),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_422),
.B(n_346),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_302),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_424),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_298),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_368),
.A2(n_301),
.B(n_306),
.Y(n_425)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_408),
.B(n_420),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_428),
.B(n_442),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_370),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_347),
.B1(n_376),
.B2(n_351),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_434),
.B1(n_435),
.B2(n_437),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_423),
.A2(n_384),
.B1(n_369),
.B2(n_358),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_433),
.A2(n_392),
.B1(n_390),
.B2(n_418),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_411),
.A2(n_384),
.B1(n_377),
.B2(n_378),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_408),
.B(n_382),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_438),
.B(n_458),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_417),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_420),
.B(n_395),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_399),
.A2(n_384),
.B(n_365),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_443),
.A2(n_412),
.B(n_401),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_367),
.B1(n_384),
.B2(n_386),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_449),
.B1(n_457),
.B2(n_410),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_372),
.Y(n_445)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_445),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_353),
.C(n_383),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_446),
.B(n_455),
.C(n_393),
.Y(n_486)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_395),
.A2(n_407),
.B1(n_421),
.B2(n_411),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_400),
.Y(n_450)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_450),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_401),
.Y(n_451)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_422),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_454),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_400),
.B(n_359),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_396),
.B(n_402),
.C(n_406),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_387),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_419),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_356),
.B1(n_357),
.B2(n_374),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_403),
.B(n_389),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_449),
.A2(n_415),
.B1(n_407),
.B2(n_399),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_463),
.B(n_471),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_455),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_465),
.B(n_469),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_450),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_466),
.B(n_468),
.C(n_452),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_454),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_414),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_414),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_485),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_444),
.A2(n_398),
.B1(n_405),
.B2(n_417),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g505 ( 
.A1(n_472),
.A2(n_480),
.B(n_489),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_473),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_438),
.A2(n_392),
.B1(n_390),
.B2(n_418),
.Y(n_475)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_432),
.B(n_404),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_479),
.B(n_483),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_481),
.B(n_448),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_419),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_486),
.C(n_488),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_416),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_416),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_430),
.A2(n_361),
.B1(n_370),
.B2(n_385),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_487),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_435),
.A2(n_385),
.B1(n_361),
.B2(n_306),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_478),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_491),
.B(n_499),
.Y(n_536)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

INVx13_ASAP7_75t_L g493 ( 
.A(n_489),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_493),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_472),
.A2(n_436),
.B(n_443),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_495),
.A2(n_436),
.B(n_480),
.Y(n_534)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_461),
.B(n_428),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_477),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_500),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_520)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_487),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_503),
.Y(n_535)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_451),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_513),
.Y(n_526)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_470),
.Y(n_521)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_477),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_467),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_465),
.C(n_496),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_518),
.C(n_529),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_488),
.C(n_469),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_527),
.Y(n_548)
);

FAx1_ASAP7_75t_SL g523 ( 
.A(n_500),
.B(n_433),
.CI(n_463),
.CON(n_523),
.SN(n_523)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_515),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_496),
.B(n_485),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_488),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_533),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_482),
.C(n_481),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_501),
.A2(n_462),
.B1(n_459),
.B2(n_442),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_530),
.A2(n_492),
.B1(n_462),
.B2(n_459),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_506),
.A2(n_464),
.B1(n_498),
.B2(n_504),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_531),
.A2(n_506),
.B1(n_504),
.B2(n_498),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_431),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_534),
.A2(n_505),
.B(n_493),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_429),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_505),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_520),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_547),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_542),
.A2(n_546),
.B1(n_530),
.B2(n_519),
.Y(n_560)
);

OAI321xp33_ASAP7_75t_L g557 ( 
.A1(n_543),
.A2(n_525),
.A3(n_534),
.B1(n_519),
.B2(n_524),
.C(n_537),
.Y(n_557)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_535),
.A2(n_502),
.B1(n_490),
.B2(n_516),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_536),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_526),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_549),
.B(n_551),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_531),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_SL g551 ( 
.A(n_517),
.B(n_476),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_502),
.C(n_490),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_552),
.B(n_555),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_556),
.Y(n_564)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_537),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_447),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_476),
.C(n_513),
.Y(n_555)
);

AND2x2_ASAP7_75t_SL g556 ( 
.A(n_524),
.B(n_439),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_557),
.A2(n_569),
.B(n_439),
.Y(n_583)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_560),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_555),
.B(n_552),
.C(n_541),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_562),
.B(n_568),
.Y(n_580)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_563),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_445),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_494),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_567),
.B(n_544),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_542),
.A2(n_523),
.B1(n_538),
.B2(n_533),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_543),
.A2(n_523),
.B(n_514),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_541),
.B(n_528),
.C(n_529),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_548),
.C(n_540),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_553),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_574),
.Y(n_584)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_573),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_575),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_558),
.A2(n_559),
.B1(n_565),
.B2(n_560),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_579),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_568),
.A2(n_556),
.B1(n_550),
.B2(n_545),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_569),
.A2(n_556),
.B1(n_497),
.B2(n_508),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_564),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_532),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_583),
.B(n_522),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_571),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_586),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_570),
.C(n_548),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_578),
.B(n_563),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_579),
.Y(n_598)
);

AO21x1_ASAP7_75t_L g597 ( 
.A1(n_591),
.A2(n_592),
.B(n_582),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_584),
.B(n_577),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_593),
.B(n_595),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_589),
.A2(n_583),
.B(n_580),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_586),
.C(n_587),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_597),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_598),
.B(n_599),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_588),
.B(n_575),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_590),
.C(n_581),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_602),
.A2(n_564),
.B(n_540),
.Y(n_605)
);

OAI21xp33_ASAP7_75t_L g604 ( 
.A1(n_601),
.A2(n_595),
.B(n_441),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_604),
.B(n_605),
.C(n_603),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_606),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_600),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_532),
.B(n_434),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_609),
.A2(n_503),
.B(n_441),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_521),
.Y(n_611)
);


endmodule