module fake_jpeg_17331_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.C(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_19),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_18),
.B(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_45),
.B1(n_49),
.B2(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_27),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_23),
.C(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_43),
.C(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_48),
.B1(n_12),
.B2(n_20),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_26),
.B(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_2),
.B(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_35),
.B1(n_27),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_14),
.B1(n_12),
.B2(n_20),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_21),
.C(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_58),
.B1(n_44),
.B2(n_45),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_59),
.B1(n_35),
.B2(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_38),
.B1(n_39),
.B2(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_42),
.B1(n_46),
.B2(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_71),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_54),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_75),
.B1(n_59),
.B2(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_60),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_67),
.B1(n_59),
.B2(n_34),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_77),
.B(n_5),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_11),
.B(n_50),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_5),
.B(n_8),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_78),
.B1(n_4),
.B2(n_3),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_76),
.C(n_50),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_81),
.Y(n_84)
);


endmodule