module fake_netlist_5_794_n_86 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_86);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_86;

wire n_82;
wire n_24;
wire n_83;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_0),
.B(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

AOI22x1_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_3),
.B1(n_17),
.B2(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_30),
.Y(n_48)
);

AO31x2_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_36),
.A3(n_26),
.B(n_27),
.Y(n_49)
);

OR2x6_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_31),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_23),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_28),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_30),
.B2(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

BUFx2_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_50),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_43),
.Y(n_59)
);

OAI21x1_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_23),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_44),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_62),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_43),
.B1(n_54),
.B2(n_36),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_63),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_68),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_69),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_59),
.C(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NAND4xp25_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_57),
.C(n_54),
.D(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_76),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_60),
.Y(n_80)
);

AOI22x1_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_29),
.B1(n_28),
.B2(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_29),
.B1(n_28),
.B2(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_29),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_81),
.B(n_83),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_83),
.B(n_28),
.Y(n_86)
);


endmodule